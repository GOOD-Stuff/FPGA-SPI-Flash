

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
icwBRV97stUfR2Mn0wfPioI0eY3zGZJF4gSa++nlQlMi8xdqEhl343ha2TeCedqJlXwUNOMTshjg
NWAZ0CnPtg==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
KdJiATwLz7apgDVo1m61iNvEkKe0M4UdBpI9Yd5Ge670sdg1t/Nie7/y7x7SOpFtKcG79N3mDoiw
bP4Lo28OJmNglVRWiKdTRUXoQr1KC8IPt4mFyf8RW+0wysmhFnEJpQp5SwugZAg4ZiK4FJrJlEZp
aSpgrgqxILRzspwvJ28=


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
SEJEAo+4DoRBD70Ek1O2LvfMayFQjSsQ6O1GJG8EOchOxWL4gH+izXdYttq1qTGn/KE0kJRFDUcX
A+ZQ8kqk+Eda70AyokFzsXsNSPHzlbWGhztR1gvMy+dW963rNBnhXvIDRr9xQxdB0S9wFcz7sOOD
N1RSFCm4eWHHRbqFsdE=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Hw6LuFnFxQVdpUVS2z8t5Yf01nLm9evFIzBt0PsoeSy3+WLcOytdKrEuHuwtqg6ihJly/jHVrfAl
TVavmgD4k59+ZTPqwkyYVYZr8LuzM7Fv3Zsc5/au2o+APxXDon/zrWg5zDCqJ+yGISpVFOGA0MAT
1rg2BXFph8wATddw8zNlEp6bqZO8wbVr8W+qZoEQF6sr6GzqUaybeo6b1Z3w1X7NKUdCSPPuX4db
QRR5bHztRnOdGS2ZkX/0nKkoQdRgAGHSPbGl9d/YRB45phWabAM6E0g7GJRxyuqw+AKvG85eSMKN
V6SyOVpBvhsf3QR2XAMBRIjaI2XLG0cVK3U5SA==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
f1rsayuAPFUtBwuAa6sFvNELSdf5C/KR4epVKFI5FedDC7MXninDZvVIr8Ro+3EmB5CE52O3Cses
OzyWKYv6YZZKdPiFqafxQGdjnlqjoxI1gThSKKHQBU1hBfjbwsxmpQK42hqhWzSCpeRTJcjV1jcg
aVPLy5PWglGMv00FiULQXmmn5GFwuKdr+Bnk+e2BuHMI4hipT8VA3cn5wgWr03pZFoefI8cpN+oG
u9Ot12GyURIz66i6gWxGmq24zuJUslhyvcG/IxJB/b9eaSe9bwz573Uy7K+hKZAT043fQL8TW7Ov
mXUYJTHcnse0uXeW3bie9BUo6EE7Y9TB47lk3w==


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
u0nDmA3YrWcfEk4185AhUszcR/nwHQHMMcbB6zFWjm8trTpyEdJp71iK4ywXp2oQ1lMSKg28ST8Y
GUH/HaXAvnJIVIf9lm4LECEiUiGW8afQ0cwQ7j8ujiLlWTcu0tDGOvezlUc2E0EMkmYd/yAwxLcX
QCiYzQrF83xIvL6pPU5XdJbaD7dD4CFOpFEQRnzHYTDxHZHUu7AGIhYCSDrXQ5OQ6te9Q4sUdPJS
/KiTKe33AZgktXIhotf5HgtgK/xiCoCoxnSbz6PwQCkJfuQJUXFVua3fEYo6DkxeRwgmhGEr+1Nx
RBmwCvu87h7nHZQ60sX5T9NikshAxtWacHhtGQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 1050704)
`protect data_block
JCS1xJDO856PFweCQJzFQljdqkFtWNdxy0PdMr5xRsFJrfCZxILhTcjhXEXuFO49lax56a2Zitm3
vFvo5DyomA8QWULvY9+48nxJKwV4jS6vNnP0uuA2km7WseCRNRVVzwUSp2L3EMptVB2Z3Hr3Fsyc
XESpBNpZEsu2c5UpWR5MjHzun33R5eB9mPXBGqHrM0ag0NJzzIGALU4T1D+sp7g5rbnkrYHXHlV0
0UyXbk3pT/KszuiNjkPbiYJpWj4MIenDoF2Nnnhm0jtg+7CfWSjs5Wwk2FhBYDKzojYZUpYG3kY0
5fCLEanND7LDPg1W1HQxOruH0ig1vg66tLXNmzbfVLgyv3MY65jSMfWj6BGi41Lo6YU7zyDb1+i2
jEROOEUOY+Z+6QzY8q4yLHqGTZYS1/CfbrlXZ6wEDwcpbksbHxPIoxwLa98lbG478jOYjTMeVYdQ
356FOJ5GS/Fck3aGc9FnOiIdJFGD06Qq0qeFc861wEyEa33jQ7s6Pf5SlTjUxEvC4rSuVy0mKFTg
PQ0ANoUnWeN6S7Qjzjexva70lwtWdH5xhiYEvACx2U+4f1p2MDTeuHU9c1dmhQB+RK9/mipAXcZ4
usfJkGXUkI2ZuD6vhCT4bTSWoMplVu/zI/AYgnNyv8esC8bhWh/ZIy1cuIdopaY8PMh7IVDI45o5
EG7Qcz4tRA7SKLldqZ7f022YV2lc/3lgWOVzWLLrJwVeU3wOZBZowmKVKluJ2XMzxWk+wLtcqVHq
BA9TNvPSSOlruardJoQj7chqyd01IXhOYv1k2JRyOFgds/OJG1Nx0GWcc7GIWjrVlK6tZKTtdNMK
OvF6xYLBWeUbSUzAQbF85NURgfdQZNIC+vDT6YpOItxdI8DqcDQOI+t9mEFs+TjnG/XNntbuyvgp
9+JuP0+R+hj1uxWKldnV9huwuqA+vOIE7iqcfBZOW5U2svyjdBaL5c1+kxlgAuFoA5L9Y26moFnF
e2KOVjZOcCvrmHdFV0RHSAMlHN0/aaHrrJzv0XczMlreEmDgHagaIczcMyYfh/WnIDoarUfllAqw
N3UJ+aKrSr+8tiWFTnkDuHHacD0DCrmUxqIKxOFcTHVSxbPCjfcDIytic4qZii45Zl42CpVPXb6B
armTtCqK24RO08O7OCJirUe+Wb7aBjVq4zVsusKJbIFDWcDmWCuiLcIU5BIe2hGiuyGQo/7t9wQa
AtCqd4rRz2cRxMlMXKharBDZBTVURgancBw1AnSGgUle4NObDv0LTGF7cJf5vp5U8D68isDwX21W
Q2iOST96LnwvudFfcgde1NS/uez/Bn+KHz0zVkW/LxZrRsbkqBz0k8hlFSA6S1iCRyZ3JcOHTdQW
FIvDx/YfL3eztrz6EWfdDGWgFN7/5uWeEAv4q6tkUuvAdbM5W/OgR41IM6DdhmIp91e/wA7UNd7w
vwZ2sxiyi+zm+jX//MSnT04zcNXJy98HthlmBkerjsT3ymybH8vqlCFTjeeYhRmdGr6u07ZX5Ps5
yIRlRLLoKh8ZyXavpgTTGvPboKolc7+p2Yzso+qbci+YFjnpflHgocTD8YaVihZilxNoMe65FqAZ
/iHoKEKq7J7mnSu6XVw5IOYPSmK8bPb8LUqwgX3gacXAJtXrnTNZ5EzVLW4qxC5R1I/OOHlpHvGY
Evf3EtM5Ul3g2PW44h2VKd6FTRa3OidiGygdP3+CVEMB+s4A9zddIYAFQ8A+/n31qQI5hiPeZxPH
Y02Tr88zk9+4INbDbtQwy/F8/pvW3dq8drbibEHnl567MgmPGq/3xu2fvW9wFGzQjAy4Wy9pHSzP
JKcJwgtNL9HshXnSxH6sKmYhKdclGgOElAlRF7KfUzeyNIkSqf1RKlj9BSyCbj586Ui47gDVNRT4
BEyPFuAtLTzE1WyyE1OEbL1f+zCl09CXa7PSY443QD0sKfdjpbrLctxOv3j1mRwU1Rz19r2RTTbs
xMrieCWIAw4ZwZPgLXgXRF1mXJA8+InTMttV6puiqJGo/YStGU/KpfNaSNeV/WXJcA08wtlQAxb0
KyW1yg9Nxew8Sz+Q5HBI8U0DYr0biTSklDAOxGs8yjOozyrlQrKtGAaE4xzDfcqF2pS6dTKlco/i
hlDJaDeewY8f8eKKzL+7LjVpC7r7WK+x6WqdwBZZQctaXTnsz/aHxAiBTjrmewAcAgp3UkL/Mql/
RirY3BMoX7zUnKZJr7Wqa8xw5HFvD7E/x6f7WSJubB1ogsCA72MQsrgUsZoGFftWcnRzRks329d/
Ul6GBtN7cmw0jo94i4zfABn06bFjbEKlZePzQi3ayQGD7eSyRxRHTQIEYGECqaCPsMrdThnT9hzE
oQq38V1M+nmn0Xs5yW86mA/sWc4RiD2xX6NZrNeOtBN5GO74KY/KMS4+Fa0L7C8rwS48E3Ks6kqA
w3CP0M1TdZETWgIfJGBfsxPwguvaH82j0E4vb/dh7xGKVjleC69ItSGOutpKKaxEmTVUZTNt+8jD
07wLN8uson90M9b4ZaMaU01gHs04Zuj9qkr6Dl6Mm0q9nm2s98jWeC5j1li/+arCEVndwTaDkZY0
1TGGtzQliMOg6UcI1RHBnc7fUm0ZTsKjDCO1038RjAPrmgKVlCMolsDH/vWBCyAPWAzo5ZuAAwzU
irA7QtlxeLRTT0ByGsK4ex/8nbmXIsAh7UHhRggiKQdIlxn/d+S12wOo3u/SZUVkaKL0sB5JeKFV
8fwpnNgFX5lS/NlBz9VM6BvVbCji+uz7KyqqMigGNZtOb44kENU5AnEBPADN8Ja2wGBMFFIZbfQ0
D0i8DEQ7tTMBB8ax7WsuP96NkrBvqsBnn3cTwERrwvBPYW09LYklujRpNJ+OXhKg7e7LMEG3aAmJ
sBmAfBD/piJELMHbUukWoSnIg2OmAZhpsFdRcZG/KHOpZu5KXZawlx2UOYbBKbQSHgOA0i0qEBlH
g41Bigk/WFNR5W+2yo6+ktQuE61R54e/OqzqyYrpTKBYhgBjYVDaQ4foXl2FCgBYjT/C95iNJRHX
JOFXFgtw6+KylOBoCfIZyDQaSvP/ds0hGbrRlkPVHWeS+EBCvABVlWRdYrMFzsf6yJypuK05hcGP
Sk6I+x7eKmFHp4uPXC28+k6cY3Nx9MxfAQR1bQygYZhHnRDo5Kh0OcFFjQf8BqI2P77pLJCKlufx
2aU3W5kirKs8Ddejh6VOaJ4kXhzfIo4Dx+XQ10zf2AZMKPqGSU/xPRQbFZMMuuxOO/Z4Hk5TfzcZ
R23V53PlrztT8at4CU2TnuAihdlW9FFRexAQZx0QZJfio6MoPKSDP+edYpzZs+EhOnMm8FJqfyOc
Q+LUgGyuwV9IBA5sEHR4iQbUfULt2BJDMRYKC2FNyMZkxtapBLRfsnCgThsNcPZNFklr8m8MDdoi
lKEHRuulKi4zhn57i4p52ceXeI8G2yjUiiS4hacuXE4ABV2vgev8E/Nvi+4+EtuP8jNJxyGI7GPy
Waj71Lgc1w8Kyl6Tv2dkABF/x2JRoo83o88J4GW3JrGJt1NsaH0E3HCuC05jQhH3W7rzHUBTpsjW
jfy58UP1EBCQDz7DYViG2jULhZXwLzEJn85HkMjlIpLF1/LlT+lUodmjm4jWZ/Ir45QLR9S+OAoH
TBzg2pXGIGc91iSrL9zjy9OpVwt/5kGYlSLEfdIsbo0crb1f6vjAjygIwU3LtJ4liRzGvorMIHYi
2ky1ppaBMQc+ypI8YsstVZSzIDtEoiAc8NQ8pe4b7Swh686+IzpFI5axE2MqjjEZp+u8BCOWFRIu
pw+Bt3gJ/782RsmWn/gyzJwmlZrXukKOyaDGpAMzYnhkrlM7mlg5IiDqVzspdv4kXEuZIi2xS2kP
tQHcCoZEtYqzp8AzTvqVfamkUb8UnNJF+Cfg286+fVfeph4nX0xJscYVt2m9WyDYWTA+6viuD8f4
mSO5pKeytFj5uYNfaQqvwiyXWb2iSu1G4bV8YVNF+AO9Kx6Py89RPxQ3yuFOTgzkWRKsIcprQv49
sX8zV6Jd8obZH6Iq2/Tw0rSoUXkTG8DW4A7c7DsOLVlT+iaC8b/F7IzMxnNTKicFvkMle7NHItPS
BXAqc0EwIugkcpOvYhvsWumpPLYdrfXTcalI7gZD2rtL2EEPT4fM4v27WpaB4cnoD/tcgeqB68ZA
QBpbnFw0uT9uIOlBW1X+QTBWRBEsJ0fLqymmYMff8rOSo5KKWP6J+xbsfL+VzkyPc1uAbkcFd61k
MF5PW068BvQYKwdAaV6upV5AfWZUEPQPwJe7kyKzXI2miRBnEvK2Y4QD39eqDb/Ta8e9RX6mpREh
5g1B99q1jT8Hg+RjWdGzhmklgsT9s5lICzUJUovMoWe5SSHuBMDZ1zFr++4r0WRVdSli/ULpyQeF
0wLnycXjvU+JM1CEmliIBl5jALWUXFWNFH8TDarv7aNt6LLO2/KKLU07outNWeXqvH7pFFqhxqrW
N6ofvO6kn/Sjn+QPtUP8wml8+RsGP9rkt7eo6yltnPW3QWba+EsxbDrMcJ025E6MnppnjJKzJRVe
FMifxEu6OCFA+e7evKbajBWyrn2taKwoHX3IWo5APA8fNa75STH6+YfABweAUaCTmZU7/3SjCLfi
Gm197hUZ9WizEf/PMF1c5jGo/dC4gHIwLeojJTSBxKZn1LVKV/0+IODu+uf9l9auxl0z9N0RRZc/
rlwfNxKSl637HMhFn4OGPGV9gkdDqdKo1BujMA+a07ky7nPEnM/PltcxU+Aa6eyVlcPh+gLdlsfZ
Q82IgCUe30JWLfInUNvltgT3se3INZ5SANx2JWkQoqHSLMQJoCP7m19bxiWi7PoL8pFoDLRM/og9
2TnI9pmiC3btb9vXoRcFgfjl5rh2Pv6xC7iryZ2YyHHUt9nZT0UUc8PsDzyrFCDPke6nYDojv+XV
QZGa7uQx57+s8aw8/OqGtdoFum5NcRYVPkzE9Z2cmszLpL+ftZkR8iV15BBMCYsgLfV2tJ9TbKQm
2OUoeOl7LTnhNhzJ7yDKSH4dPflkguWOjLS5tiJM2VcuuBJjpcq1BVIzOWfE7AxOl0sgkILOA1+s
1xt6LCV96syKPvRLeNeCAP2J7MEBZWVMuNPIGkrY8/yZ5BM6ceohvUtrjs/XLsGmsd+HGWiQtT5U
woJk+VCEby9HGpMPHd7xd6Lqil3kSkV71esFaQpZuMbk+SvqAFWnB+EtHQv1mx4lxFKlfPODovHx
5BTxXKheteC5d8SOpmcgQExUFulp83k//FhpO1eHnPjaKaxmdtBw+4scFzzkULo3KWVbtic3OHYw
CykE806PXZQNaOaOcmpfkKg7vwPIMXNzPgfy3DhnyTim5y+ISgVnEdarOb2XLUdiqkjwKlTUex9i
LGQji4L5A0Op+kxbarCISI/6ZU/nwLa+3yTuHdaPex+JLmvsfl46H/wTf2eUD/4tBCeF1Lo1a9B0
QG5AdF8Ji+GhZiyf9GQ+aLnPCF52s2zHzFT/qUQuI10xvUeax6b5rxf2Exrk2nA7pHqbU3jA/O2M
irtwjt0faZFI01uSp/LaGPP8FdrU6/13CbsxZesu15gAIYGrYSAZGCF+yWrnFhx8rw538RH9B/Xs
oawBA7/KU07mxTQetVdTdEVWuZPKSnYuH7K++59mYl6Em1MvE53MMvjGcfiL4HOZ4zhb2t7crlrL
mEWNO5WDmYlGUmQKfc5kI2Auc50eH6e+VX+93PGJAFNrd+1cooslxtTU2t1WmKLC2cKw4VHkVLiS
7KSa/A8Q57BlLjY4in8lsBy0+vkecefcf97X+yqhn9sx0VShbSImUU4l6gHVqfhlrBk6pmNiI2GB
FCFi610iq1qasc93jEwQn9RwpH0U0e1NMZ9nJfFAO0WTK5p4baZzyMYiD7duEDR6E39ohJc3HIUv
fiiCqDo2mSNzx/q8fBlwJYfx7mT6k34koRVUNbEgAj51w54Yk5NxONPxJc2Pg8Z+E7EqPj2/gZjN
FGtsU2nVwNdeCEgncFnzKrRsv0ibyjdGnai0Sz+fUFZuavGRCKXrDR+iUTqDln7aXsS68YbzusQb
aCU0IQhfk9rqfLzB975SnW/fsVkAjx+Lz9JQZjUawNQfN3vgWLX1RSbQKrgmgxi9JsAJ9136Oeyq
CvbnZWcHYoqQ5azII4XAuN/fkYMqYKmeNZzxjsP5OZuWKJ5P/x7edOmOoGQyRpZxFkc3mSE50AVm
OGV/bxjMrwNYitmrorcyq9Jk7tiECheoc9/tc5G5T+dvecuuGQPzAdVPRL9hMksnsq37NbEA/qqF
ciI0etkXLflbgxp6/v+eI/eCoB9p6VwgfEkiC9Ogv4euDtL43eZpq7kdohVY39vSPwPPOzPysuoE
kdUgLenISczN7wtxZV5sCZ3XFTtfa7rO+4sXITfqEcYGGbLuTQ31n6PHlYTMeA82MUFAFakxmE/b
Nk0J5LU9PNNBLCUIY8O77Z3NYKB/b0Wf+2izIEqKCxTiEYtLhHWgyz/jfuupp8sm23a/tpHd+y+O
fjziIWVUJcCth9rxPuLdYr+FqmSSKX5fkUhvPI3pXYm0YNamLP2nO1QpwnV8f3WA8bJcomild7wr
P+nXIgMlwA7liNMjt17QlBUEcgFWyh8lG+D3o0Lt1H2HaM1bD5kU3ovj9We14yD4Xdi3BUa9VE5z
6ieneD1mZsi3WMVi1ogUw+sV3IQQY8VCBENL6QFYuZymI7+PWNdW7aXl34dDlvshzDLcqKax3+AL
Dl9/ePUWBYbHDix531TnCSoh2/ii/zI4GFRE4q2K41MyY293F6u38edVwZ3F7oCD7M1MLB1LEVAf
IP6OMASVmGhXcN7Ke4JsmcpBZ9FTblxPDpD5ESfS0HIeTC12Z1lQ+lTLF3cwkpW2oS+9sk4kw2v+
N+QPA7CVlBXJ3VfTydexpr7PKF7jspAn1utpKFtiBdF+PF1brTfhmYFlR6QITusYmP/cj4J/GMW0
QtthSsc8RWVwCTz5FNSFDWSX2lU1DFBqlaCkaxoDEjru7/Ic9swmc/9ACYWDyCXPDuTBr+DCkOVx
0A4Mmhzvy2n0XufEMYtWnNR4Ox4eZaneUQAZel6EDL8epaOilZuEBHfjCxcfG6m1eHp2nHd2Xo9Q
bOZh4e+eEoD98cd+soV+IA5fWWjc1iFRXI0ebTeKwjdubpReg/lyeWYyFdGIE0AJIITxx7vz4/3I
+HjySY4t4vnBHvWp/ukdUakwYsBrGvWt9AnIPMfZiy8yloEljiggPepE9dDRHIwibA6bh+vKXyW6
P1Zlqyi9cynznhhvTCN91IPsUkfrmXit02dE+aor0ag40qYWmXY4lGXMiUF8l0/j1KxChnOOZfxK
UVcgjIYQAKBCYdkH0G2s2OxFGDARBIph6eTtoyJQyVlYs9jPHqNzP9O48GWDXyhaR22l5R34BtC2
QEejzOHXSd1xmzCItM+A2QAARQ+oJ00QkQdHvc4VYgKQRxmuiuJnc6BbQtEP6wNlYeYca6n8Dn83
GU1+6IMXywcufW+mGN8mWLCqj+2jzNwwAQ8snAgfWCOxH4Xg112++4v/O2M8jCbbAENxw/kwvXfh
THT01lSKCs7utxes/MWAuAg5cZjmCHIyF9Gt4O6lTEGxtJ2hV+3PmO8CLp/LaTw2xPu4rXjosldg
i9Pj2jFoWsSptc/mgQ+DkolTK3QgtqdqFd3FI2lXVAN104WeUg7v/eIGf+sgBmyOrmg0baJY33up
h3YS4YDi5u/4+TeHXVnyVe+jSFkiy8yWrQxGZYnScvg62jR2cxGvEGWsZZA9mZanO76niTf8Nomm
XLmKIH4oYHXFzd73BNaatcnHIfO1D45a6IiNRkJvrky6gSXnb4NmHel54POupMDo2dzd1s18cFr6
A4cMcamtKkO041wGyI1t//7k9ig74sHKmD2FXPdI+RmM5yuAoRbW/9kItgPaeEM4fE2URCjERSl0
GMbLKNcZyMDstTvMHz91QDy4sqTDRMD0Lg/g8phjmKWvEwnIuLSfEo6M/lgkkbE5FINKC+EttS6k
u795iLm6HxTr3yFNyuVwV9OmcTX+HBkdXOgCWdolF2JL0zlrWIVCqSLdc7JxBFmWgFmTpbthVSkq
hMAN3sEj/abOMparIkzrzPAR8PE6+XsMxXbD3PAp6n4uvZ+052tKOwdRp5hWEDbhMbmNUQCk6AlN
yZGov2/YCg8yLwHipraOuR4+x3ZKGSKLYZBD4jiZGS7H7pAm/QJkTQi/s1jArUerIqt8X3oed27n
c5rdswZX6T+840lDATRek+S+MbLWNOPa8r6FTbnqAD4fnERnfVkmFu2D9Av11Wu/+PNa0Wg6hx7O
k91joRdsXrVWfYg6LDlfpJmDaWY95rDGBKLj3rRLPI0tppNbDHEbqHQqE4NfwP0OAA0YZBFpdKaC
+tDDaw0uyu/DSOfUxYvuENeynqmhAifa6gBP7RcWNGJb3dhiR5U6HwZStP+yh5S51QRcoZi1u/Qb
LVcQ6jJZ3k89xVn+4UKhtOOleD1HtoCQajiOt5jTl20eSb8J1EOP2c8I4VBDY97FVgQoHRGw7gUM
CpWQHUSpE7Y9L7BAu5KAJIp/Bf5S6YsWfI5DXDkuAes+t6Y3AylrJ3y3e3F7zlDe3gOGrBJL4KGS
8EmEiseugJBGoH08JAkJVSk5mm7O6AUqt877g7vLRDTC5qSKb0CcBjw/AZ0jf4qEq3IP3F06yyzZ
Cg9Ift8eZmIMOmjffarAfatWzSiYnyeLqe85wZtFwj5NgjM0jP5rDC8PTxCSHUgW2XwLT3Ys9phf
TtQHi9J/7aZ9R5KnCACN/H5YR1oZqxyMzg9DnNHlp3/9hpomUbLo3g8VPiENr94/rSXa9aq0wqxU
YhgYhBv/7hLr1EmdooCFmNjjDXEdrSxBBviXE9MiZMqSw49yYWDnXQ1V1Nq0BPhaqkjj8swq+yq2
KxuG66+ciMlRbwaGKS4vtLWBVKCoRxb5PdWEnMveZp3UAIDOC9rlRJKHiNxPhvZ8hvho23V89Jv/
9KKKSqeftke+BSdVVXD+Gwai5UA84GksBDxBPzy2BVJaENg7k6rolDCQR65+LFnzGiPLukztprqD
o6L03Nu0qHqZPDWSmpz6idW0eo9BRK3P1fCYPozVRAWR964bP4Ysq0nGki6vcMTutsYM3jMtOPGy
5GEukeZGHnGS0+nNE7oa3JIvHBvLGNDlQbHSvsPw0BMoi49jPful6qCpL7jq3NKFTleTmxAl+lEd
r7Natb/GEKHUGt8EjpWlclg6ub6Z+7qXGPAWfRb8OprqLImGwD2DcPLTSB1ybSyNifQgcpl8b/JP
slp/mv1tOJmZ1VrVtFY6vae0UVNl+5tGEnXDcmMpu/HIeCKwtCXVIetBPpxzQHQRGWGlvmUveYWd
rOgEQ8zlEqoOi1V+j2qB5vVTAVSaK3lDzU4yl7tDmO4uVf+tTW/9CX8gfbFVM+sZUDa5zPK32+5p
0MQ9Fmpp0ZOpGj+NmILE2xRJKuqbfHBzKd7chQrdJMF68RIWCIgp37RZhGGZKad0o6tBXmo6P2Bu
slBPYe9dqGgnhv02jcILf2UOK2SEdptd7HrjQBMJOTW11YXCmtYkjcXAVBICXIV0S/sP96sb4q07
pU/6tYKd93CJ3MnzjbrvDrQu8dIMBMeJO56yLZzs4ZNF8AgYQ5J4KQKgb2ziPlagSY8LmPQvoXvz
kTNTXIVC6VFk5aMq/zgjGCv6tF/YWlrJWMKx2czOX+QjbrEQkOfsqZLIO/rv1OnwUK2rQy8KNT5v
TU3bjRsNQImUBEHpGleiSv5x6hCTuGf0PR1c9jO+HqLnAXFk64y6d/IP9QpWaBEb162ComIu4gYA
jItIPho9L9SKnOVPJgyJnPq+RzNRJiQ8UXDcdOnbvC47FQOXjtBnrgnFxu0X/NoHuTd9O5KP+3tX
y1j1mto/gtIsp8QDFqCzIJoYZmNSUOFGgSt4NEkevKLzSqr5WFqwR8K0KjxmLeakKjf1Ci01R+YS
zso64ZM4oAqpmaY5UwJgS3rHwd5i+1JTU8qXCkyQRLfW6v3A0RMarJSpMg1bIjFoCyBUMrB31OO8
U8IsKcQ/HGxpws35OwLRhcklXIrc7gvVj2oUiruiG+4FnIuMNUw7YiCgITyUQqkUn4dV8n4dhSRH
ecA+2Ljc83Ez3E6O6qldGUm6sq5Ubdq3ZugiBwMXl9ARa0Nhqm9QAdkKbLRdZxVCwHoDvzoFW8qJ
xFCnMSoBzzAFitREeE8G8RCm/coVVJ3NSO1S3e7+mO8nIuH65OKX49jg3X3HLswv2jVGP9HSZZ+I
hUlJCX3Z+HwyE/C0WMXxLcy0bb8ACz3r8uoaoweJh6iUcvx4q1HoHdWo3/KWRGXP97Xn8XH5oY2T
SqWn0x17NKQCqERDKYIHfRb3m1vvVbTjuvwXFOSen60rMQM/Wor0atLNbY0PLhXR4eRhRopHHTrV
7NHik3hOA54Fvr0g5Q4gu9qFP7yVVbpJ1xLafmSR96eh5ouwItbutH5kvN3ZZZ+vTW9FQRge6SDB
3ieIzepFrxlNdNGNJZw6X5VaOXYn4JfD1Fx3Y6dadzOOj+8WBAm4x1LG90VbcXrHyE90J0+UQFd5
+Myo500CbAJbhk2Qz6cssQdUpd5P+/kT+w2HLCcdV45sy1to/yyKmZEMxvgJ0Pwhor20+7Zvz1uz
5YEy954N/7Re4wZSD/SGx7BH25w4apZQar02XxlRKW261zgDSg6qndoYwYrZd7sewYvoUcIBST2B
ZBaB1qsjNn/rA1VxfhUaSkwlpYz83wzbJVnPvqzRFpUyh2HRcx4d31oLasBFkO9nIGxJG7OEYEfl
vgunQVVeIVKTOe42LWxkUkRrvYjMQqs5dX0lYic3V8Q+AYcpQNilAKy4rTEF9vluvf7Qa5wtcgzD
hRn6dehIGAaBB4lVKxXu9oHARt8rkhdBfgFtdGjCeeVb+Grg7dvpnL5LarHOxf96gaWGKvHB2y/W
LkY1hSMEi30Ue3E8SuRRihNOhl7DCk6zGyUb9RxEg0KkMrdYP4BJD+aGSmQp7YRL2JrOZp8Eu+fx
m4iXAovKHvBTxpsKrwXjHMVZdG2+rDy6362B/G3Qr60Du4Z99NWFq9Bt7M4mSYq9ltl4R3L7+xP9
K7JaHWgWCKbzDgP5Y1MKlLTapR0AR51Zvz+SNVrPJsyYedATjihxMcphLi7TsbFwTrUcGjHr8ZMy
gr5TwmiPWIpWR/cfsZ67UNlFqC9ep3kF7OJRIBrfULC/8OKI+xJrxRemrOGRZuIxUQrEG2dZPbeK
QzVV1lB1dkxnRZndVYslgcqRXuR9KrRwUtjYFLsHrNeMBssioWf8FXAacMSy9hSMh9mqH1xi8HuX
F282rUfXvYfsXHM7Y8YCmIYLr0DI2Ugirrwp5z9umqVgeBJzmO+gLi2LHCGzSxaVEcgdFTYFUwHO
v0qt24MJ+eqr3dIUSd104ouuQ7Vjqgb7GOgz+NH2zQrEgx8Eo27KER+JpdMW5ETJTORM6esf+eOy
8pZrjTxIH8fUmf9/uxViGj+Rb+OYKYRDak3a4x+2ZGC/5TKEkpR4arlUxrFOMQXIRg4IgrqOEUhC
/uzZTGI3JMmEv/Vhl//EqWR6t+5Dvzk+bnAjAOtwXLiFMi43Ds6SS6hL294bZdPlwhES6CrjCl0t
8ziBwH+nw5myfV6GU3+NMwzyRObz6k+OcHBZEcoyrK5sY2ARqIQIgemCj/ok0ZpXXrxLMknumpPL
M1XW3yYbb+jj+cfXb98twsPsAE0zEvypqbaxjcCTZbIagcnA0BpAafiraNPesWbdBzQSWiPUlDrk
H9Og8LlO0hOrp2x2qtA4PnYneFhWHUnAQHRMpde5iKUfpgInD7v+YmoGiHSCLx5UoYuUNhPK/qLd
vzGERHhmDOtjN00onmVBestZG3g7vWHp617eGfJMsa706sSTYHAsm/zNd1RBeLKtbxEa854Oq0nF
sNEZyeijCH4s4bUzm/sKRnzhVg7klVtEh8IU5ojcmCfWsOqUlRFd8jjbxHgYy6+xg2WNzi9B3Mgr
GKcQTtJCGLqsa/ilvRKVTq/YgNPbTtyCcNwVhsYUEdi9Fc3TmOoX9zxyWPKYvqzhJq8rYwBhYV4z
Ey2GmBZhIA4JMTeuzHD2gYxSwJCs0TUfYKUYNpzlfx+AfgVGk4P9auL7LlkoG+4pDSxyNz2PKiIi
PMIqSqnabAwOTvjzd0QosQSUDyuUEBzr7W2TK4QHnMIfPPiLGQuaqrixzB7iaPQ050yeazGCmnbt
/FxTWf7BDyOabIg+8mSSiSgD8PtOOsaXfDPuuJInXgyChG/FWtM6A1jHy8dtdbXba8NtUHZ+oOzP
zy7FH/uk1MP57Zt8bN4DK7MbcE4f8d8w4ZL+kaWAXY33D1wG0jzGKdmatQk1ID6MLkvdu7Dc0+M+
AHToc34JdSQ/2IlILjODx1G/vlRjVp8hIVZt09+Ns0KYQPOWdht17H6jLyp1zF85KO8ZLgKTg2hz
Ohf5sKJo/evzk0ZwB556BQQJVJyUFFrHSK1n4c3lzVDlFgFP9nD/n4CCt9jULqRWoGP6S5KDoIh5
Bdo0SzNI1CzoqdfT/XoHwkM1AJUfmofvfuUEo0xstQIQEArjBvMffn5Q1PELozRXsB2vVajJmZpD
ke3d2e+/RFCvyLJeCJs8AVLheTXDWUO/KTzfYkbBNweYyMunHl51NrRrdbx8RZoH+a/AIv6ydE3Y
SIYoIjcZ5ISYBBcFVfXdccQajPBvKxLLLARveysxrDZKAzQUMMi6AYfLH1UY8I/rVuQYf81p+MeV
qxOsqVW7VlW4/BKJw10pYimOkdExDZcKQj29wx0CerooRm/w81k/9UlLYOm59LtbAJC984wtIOy+
2dMIrM3eDc7j3UewRVt8JlF20qfnxFMgHY0loz5YvjCSBT46saZcAs3UFj0aWUsYw/HsUebAbKrq
IOlVNpYfomMzVLnZeDBXFGgfRv06zl0xibaWss0yxx8s16aC2QvxHmGPbdB0jFgHwRgYguPpGBCB
/INcaYv2NGS1cn07skn/4W2pI/sQuuz2x/9Y6VV0eUY5Nqh3FCAfHIzyMHz6DTxLys506JO1JRtT
rep/hOpa9gcQE8XDipQamqa2e+3RTjSzR3xcwL4bree6cKkahyJEAOOfdChWnvSSsj7CkjUUGpka
DUWx8IIe8dHhv0tb14EJ+yJ/l/RWcIfDG3rSFBeVjhhfMtYjsYCjxZl3S4HdBqcAHYLaEGouk/t7
LUeoHIXdNkaniSQgF5edAFp0O/xhn0WmPHMm1tgA5q74jfpXSmpAYIMAL4iouxOQx4fKyXi2ouO/
sj8MqHZinp1Sg8l8/+Vu6QQsxyf6yDmLV30DN3+kIo0Rb7COSqJz8m5NSlADrYt4eI/hjYDdgutH
VWrKEGiLA4u+Ew2Eh4ZVCq3f0s5yTrPrHGeqdWwIjsmwMer5SfKFx3SA2MMaa5PuukuFzAi7FDyK
cppXidecApnDCBoOQRVgv45qz6e3DKpSNnaUVPPDNkbNvJBx1GGvCcrTIS5Or9uT+kzNaO1C7Qsh
vu5dNt5qUFl8+3wT38DClD7L4lWlUgTxI1PIVbEdfyehlqFFDf0ZUJihu7GDg6L3TYFh15CB3ZhG
9Yl3ZXbBR8thSyXqXzUOUIIV7F7q1LUbmEbBmzHv2qqg9MzkoK+PCqkmjKH1BaFSaJwSYWghD0bm
pmpk/mqe2HvAJfPj7gcZ+ZqDZG2v4izYjqB1ChTyaewdeWaWDisj8yQXQNcdlL/vgB9TQ9y+uMZC
ON/4wVLvRNdY1DBS0G3pOSn/OK8wGIci399SzJhJSSg47mI86Z9wPFchpqRxs1e6yJfNeyiJs0gQ
wx6YOwE3aqI4KIyuaGkKYOwhHfSbMNFyM2pZrKFtw1aAs1ghZkDowvN8qS4R8c8T1hACQq3xRWZ7
ry/GDUxQmkgYMJZniNgbFBIzQKhpdNf9a8djITJSCVPN9cJoac8AaDJs4ZJSojCTAr9k1v6Qkcu/
lIYU//cSITUzPp+yfPJrjt6Qu3+rREpRRhMY2L+XGghkFVaqfuIrX6hDVvEmA/WOeX+AgSffy0+G
yXv6GGJ7JikTIoy/RtTieB5pBSMvNN9jsV4MvdQL4ZhoyYxMU6HvGoO62/mgcydK9DTXcBOuHrme
uYImI56+NAIWNCamutuv0ccniWkRcU4KzTB919yiotQNvP9XNHzj0XQ6lfHRSbYBZMU6Q288suse
GhwxhxBPX+a/Y2C9AeIXU3ryBhGmOjs81A22ewEULMVukOpT+6iqRmZrXFaeKqj+25SWUzoZ2Y2W
NgeU7SBKRFVT+QwUNbwa4t9fkHh2hZ/ErXYxPRIQB5awh2CeS95rhdl8KdHBjUKxK5MvwbDTUcVZ
a9Lm03Qton8xKYzpkkijq5t0AoXLTUcm6ap6iiroPG17qiGq7CEg2O6Mq9y4wD4PILoAsEkDIzLg
th7nJeC55AjoFJz60bFOplNzEjG0O/DlvU8dayJq13l9Xn8Qd0FLmGwCoIJhXlgzb5ptaxMXTlTE
aDd33ElorGPc8c+WTf2PhkuXR+uiHbRVNQflEwOXUTyPgsziLMkMnee6LEQ5J73fxn4Oo61C4ERI
hqSAg30LfDBjcQWwogCgdvRT9fU+JoBVV+MkIErDsliUolh3RszkQYquzJo2YXV6Yxs94gcvYkPq
5LRiRccDemf7iI4wHj5YQNrUX/0xMdHYOTCXBA+SUo61+DeDUdZ0/EQORlYLdZUK/4tNeLN5XX4Y
fVwWgYkZsKPxZ6M4nrubHRJlzwMlvHo2Qx286rZ8Wjt0D1vWCht2QTJXt4djDPIq9k2WKks7VUxN
Wc2n2TNQLXnizVjHTPbPmVSkK9ygG03dRHvk0tOap6w3ZZBQziPii12GJrZ4yoswF/CgmdWSTkZM
RdI8dDVvRK52CRU49jJlYaw4xn777sXqrCRe8kGBhC9KuxgOMMg/FPR3hHc8SE/LAN2ZM3tVRq1Z
H7PLT+R5N4T6s5Ew1+ysw+fnH3niafFQd7+o8tGDBs5HP6lRDCaZ4bbia7QyQ/DywC39hy/EjbdU
wfHGXMANlN+sPDYYhNyyETpaPl9W0jWaonaDa5DfLt1p4CRGcsm0wBMuB24fM6zhjNWornXXVY8o
bOkIl5HS/15PCqolVoe3yRkuczrt7XEHt4Y6ftl/vuoZ8gvUyCNFJDP/plUav/1ar1JXWTz/+tz8
jsHo5dy6w89LKU7Glhr6S7poyf7Zxhv9Mo0RN/GJcuZMu4WHuU6YTkWubigslXsN+9kHT+enzFR9
MkJXhXdPFQdSXDU7gZCYaB3RJPbmABf/EDrvhQTmAWcs2xj4Pq0V5hIhsU1ILC7wtMcCvfSn0p4R
RtCj9+0W1Ymv9qzF3hb9M6XEtTPdw/5Op+y/17P6Qg+fm8C41r4KuXHm4cg5C6IqWdwGErU3R0T9
+maX1RNhYnsLJvacIMAbx4oLO/g133FwvH+1AqeA4v+DJxjb47cHsG5NT0N2eXqltuCUyh8KVi3g
4zs4W54ohFJoZ9meRDwdvjoEZVQmRSJ5SSB4NFwtELEzCUhbARsTZVtSTR36xlZOLLLkbfm2Yy4I
ynPT2Yg4cSCIM9KWUCitEt8dQpH7gAF+TujKvixZ9NKTxC6QV5X0cEq9pYUjHx3qrgZect1TFOy2
N2jwtlXhpGAIqC0IiCINhhO09c9M9Lu0ftZCwz1BcfO/vB8MWD/VvuaQ4PBHTRqksoEJ28NJav1G
UudM2mhCloCZtvCx6mmIWNEePT8JnD9A77yLb+PjVbgH220xkQXUwhgeNB0zZ66H2iVAzTes0Qpj
ZYwq8QwBz81uwcVfpcvdGEa19sHY6WBddTUvi3mqJfPbw+7FdNJn08Klgm5hlNR0ZNyuleL3tVLM
51gHMjx0ZAUH57vyj1TjF7WeTQbNdUscc8Pnbp66hnamtasJfBJHDBX1lZWgWPYUl3UIp5r1Z4ny
6FgzOVCYpOYm17++K3DTyPurFTtjTcbncESLKz23iRB9IKgDcAmQnJN9qksYQb0PmkNoiROPJNMJ
aMl/XGhtvWRxEChCPCwvmKjmm1AAaBie+2VJCxSZRsypNG+MdPEEIjU58fN1a2RwPDpOxiuyesA8
hPlDnZj4vthqDB2ZXsGOZi1NQPFuDMIDwiJs0e07PzHPWvIqDPrNEYt3znNhRs+umjSHjmjeiztZ
WTvP/gX6v5LgqvI91rjCcHUZleoFxnKC+JjaTFt6ShKyUW6oFJkIGpTlMAzEvwKFT4h2PmcfHijr
diJDNKeV2VPtv0Vr1GkXZSTK9INceQKRblkxgE/GHa6FfVKccaFrmyjA8s37br2SoNWEar7TPHtx
JzhgXdBRYZkvNHY4gVycMhpqRz0jfWubY2QwMjSoD+qD2FwCLrOlsAi+cmqDOpjcECqqAS4lU2M3
RyWFqXaYdNeypHRlZ4sxK+KVxELzihcCbMSgSQw+k4ZLsRIiIBgTd/ngfR2Fng364YqeEC3zosnL
pV3oUR39FQQWCp4EHQTw06kmIYaoBYvBCqjvppi68nO1kH1fY75Yf5pvxnLgEHh39XgQeFXDC+x3
4OxtV+Qbhh17qor996rVIXbPxabGlYCYz0h0WCKrCxoc2kbNCifuTqbf/x/H3Bz8ajpj8+Vcccvn
sIkEMTy8LurJ/njPkWRa1HAp5hnZcNX/WdmBj531ldhddrX6Dx2WHORelTF7ay9G8h228/+KRrDJ
7xnqE0G03eu6xkhhXOZIRNLMSnVoNdA6IlkZsQ8t6Udx8UmHsG3rQoV32o/DlYvnCJHrQqSDTDWL
R3f8smCgnGb7eFDpn2iMsU/FYxUSAte+t/sHcSmYc0EApgxQzjClY6r8lGYlqBQJV5N8zcXRsrP7
PVycEg5jEuCJXhUbxn9eSKCkqO5ANrS5XA1veai/8QqTQnwJhWlCCMNeMdzu53roTrzSu82kJCc0
w2cWaQgGB2Xf1kUSFvB6qutD+4RWOeuAY3Q0sH9+/7kvyfH7zCjl3KUxaxaD2mkwUSuEbrrpvEzd
ZInAyfgf2mVJvzXGw/qO/yirHlONxufTV4IC/jgD9uvuLpBBPqSJkugBTugZMrFfsjKUyGUNsk2V
pN1uHvn5PeFB/BePJzcpJ5FS6i68iUbFdPGxMwB8LI1D8nV6oVFFJ7Pg9xsv10xl3JtgulhaOIHl
Y3zP7EoAjeVmR7TttqQvXGHUGdvijB4tvmqYqzE/rexZB2MyOl8UcY/rXGY1VcIFqHqyktqWtIj/
Ezd4RhJ3ev3LIKPcR4AMcU4YnxIWK9y2V6RUbX0CspGyL5xjuBt2XuJNJBAoEX0ovImz1SE0uv5k
vbls2TI42sPMC26oXldL5Ax0I6z3abwavkJZYBuoBz2iyZiA80sOiT7cr5Gvg/clQcBR2Jr+3kbo
qOjixgaSKCz96JfmtULcr7K1av+gvDeU+ORovmVkdNoJgf/CKuCJ9kBxIOgfU2ZMvzTG5SBvscUS
YaTm2XDSoCb7uMKcZJqKXFX+GVULfC44ruEVeCH5I4AJVpsj58xIAKJBv/n5G+rNnG//TTnOW1dg
VFwghhYmNOVGHSITi4aqBWP0GCGr1zYPwiXGmtxL1eC9bNzoQ2by/FtKWDdNrZOhosXw8aAWQEtU
+Xmp6kzxC3WvSAxm88mt5dlJNYHm+q5uUn5GacN3EZvn9xi4EGTuOD5ymIC/EwkZoWG3V863L8n7
8Y3QFnIb4TM72hY9n0XHZoB7eCAqMwZQagydHyK7Czkgfcmt+jnPkZrPL1nVJoHPXCjr1iOtSP49
kXUpTOdadLQJEk02d1G59xzs9Qkn4QpeZxYDl0E09Cf5Lui7zq3f/utj55MxLi9JYuzUxx3B2sns
q8XWpaTEOwtSlIEgvWBYQfHJO/LnPd2w2kNyfftPr4gv/xOjHyM6zU3aR96LeojOYR+vu+QEzCLV
9CBYsG1DZdLSP1oRwmK8bCVzrqVT8Ldl/Jzgxtl4C5/Fh7KsmTnYoBZ+wxvFUcfYE9DeRzYrOSQD
u//x29XWS+7r6x06mnzHcK6cZjFUnFo24K08jtdO95uL0v/alhI/ZhjACrW06/gieXK6uO61wWIY
5Zy1lbGpKfbvxGjs7W9mBzKOUCjtnb7VGKYQw5Ha7qBZdfw6ALb2WO3Wg7sWyLA520GJ5n7bhDgp
ZCWTbyI/1mFg0Au1NVmqgu+X2zHcg7x+5TqjgfiSh9OWBBp+HDx2UL4Ni/87LIowmd+EQtLo1WdV
cf4EMP6Sqe+ucWdGTfL8UYstpoe3ciJsv12MbeuPxpgJreFhLMzehvOf21LnDwJ2Eh7sRyUozIna
Lt4TC8VpCrYfBM3dAG7dJo9pyf1lGXyqlJnDLXJVwHs15Uq4hrAtrx93vxM0LOnlVow9FzFIUz4o
AxwT9G2QIg2ZFOF/YjEE1dWMWgOvPZrOtOcGC+SGey056Kxz+9zGPZ3tGoW73gZnKqQhA8CmkHJo
0jyZsBR+aDwz6glFu0rdvHu6Z7EFxpNbgXj8711Y8uRzyei+fC5baVUnffLEmR+WOYt5GYEZU+b/
Kg71SOPOfLiFzZai3EMzBz0WAhCuPZsBAAwnU7IluNrjJ+ansnZ99lqYUK3HQxHVyOpTBxu2sPTb
rOTIxn4R32xWc6MDZ7ZnMBEUSVQnE5viJwcqNBnffwigfhHCVLKwzf8IfuU1u2jxudB0GzPCdpEp
ZTqoUm8itZVOfB/7vIgXI0SG91AqtBTUkqxzIw+TwNLtXI0n7o/JIv28MhhZ7liDzX9j4PL1e/49
PrKuOg4OqhbofUzg45CEMCftiBsT6oCAUfuBZjX0RifNh4p+bIefRqKnmJ8zLzSMWN2J0QH2xRu5
/IeMvUc6F94os7gA8ExJA2Hi0/V2kFzS39LLmFN6y7PAk+kExtcnRy2wYy2dPiaq9aOTUAio6uH8
0IsFiGeT29BsvKX1tGq6SneZDHUocGs74Z75iBz81zpJKNdLt+ATYt2zqzS03S1Y5hdYKIrVQBBN
sLnRBHmmFAB+EQI0BRai+Usan5STg0ux4RpfUX48RT8f+fAuEnKNNt0KkbZTJZoYo+zbPYQEXc4u
JMibJeIcqBjCj8V7YZNWdry3dK78Zwh/GmZBGHa4MBKl4Nli9q92nolpkn9sjTraiLZHazKiMg6M
k1DaSMM5PE7ppJ+UvBVvt2F6irjdhXLQd4PhMABI7xfD4cq8W2o/DRPAAN5CnjXZWILr6R54Ahnc
+FKQyrOk9h82gwX8G28OeEEMm09itj44dnfBxJ8nIOdud2SFi2lI0pMR64ZCWIL3g36kB4fr3AjM
iiMH8TfrGESeNzoHXjCc55tlLWOTtQ8kdEWFdV97uFkx9oyXPRWAbp+A/FK9pRdw+fs2vax0J/Gf
Bbx8vh8coqbFRDNYKjIeYCLZbu06LFC4pHF/GeLNox8mdt67Mv2CKul9IiJQC6FLgBshyoxDwzIg
loyTMDcgdJ6qSO53k7ku+VryuY/kCkRKxMxyTQ4C9iKmuVD8Bg2vssPydRDIoLrgXkSwvh6s7EuG
IFHoL2zzq1rbycISE2DtxMXgcipzrU/V8a3lMKMg4wQmN0J7Lj/H5mSpKBNU0xXZbm0m8DlS61/l
4hBG302LE3FEJ2pcTrzzirMrxkvZsl0pnZG+qiTe6b+PZ7K1OrFX1vIEpEd/rZuBteJdQZj5DnAT
rUYfyGZRZOn+RDwENQEZioz1lfNRKD9O7tL/rgLWcD+YfuEMw3is7sq4xcbe3JeqKcS796VrMV9l
RaiuF7HZgYJGLUJUWL+JeIm3d242j3JkXZizaB1n5YzYW1X/rfZwoPlEf6UeE7P33qRdYitIYBkF
WGCkwA3opRx2mUzY7/JSYYG6Qsh33MzCo82NOI2cmLxbSdkzng39etTgWBAgIBN5EgOl5knb2149
48YXIszl1pYK9ejmxG4+Bp2wb/JeoZozyGhbVOaq5zXj/SGBACrIg0ubs6felPSv8MnLixF3pEDr
pvSZLuSM+O+JO3sdkDqn/yWVxyDeglUuFRBxgc8gFcd9IeTlj31nBlYN68YoRCk/nXOZJahW2D4L
KOSwf+67QgFo1/U51wyfVxb67RAbsSQN1OR5tiT9VvimoAWi9sPjA5N8Vs7lUsrvwPYsJLpMjlCc
j9/gOfY88orD5fZ+600wAqZftv0axVyhANSKU+xObQyZ/0VTV7/voiJmEVgVPX8bsmx5H3rsLhTm
OaUcPYgrdnL0mtr1IZ9QXfikjDXOmUGoZANDXbY9VZ/s5ExaqzsEqHfDAUBVniJIMOiHJLs8Q9wO
ObRuSUiv3AmD+jNpWDg1qpZU/IwXwNKrCOkv99uApvvb+34ONP1sbRxpGsPnWUGiGUma/9tiqr9L
VY2ENGE17iniZzgKeunFDJLDjWEL8xu/ye/MM23Q55sp+DtsEuUlH6dh2WIclkxIGwBVH5ILTEKR
0oODjLxNdtmjHn1ukE7lIH+XOrqMVIVAynhwV8qe4mCjZ1IELk6m2e+ckQ2XzPBs8xLij5kklPnT
GOck5jtPdvjPCb8qi6Tspt9IIFY3EaVRDtC+SLTxGvercgf0qY7kHoOKqUDhjL93DgekF3ss15TP
OpyarLNupaRXtIT0ERjsIisOZax8/0K4aXui6n/VcKoRzYdyOdb5KbxmgTRmLAO9uDxmqtcO1rl3
tP+8zlpRKC2IBNgUzXonIA8VdTkqE2gZ8yFmH6gai6CC38NIe+9/Fg/EJmZ6QJFq3TfLEbdZJRRy
7GN7jZkNMOYDt2QX/1yq05AZ3Xl9vgTi09682lkXqeKRZL1jlxVR/ssoQHGWFhcrTeVzfb+5dpLX
4cUtlSyuqxhN3CC7ltN3Y3/re2VKM1tQjpKJH3phH2zReK+NQ6PtN/HGtwCqYhLz3Hfg/3clMpGR
6VbIZNCU+6phxaQ0GPK8wdafxC0hvKN6wD8HNstBbr9aMp+4/XEOH0pA8vGAlZ0Q33UmgrkGrJsp
BpEx9+DcgFd86+eJWLJLQNeXnvG+9Q2Bl96ZufI9iWUsoqJHWLc3JvDmyrc6ktYCZPfPJaeDkxJp
Jhl42zGgjv3kO3SisLTaCBe6ZFmCfUoCXamPNMolqX4yaKIyYPfKlU5/1BPcHuxG6KqFGefaFSuy
VRwU1QNfnwi/zNUuo8syxxVujBquXC9sPF3oFWq2DVJkexx1P3GB1Flpe+rfr+uGdIXYiTVpIww7
SjfbVj+d/teHlzinLXPJhtgqVt2SrkMil2zlLbDY7Zd404stBDpSc6Wg8DB83DpS8Mm+Kw3qpx/K
+BbyI9wXpozjTTC+nY9pI9nPEhe+v9jwKeHLiEblY7dhH/pQNiQbsyMW4Vb+jQqjzyvUZQd4bR0s
14kYYHX4/mgjr3Zf5CPPm52ZPEHhyW7FPSkKlcZbOGOzMToNbmrPrafhM42Ju3vHsiBMMVBlB7sX
PxJ8YrdY+TTCs3rXVnXp+hUf3zYWPInmT62h4Mz/rwpb1c67pZQCGNfPgdLYIiZNGd9VrOwvfigX
jM6Bn5+VmK0VkeigKAXrLgxo1bZJn4RNXodAQh+0g4ynKPemz4oy6Kve/TPBjx+R0AlV0Ljdoyh2
LS1gLqeihXqDDUQzIAM65qDZx2szWJcw+TMOgnr/0Uc3IEZzsVor2lWEsF61yj8VWhZyWBv2KW+W
K/b6364CKVu3frkJW0XzRkNpcSWfSSFytEQPyIUjAGKbCDe8Qum+j27nK2xZ5Nv6chEPuBngZwfq
dDa8V5DfAltQWTsVEGdNtIQgVtg9Er8EdGVQmdJc8uN+NK+iZaeg00X+YPtLM8yZN+ekixOPPScB
QlXHhqIE3Ud8lDM9cbniO8JWKJCc6dxfjwZJYDhyv8lR0XOd+9+1mmd9kZdOQpnH0h+8PZiyzl5V
IaICuyRJpGkQ08xUb9kE+O0blpo6L2SIRAS7u+zqqrjvrRMcKF/xT474d8fekLUQxvXo9Cr+4D0G
BP1Cetnv7qNIJsEWjW8IBzJ+Dk3YRDlIoB75vz03axLdNNgB1MSzmAQFR++FM0t8ujhCsfqgyHba
TSixxKjMm7e0U7HGLrqooizMih3UMbYwDlRRdFGRwQ6I/q/Eyeh+GPEzR4OFUpO7d3rM5SpQAFT8
aw9Lj2Cokn3lwRUXTgP3YLCWDCHdEuotlxeCg4t0oCdf1NaT7n6W+Ajj40Dfdya1zXHl8JEG2Fco
pZ2/xlmrdsEonUSg21czI9RKzvoVucu6Zsz7wVGLkPcGJ6WffDefDjPWd2bRk4uAnU2I+UcNSsek
SAN5G9mEc1h8dJt6CpTbgqzrg+gHlVvsoJNi5XMPFO58NS4evavsVwhO86V/F8Wp1vMlh3ec5C4O
p/GlZkXbZOfjbHZ8IESFK3GNmD+hw+0d3Vs8uRopYNJxPPE6pYHfd1SZVTeQEnXJ5O4vEtlDn8Dc
vjigWWiJuGVCzROn/EWew66xzKHq+gCCbvjDXVBf97/f8DpXt3chhBmALCzbx1czbytnasAZkf9g
c4XYI2wdthvmvkId/wjJ1eOZKQllbb8hNAIQxOLicQp9q3w0j63TISOrS59JZfdhZqMBI5+kxNaz
FOm4ZN0Yns2mpvaKnTxT99SmXOSJcIAIxWQrFcyH4veBR/R+KVsSYpV+VJdSsgrG9rHmqdAEtz/f
pgR9o93AOsjsdKgSa09kdwTveJMK5JF6G5iM01MnKssPF3AqnBgmMZLSiCmD/sPooY7wpWNjccFy
7eLsaOfmDh9HeucUqeejboT7RBb/jvlwQbgXdiiGqoIVmo43ESsK+ffb9/p8tNb0xfZjCGGBr9BU
itwn3XTrtG7ez43BUxxJKmciYjIhXuCz1+r327aBPhUKl9YAeOI5Gv2vfhEV5gSv95/62E6S52Oc
K0t9hUpkjYQFVwo8l2R7muWR/fQKizMQF4SXmWsqJqtebf5yD7H9LBSk9BsA6uiDc7Ud8CY9VtMa
swSLjaiEBUQaqm5fv2F4NO+E70a1JLTLuEFzAkqM5XK2YahAihNSth+cWRj9at3ZSvSJGz1kTps+
Yh7teaYZLQiKrVzZRwTAPC6eBFhsbErOhTUVRr0iLEo1pib8Dr8dNUal3OWoCcH7QoH/hcd28r7S
Vl0GMmu8ZgWyhX/yKjG2Yrq3qYldZX3oUZo9y9CVPA0QdHfp+dMzmMLHFzwmx5n3Du5ZCP02gXoU
pZ0b8hXUrZOOjxH5JwSkSjeErSwPyaEPogoVXsShVfK0zfJBm8EBc9OJlBZE3EcQlgA7mLD/AkTF
JLrWEA+PlF1ZYEHZoq2uwf0L63WMICCkXX7qj38cdOfEX1EfurpyH1jLv5OYkZPUkgmZDtbZ+pOP
O+ki5Fn5N7DxWHZX+8eCRrRa6s8Zh5nTerGfYXZRK5ydFhJM47WiQjMnayfZp7ve0KwMedd+uYdZ
IleJDLvwCdQn0kiOmqrwjXEVYy9TxTkyucBpP68tf8ep9QqEpdFTJ3/gMGkSCkjIm1ZefPpsH70n
kKZXqr3OXL4BFDBsawPk9eL/2SG7EXy0u1bDOa4Hb+LoSDOdQUb2kQE4kJC7voDWoUSYrLDNI36E
YVjY4HT2SgZ8Io8/qWXl97pLNRbMRF7FrpBqySwCzHWOJ1DiCExwtrpkXBCQnvrcO+lttUsvyNGD
CLvNQn5dxZGo/zTyGOhn6MMXryMr89UmKe3LWRvnDzvd9iLqlgZHnsisdJJI+Fwm46aHdVLljM1C
/qbUJeKTm4h8aBbuBxnbmLju46MSsgHedwGbk0K0N8993Ai8KwScsaliqxMm3VjsA0Cd4YonTK1s
oIzOXpDG510WhxDIRYkqaMGrEG79ZODtS9J9OyUAl+T4wfWLk8OUSFUeFdyAnq1HtPA9MtfBthWd
oT+MYCtO0cXDdo7JHAFkWQdJ9UpPeelWmFCC1Ot2FLpAf+edF11Rcks/TBPWU6G5S/jAHRTgv3n1
y566O31mep47oVZlQEH52STnHkTMqRubIlR1eOYVg1PBCo4SADSBmbGTXTptZ8E0cs+pWzyceru4
VMqw+BvKhAo07V5PfK5prdN5fMtWGVXs8b3sGUam3FJY4yUWHaD/CX09UlZ8vdXgVHaeKYe8j41T
jpKXabOVshPOcQ40lRwuR5WfqLe9JvKKJmU/31kR70+rEE2vjMoeCTav27kRMpFCn4aTBkwHYDLQ
7bsAFJRvEOWvSnRB13Dob8gbBiN/R/zwou8SHYzzEbXHul9wBZL08YCgJMQRYyB/klsKSz61J6NE
sSMjl4Hmh3NDMMZGQPz68ng7yWc4gpgisvWl/OTar88ptcMlkWuUTslsHblHvV7Gm26Sjmnh9rRu
LW2CcQn+LCk8y5Un2Xpjp9bNTLKp0NwwSFgvf3/huWS/WEXYdauuMUOy7ZUqKWSdKSd+WZ8FAvZi
vrKQy6py8kPBghc11YDh99JrEuDMXhyZ3hpYXBy9RtL8aOtbZs4UGagXMkUulv80H7pl7H2DNk4Z
cqNZFDVipUEbsEHD7tEVmVjg/EeKovZLWZcLKSvQv7qsGDz2igttTSCKXuapSWM0io3m0mgbaTec
cmyX4pKQwrdrwhprtd5D3hZJtPT2RVSc1ugVEhRMD7/pCNY4StNSf1U26bgVZFCJKlWBOux/N7fE
GItv2UOifZhm7pg4HwE2oXzxIim3x46W4YgJFjfhOIGq6pKBrmk988eOsCy4h2+RNRBw1Fri4T2R
pyTpp/cloTUC53k0/m2gQpUfb8FiLLqtUYhEIFq+u3RuJxrryviJFr+GdfmH0VXsQ8M71uJ253Sb
LqOETOAOZL/75hRzw+npG2AwPsT7t7xOPXI646w04q5A81nJcEWrGr3J4vwRhN/2ezygYA1YHuWK
qzSAh5ImXlvY1rS/0kjCJE39XLmGtK6PTDRHl3+Ow4HJvvcEUwKypZy0NF+plBqeQ5Sk/o86rYs6
lRD2ibYU6tlFl7PoDb7cFuIR8LPqsKD7Z/vPfFVnHzYuUVyoKq1HpkmM1NqJgmrXMV7odx78qCsF
F/75IX+SyQvWfqlb/R3fBHzLMwOjjxtI8VRlfXp4TemAJSfA9uZ6Ms5i2H0KT4u75jhOphTkMJLN
BSqtSTJJ2wLG5+yYe+RYd0OcV84VElUm0MnRGLbPQ2ulOwycdpbgmhO97Hh1u34vfSkO/o05zRro
PnfMdErhUDaLsJagL5+3a8O1/Cyf0o147IbEpvlnHztnhlSfXc22p1XwLP7S5FuE/qZoWvDap5x+
foeFJpJszT9zWqOEMJhWWDFzNzMLK1I+PGhYSYKSU0TCLr6RwnTE1WkLo0fx8mTc/EMq65KpzAfg
V+C2D7nK4oF0O0n2sXhKZajfFd6QKxwdekTvBNnvpDruKEZHo77ZJQbUkgPUJ74Pd8QHGKEvSD4G
+gIiLNa5+LaA9esAfCAsW7++1d62ofz6OJoWOkXZe7V0hx0ONC22hw9nme+vz/kKP5JX08Whrzmy
apId6eyfEoTLHPi6puwcoXMTcMpt12i7671UmNdHNxF2twVi+Xp9FMmjvOjtJguonw5U1UguBBVn
ARsZNSnwKmm15bECnaexBx9LxNBK0xxuO4g7qTCkrxuAB3ZQ8XbaiRp2AkD5DjOQG2vNgKFS8gXE
1pSELwNVRhjTMiRAC9qOnh8D7/DnXhWH91MC32PPO1gYeLCBUmGqxkdILtS4GYk8YX/8qsQUiuiC
hiO6AzxEkwrvGRr8GPsGNwttu9dt+E3rI2MlVXsM/+Bj9cNWvgJ2unmrOVIIi3q6M83iE4VtI+hg
vAU2rDmasGj0ConIdnPzF8gTvxMGUs5SMHqBhVuO+T8i3fzHlAgtp7eSAsW+TAk3cNJqD4mDw6Gy
PKCrUYxDKcncpxzwsrnWFgxK7AMZUk8kQ2ozvU01qY5DrGUrV0nwvOfokL7Kb5VzRmAsWzp6xF3L
Q42rPMLtHIkCf02NpxXeFYRLqY4WaERWt23hyqpg+ohz68RyKLSxK2oMcS0zLCqFYgTgCUuR4FHA
6ewWWZJ0lSnIpLx8dd0mqzkF3Ptp7RIx25rHB4K+A3Agi8bXU+m3Kh1mbiXDTYvOIy8s+fXdb7ap
O8OIGP5OzSJ0ZMsvmmvQrDYe80LwKSHn+bnyitb6Nhq07kt7AvR9g+Q2G/+/gl4RC4VIF7ANB7T7
QNV0O3OC0Rr2Wc5tPLrIZiZ/eUWgAvfyT11nyGYxBKHuinVYiC3PAuoFitGlcU5pD2s7zKSKJT/H
FwUUe1yzEZgnX/nRZ4Pvk8TYRhjp7qFx6CqoMXDwz4XmYbvk0MV2uF+yqT4H0Z8K3kWq9BDwkrlf
YJqchv4ptymNKZO+pbRTuKkJzVO3j37nfee2OFcCBssa1SFcKo3O2hf5tXycwKS38AUCREiWT0aw
bZ1wLQF7nIMYebEW3I4tG0lbbgUjLNcGhfEHt6ZhZEhkUvHkK0K1ArwO3ndkAiAM432yXQhwvd4d
xrBehtVuC+XL25oM6nAsRvMkQ5+2OcFExQk2R6QV5hX26B4S4fIMfLluq6+BFql6cwOTqRUzLPg2
2xn7T9lhDj9U2i6sh6ZmaivsZ77OgVtYd78h+Lmuj6tKr4vLldk1aIULW+sz+36I8cyVwfBuh2tH
NTK+ZYS0inzyWgbE45EzAwoH55N3tT6jq+vTzzcndKE4JSfSU9GMcrXRbq+KdBPn0P0xfd9EYsS1
ekrJdwrYubBp4Juv9WHxn+MO6jTT+PwXw223vGmn/ep28T1ot/lU0d6g8pxUN+qqL1gR4ECrorx2
6+fs2n7W4Dk5Igtu3nCbLN+bbB+KuXQa+E88oEAQzSG6jjEyR92QNuaXulImmFY+aLeeM3Nkdgal
O/kX2sSm0u3zGvZGi4FgXgAWTDff+10v4P0PHW0MLCR/ZKEss6l3kIFubN0K73P3XXZjR5YTbP0W
PPiTVeCGdI5PLlwjx53vsAcGkLzQ1aiz+85le0+W+00zQDQemTJ0Ra2zMfSsjd/a6DYaqOQ8197T
JNOAA4urlDVuU6k3edFtGF5e2OS9CTA4pFGyVD0CANxr79PGsoAg9ZInLl2sEtnj6c7WbBu0uFpu
70DcSMcc52Ewgn14SV36r/T4l0mesvkxcx/FPsfbkGwneQdANs3i+nuKCfAAeXObZCIVpSAIcN15
ipJse7Sf7khakj0kxF/RTfcRnqkPs4k1NM6DfSNu9jWMkKFoyPohnxxUlxKryvCoBg5OmVi0/mK4
If3s5YyBiFBXSvXblz06W6LTvZi8G10I3zVdxBmPPXPQ1M1xpiLC7eomWjYyUgctHjSwl1+JRhlI
12TRiZWHrl7mO6tXhdWVU6BNclf9SkOuWoZc+IusvAkMR0jyXqG6OJLst0iKmCJo1+tNV3CxSubw
gvozYdp5sMpo+rbY+xwkmiU3oCl1QBz587VnZqbL4l3MmriWi6drIGuec4hnsKpFyuaRGXBJiZGm
xFytaem+jDlsSVvTqw3/FpYAPYVq1Gz2wYtJgx0+x3hnOpyLH3tKgplD0wZnKxiANFQW2nWgxpIf
m76GTqevDx5RwbS9qGfv4CvEQXkOP0u4ipWjY5wLFxxNwIHchZssn9zwE3TnKjT0+Khdq1/f9+K5
thVLXf836k6DLaZJu4FiTxlCYm2f5gWrVEiu2O2t1UyVTlmDOPgFPyAGBxjZ+JWZk11EqPpF44hN
d8TQTKYAz733l5IXN2Whi6XeVdFrEbTsj1m7kAU+Y8pzQaEr8+3MJIzC68K0SYSoX9saiAtHO55o
zPwxclxrkldtASlgU6UJ6GKI2n7gck42WP4vVdZ3evL9EK13atOyi8sMnUDvsWJ1S8+I23PbBJi4
UsNeA9OlQGt64bc4NSOP8wDgb8f8AftDSYTL+yWGYH02joe766d1hA4Z86FM9Rgzhq4QJ05i0PVc
ukhAAZ/teuc7pqSNyuZ9ju2N1wvDs5i/Sq8HxEGJPQYRNh9omqdfYWCgCjrgzklmgAhngm5gg075
w1LvA+IqeE3McRAAFC7naxWQfhhdSMWSxPgZkMyUCMj3PiEyETfsuUV6TiyE0fAwIwD6LlY2OLYx
3h6dQRmfG8xsp5by6fmhsVQYX3+du3Ck77tweEBcE3H2X0NM2Og5kDqDd6BSOlVucminZtxtzq/q
tHGGF0Bh42ks74Vsil2f85QFi7fU6k5mnOW+/Xi0ShsyAV2TItH0E5hd8MIPJc/7zAMAxN58cACR
MJKEcjovspx5UfdELCjHrpzsonm94M2hy7C2XDGujuP20q9eKZ3mA1us8knrcHZ8/wqOPH6ha4Ya
4jaOceQ7rY/KDdDZbolzajGq5XGfpFouclNh/xwgxPcA0xNQyDzyIMAWARnWXxMwxE/OJxchnqeR
0Dyy9uMb4OTvJ72JnXbcpVjO7w1R8D9Q6UJ8WAYVKUtnWes2QkM+oNqn+5M2gcljr4WOom3k0U9w
nayzKnw6FCmyNeeDV4ffu8oo+vjL9DdsSOd66yjT4N0LEg/fVjbQ75NLzJx8CJeAc0B3E9FRjO/9
GCc7l1gZJtBD+LTUcS5hoZmeLKMeGmbWYB8ejFMtzdymvQV04q/W9VuLJdjWTqpDBAELW7RwtxJs
Im86Ag52yQRAlvqX3R+aU7NaDwLgmB6xaukzfUVQX3+oVxpyV1w4KGbQyX7fjtd793Hrnjk16LpP
wJaz6zTJlgQC8gTwW/KnXumoHKxmyzfity3HlF1MoGXOyZkOiV/jN1t65JYhCSg+BchUMJFmjrjg
E+eawMZW6KI8jkcHb1dnTPQWYbJKFnMzrmjzCmdNRD9JEj5E/GMpvI9mm90Eo1Nu3t2gGIURKT4o
2U0zPL4upGXZlHvqc7IiEdr7bWix0XC6tKJjCDDyJsDmtE3YQtffOOVZUjGOvQP6zA1Ies/y2m5k
OAURSkdGF1KAs+KdNwapDClA7wAS2K9w/F/Sf/yZ6s+UG6CgxGM9lX2BT5swb/x3bZcjD+wFJfqI
nj8UaiCOM65IKbcl8wVACISPSjhLoQ7BE7mdJ/UlNZ9hjpbQR0VLP3xx2yVOJ0R+iyo/GLg6ikmG
iaBy0fxxhCnaOoKvLCftXBab7+9VvBoN5ydpbqKQMdc1CZ6RFBmkIbQvLTsiVGt2U09aQJuEI5vc
LrDWq4Ss8n+1uTqFwrJYZg/NkuLPa0vGv6Ws1tfMV4n/WKqW7Va3P9uEYWr5oSPjAaWBptdcetef
kN4//pMmxDu4QqUC8S4UH5O3/Sg3Z+Tw+IyuOoBSKbIRagI8abVnPeD/pgvpkqDsZaNBqPIE+WsM
escAzeLseR5VQMLsz427+zvUriIctpGZHoz6AeU+LPrhSjVlm8f1qzwFVa2XEwA5yimfMFVBj99c
oybe1fP60LvbSHtHFuy3kAgqKbXVsaTTFPpowAlpJABucjS/KglDMTyt8O9/ViT2wyXxwfHaXMju
08+rBQaAUnGWH2/aOQN7nO2LaifeAWXzxLAObVEUGNd7nZrYxTa8zX/wRYnEE1U/ZDQVw980wGTH
RgaW11UuMNjaq7b+2m9Msrzd/bx1JUdc5gz/6pBbBdYcLqUIQab2frAtO8zI47pZLWZ1W+izCB3b
5+8bDwR2LggvlliUAZQ+DEBdebneBwge3tyoTwLmukuPTdsFvy5nUzy8v4u4k/8iVYi1aZ1c0D+h
GqIq4+e4tXvnFk6V4jGVbPCGnEXkMoKt+hPFLPvxl1Hw4JFtB7dvPXpagtz7ZLdFtIVxWriyqnfK
5jc70u/wzcrTDkR7pDyN4iq4qHVl7HGOFAdcpckYmkq1Mj/zeVfSjNgUToTCUp8i05ot1eWR3EXe
jAsfsVw/aoR8CQ7ZQYQjCspUphabD0xL9j6YAMdJyTbOoWQWsUhhwF3AjtM6qNgJQD/IpDc5VZoI
ByTRx563upBf0Wl6pbe8ebpQXnZbSeiN6w6KFfrWeVSC8And7Z1wKLBJU/VOme9a18hgfHfVpa54
zHVPAZZuQfqliL5kcQLZGb2c+nOlbEOLQvYsWVu6L9JZtG8E9nM8WLv7p1g+kl8T6nwefAv6+vPT
WpRHm9cSh7x1srg9l2C1Otr0CE6jVEBaChWQZHDnTBsKRzn6RdBQ/nu7fXmYOEww2c1zS+DfDt2D
YvyM4Clw/rKFvZX24XboI4Rv9eflBdMxVPa2hX0z2XAYode2nFdHuVL2L61H+wS5ypuekAoqsraR
BL6eSG5dq/BbFSYZLPIk35PXl9E94eo/cZLCIPk0wDjYbIwvrGGQoqvB8uSmI1ADNdMGS55tKUHc
ShdcwRj19hO9UVeCGqervnFF1HS5/iJUY/zZXcBvtl29DLG/i1199BbYX3rnlk3Wcxl1i1ZIKZnG
bBhRXxyq8eeWTsQtgbsFof/VO2/5QvILZ4eAHHawHGxTH0TL3y4c+162pIeSJljegQYOoNJ2XSwH
dqseDbxwV/hNIzR4PUnBU6GTW3pW9Ct+Jv7TgpIHIWetHipLVfx09bUzY2OpAiPEjbfhrxbckwHF
BvIFyZCjne+ojBBlvlRbCy4GI10w/Lnr04XLzBwxa5Ms9oB9rZf2Y2KPcqkhmLXg2kwI6aLxyfDL
ge+OkmZ3mPwXgWbuo8ravDsuHEdD7eYp+5t6XAuouP82qOLMuEpGa0aGAJ9QgNRUD8jPxjlyOf4n
eS7KEwJ+TPlQBMuBZ5aFm2umeCL1iO9lqv3UD+rlUFdVEEmqLRikEKIT9OpslzdVC8S/ZfECl/u6
Bc8GBVi9qRqzrGzHg2D2xThQgDbIta9tRlKTTCIwd/niC8I0uVof74BIUVST0JRvWLdfNj39rU3E
3GYkfFpEkn+zc9tdv0GZVIpFQhnxncSURQNPNSgbNHycohhGiyrOQBpDlUDfD/K+fFCGX2r/rbck
zFrE4n4CZAFK8C7wqClp0lPVjiMh7FUBim/2OSRkYm+ekfaO24H5YhiQ5Gubji8hxG3AqwvUZvUd
P9IdoQOlQGd3QH+nWYI23il4MddFqYeBxfhjLTPQ+BRCSXA5yQ1bX65gxkSpSF6kJH75dlEpSyU5
5r9x8g5hc/sIKfRAoJfUbKBdxiJ4nClvfTC1tVVLpbefzeNgkrMHfSgJJpqRJi4/fll6FWEZXxkF
o/TD4VQ9qWODy+ePE0RgGagzfGLAya4WHnhbU6z0iZVOv0VALxrkk9ihprDzBL63fV+cJ1crXfnW
Kt8KBS/puh2einC1jAFO5ABvnxee3g+FAQT3+E8Yifl9VFnFPhXdImTQA9IfZuh4UF1urS4dFjoQ
WDOUfY1RlaX+JmwyCcpCQmFAYxuWsnHy73sw9UvdQb+4O4SGcoq4wB72KdnLRL/SiEyU3r6HRwgY
e8PM+5F8xn4FcXh3I3hxbtpaGHBKXyUFDGbzXqVEhXK8eyqgkxilvbXTyiVO8w8XTLKCq0tY6xZq
CLwjUQY3AQrYUWj6nsK1kuNjoMEiGv+PFE/irDCSOY+OT5oSPt3Nn5cO09q/jcLFai3lcweYQ4Fb
PAydHukhRaE42vf1OY7weT8O3rd9meFeO1soS+90ZqacGCitnq/s74KZ3+qCSn2Dih++IqYKrtzc
9CPjywZyzcwrd8n0LAbS7Nl4hpWQrlXqsHUA0S5e5PumVxcNpvkaS12znyDWAwXlfVbp1IuYEz39
4OSkqOMt7IF6iEUqQa/L64ApMJlPj3sZP+4/vRvUEGYMOEe/pWnMxe6gs1YiYyOcysQXkA2JzrmH
trzSj8yheQA5MyQWC928Stwy4mG8FoHLdP0xL6Fxhx8hCQFzfT14BzIc602bGXj/kWEpIl7fODMo
N8La5Dvsg3akpRmWhWKQjZHY1cSz7bOr+KERuhwH4pa5dlMVdtYwg8tkIsDI2UlarS6EyGYnvA6B
XFNye2HZ1hCnQKEKgMo74l13gYOMi0yw787lTjANnjcCsxw70ws2gvuweDMotBAKMUt2YOdEjpQo
hotgvWZRFvvbWj+6GzoJW92cJ6eYVeqRzsFoK+4ammO7z4D5bpBKw9+6lzA1wmde56c/yTkleh63
7+pwL/1hmdhxGhA1PJRRr9tAGEfD3UETwRmxe4NR2gX8SECrKRLUIey8pOCUK1fy8UrFBLIhM754
RHGP0i3fg8D1vQGypjEYMSCdoo9Su7NZ/dDjEAjn1NkryRioYoZYNe2cGnRB1m2ksmqyaKQfQZG2
hfPkqoqotLKy8L5jtUq2I10OJheVP71g3OydBzURNveOFzg8AFPQrnfRyjww1BEdtycNYtCBBMVO
tZjbkAls85uIoP/kEQaW20EPziqr/YbF9phIj0eAENa/3SG2VnM7Dq++KswgagltCW3N63UAug7S
2V75sJDxdQe7/EcQ5vj+auJ9l61MPtkjVntqR0qOPJUERtW3O7/e7+8Quvo1FbC+394BEyIW8iMC
bC+f51ZnS7gpDpilDyALkMZMvTDo40QmFN5j9qXvoyBRT7h5moO8XSt89IhHx7CEdThbfvg83fnt
c0giWd1L0v2ZlFKSnx4ihLS0cTPSmNtRslS+8B97F05Srczn23FouLuEbPfjPzzPoc7qV2E4ro8U
/XLlGNuTVqVx7Vj3QXaEOgSVLCupL1J7lqYMQHdvky8eRoTuU4DGXTKy+9zjFdtp6fifalBstLe0
+P5G1gFHYnygQhqQ9LGeEShBnHWFW4uN1xEt7dMPsfc/lzRkSIqaAcPDvP5OX8yh4Wb7Yh3mn/uV
/TlzSgkMWKJzfu4EVN5bpCWbwtcc23d4+5mUy3dE5fdXXdgl6JTSIm7KcroNIjZwg8b5K38ChXLz
qbSEfUkH11Q1A21tH02Bqa5s1Yd0rLb2LsUf2pzTOkvbWHFzIJVxzMZwpGvez30oM/sGSD/CUu0d
qf8BDcQHDVYCXEUL/f7MvTX4G5xF1zQ+/0c6RMXKtPOxA2PFEeZHXzYL4JJmCTzCO3gsUJe4SLXa
crDzWuVZj4gGfFYAAfGZvflhIUMmYhPcitMOqrwMGGNQIpwT7EwdvJCBZ48yJ7Zrhzje+/8Yzzy3
MQJRsWX1SwvliGgHPv/DqPh9r3I8Q4Ps1yzvSCE6wMRie+9PSLl8cdU2TU9U6JcbHPt51NQv+qRR
WTEjaXmv/ZlPJwgJDUjGpDSOhinJCU90Ba+XD6SqrCrDtJf06k38LW7gbH53ELiG+yAKlAyLl7U+
8/i45T0Z467qiNlO1msIPPDBM7MhG1TZdUqfQarhXACDnBplb5YP7NabgWVL1XyTDJc4dUAWY3V8
i1e8An+Dad+5EtShmDazkdds+3xEN1yv6vWRuEsqD9Pc7omQjaVFiBgyaycLpc4/pU2FFmHRU8po
mDM0H0BPqyB4u2iHIJLlXZXdihG9DTjDq+KcSbK3gxOU36WweMz6MZvxym2CfSrYjp0mQdx9MpVl
4oHs+O+2mTB5LsjD8yUHorx1QYLTHW6DqeAmm86Is18cklNSFLUtHDOjcYEy2G9uPKsr/tKPwyel
PUF/eLXd/Zayzz/dU4CMauLKh1RsZvMCVy/XGc/Gjr1+APcP74LgiiM/Qbxwt0JefC7LdLDsgQ02
vZlzGU7AuZ5Mcd/8iHg4DAD0yZ+kXnMO//yHnUmgjxMct3+MLCRuKjMOF9sZZaUjra0x0wNbyRaf
mAu1MAgVlqomv85uoF2rcZya7FMgZ4capxuQvU55iY3Di92T58rlIhWBIGks/+fp88cWanVlVFtW
CQR0fjjjdi/9YAOtIkyCs4SAKoXFixFxNB0TeVF/PP4T4l5ww6llcpApUaKjNyXnZhi53XSUCtoB
6lYhjb93uFalqRTob0sNC9mKvVJmf22jjJyjT4ZNKOCd99o+cpsgf6hV0dgoMNMwj1bXuviO1ZXL
H/8lLfBX03kul63tdNTEoD/DPn5bLcNcvh0gm/o5c+s14oA4GVg8P3afy+cfMho6Ye2ACDXvgggD
xIPVykfIOCKZFkSdOyRTN4EH9zQ+r/Zt926WRdZ2QSTs9eHI5Q4pC14zLO5XETZ+IWzh0xHtUAOq
PRh6QYhSUKQQP/kVOkzBAewQRE0v4ucCApDHt/hEiPK3QNeZA7qBHmrxwlugf1KHqcEBg0iktCFj
WxpPsL9EmNJe7gedr5im94pI6u07pBRvBknjFH7t1jDZrW022LEFHZlc7MBtVa1Mp7v3nVJNdn6i
hnFlYym7vB4fEx5fyCLY+TtjvNteVpXZbQZ9c32Oeu62AGwNIUI4PU4KZRoModk5dRebUtmmg8Qd
6nwoF8/aa+H+oPDbUt15EFrjEXoZpxed4AkipJwZgFMoWlEW0qpSWVKZ98l7lsuV4Ek5xlzDRtny
XpMWc7UpECYYXfTR/IYWjLhNspMATGjb4qCKPHWda8taYDkDTXwUaqweq6/Lgkc8Yep4AJNiPuci
R9zGFcCSfj2ZMpYaysVEjrp3M4Hb0COZ12lkSjUYVu01q7L6tEisjaO9MpRyzX+J/jHszoct+QLe
DzFjaHKHylDJA8liG1R9/MfrFQ25kJ0kZ5bp9asL20lAqRFv0VgjBIlnfTO3eW2H1tjNrPmjvbML
DQGVaGjnBTTZC6q4f7Q6Wr3Tn0VBP87V57xCj5id9y53yHNZHpd8GE9bR9gKgVwZwYdKeYsTJhLw
c0E6F4VPp4PTG73H1L4te1h4O8yZH21/EdxfpWOcr0djIH0beh8guG1p9ZhvJFUtu55uYnUnrFbL
CzHb3gTJcy+lpxbtItaxuxL/8u5NSVhC1vblfsc+xlCNR6OCFG56gahXY/bFdB06m6lwYAhLkcWf
Zchqf/XYcYVXwwWknht5o04MMOMiAwKAPIQdERC0eBpWXMxHGJk2Ib+xmblgNmVjpwPj+chSgN8Y
+aHTWaLppPWvH6G2jvQJDUWMGrh08HP0GybSdgr64LOWx8HclaWQo16EVccsXalpHo17nd48U4oE
ie0TCoUaT5kApBXEyR9BbG4JyIIfoJMrk+HQ63WO6DKAy7oQWKkU/XNq3Ejw7HCtOVumTJUdxAaI
lRzNhs9r2huwGScF/BjiHNpfFglPN86orEHS9ce0rZpW6oo74tFD6axgqm52X7MVr/HByMtaTNoH
NqPqIKvC4R4rF3IWNfpj3kYCVfPf0+gFXdR0Q0gyK8VYLmWaFNLzRDJfkLUg9gA7nQwot2FijNfK
98wMgYlHR3MJhTtnLB1w4ZISKfydidr5dF57VedRcxMIkeet79ojiQN7zM7kko8VCjdwafop/6tR
FlbG9S2FyabIEwkY6fhgyM2YZc8/JBcEJFH+rm/p/OTGab8SRUCt1WjXG+KOWSE1/Iso6qu0yIFI
/NqxUylCZ/DknzCYZKH+QelJnVbGws/IkUUt+FP3lYWv67x/a8R6ZTtsdz1j+fpRSqu+dceIpnbS
Ebv7FD7qPcmA6q6kV3sij8/gOYCbsej0GZHJEw1OPdcY2C9Ka35T/c5qo0uvqRvErnMBWvbfaOlG
5omRl9CtX0Bw5DLv9YQd58gHPM+0Nh4KyPLpcuIvxfU/z+Q8YNottGl7uNyuxOz1zp5VNJ8cYEWz
I4rDFzIA85mVRKw18kGGJXtyF4H0Q9hlzYIQUZP0DPAapo28WCufv+O6RDjmN/wPeU4Xt6Pkc1WQ
rATnr5rYdkZG+yKfr5dpLFkoGCniFLECbdEG+ejIRGcuTSCyMu7yK++7OdGjSCrciDxLOi/pWSKj
F5qdSlIWrOYTKjQsCByuw3I02dN6ndjJSZaV5gq7Ayk9iUU1ziUFnimo925ZYhmuOgkFvTB+avZe
2lfh2fvKRXvqwtiV7ciF/pa7TGjpD3eB3kgLKqaZ2yswQZcGniYTy7Ww7+xAgDcPXiKSelIM2nGA
vzWWO/gsbxYfQR40hkHC/1X0IiVYNMKpBI7btNoRxix1HczcCVu807pNxOlIPwFTsax0jm9ZX4Rg
6mOb2FoWr4Ixz1S1QaohZF0rV6bk2L4XJ6R/lIj8fkgKOMBiO2lhcUFs3mvW8iwkwdcUkIjsFikz
lfDuMu/sjbUjPHv+4s3CdGOxHcBnIdBcBAskRX8/GUvrGKWwkk0k1Q5hlJqkJczN8DRJku25S3Xa
ByP5PJk1IqEU6ramOkKfBOwNhav26hG1gvaH7Z/O6tC3OEWJZOjiHbGtDpgsR6ZkCnUiR+TqKiTd
jJuKAYyBqv8HmKoj4DMffRV7Cgm2d4xt4idpJNUig8t/7zhKanQRr7aUBQBX7X4uD7qovV/dMRgP
9fjGLqqQqZvFXRqETjqasu9YlFTralxGTOX7DyiUD6hMjHGQosLdlqrzCjEXfn8UtmbexSYTae7f
uW5SFDb1uaOaq1RMF/ZrOR42ch5HVMRV+dT58/FlkIUa5RUiLE9Qq8PZT7LABiGWH31nN6C8RKDD
xzWeC6/XZC9+FnpAXsYOX91rBckp9GCcAcJ6+100m9RQFYzCDEOQFDTjKWokxFTiLcehEQSf0kaP
On2EI3urIsAP4jb8Px+lzHIVZ/eQz4ZdICEYRS50cfHfXgcY9eira0nhMw4I1qu5nkNDk0NlwPr6
57f/sWoesiSEPje3At9fKIS3bkOFt6iNfEuCQRo/duPJabHF8l4xQiAykRZfsSmUlV3KXKbdYHIE
rkDwr7dKFFl9x/EP2aX/VLtruEFLbnR7yjjHOnIypGeOxA2xKApxbWPQBsRCgRZnl7sJbetU42E9
/ZGj4AHt+4sPJ1FRwRHUWKDj42O0vfqWPx0MnavmKOzwldh1k1n2/9cmfSTYJjK+NMsNYXbXQcEO
lcUtCdSEyjD3EvFX6lCovk8Ic5SuQUchcU7Z9o0kJmiCvTRRQq0x7uBvTFeBS5xnwiKDhAplHrqM
i0huyXRYxDl3alGPLAswGQBe/7kRMaYcP2F6AErW5Q8LN6HQ7X2HLH+zyuzpoOR08VjRcnToDZ3p
vat6HsrVKVdgzOj3JvGzgbWBUvoxukLa8dbbXzjZxDEzd7DvxvLvH7tQu7SuVxPcm8XJQZi6wwRr
eAO4rgEHJJRiFmrqQnJ6uMWMXNJ46pNV+RNoQwvOvverYSGpB+Aqc327wB2oFeA7COE5Ej6kXmLO
rYI/154g3dozCzF9QsZUCw/ku4TDMB5vTBuPWkd1RoOQkfN+6gBOS6ls/zaCQB4nLND1VF+po9rv
avHpvSGHKklaKczxGekC23nA52fkny94LckUMdPIIF4XYOsHDXf1tahaI6H7l48GyOTJJvfSkPuB
RvUYsHg1LIX28Po/XH1rZ8JGSsng/WkgFtQZPBOrZ2qNUnSTbIPwWu5pn8/j5iXzKYBjbbgJzbOn
AJqCrIrlGupJ+JTxhHfeiyaiH9vrRR7gGlEMj+PLeUNR3sZPEkPu9RQr6HCnDwBgKhnyYG9aLKTz
4AU8lhOJRPEH/1TUNCsL5qTfZP062o5KRXakmkIgQ2YpMjvbf2Nis+lwjzLIZPIHc+zNnxf3GMM9
bcJ5dQeMFiDj6WOop26Jz9Na9/6iCVEDc5vkXefuanPeZgUdzT7sDdzNXVR6smGz5RMDPPZJCO6V
C6Xo5KkAjZ4u9Koz5MaqyybKCGlW72k2kU5hujK3rjDCnTQTPe2VguQm1kHe2rbwDjIsLIsMGHuQ
qDDBZcQzfVyNfunbObSyF2hmcImid58zrgqUmikYtu/Py3LH5z/hVSOCcUDpBaLo9ZH3YKSbBAZn
LxLBT+2LPdKrxqeLjmqX3vQA7VUslQl4nCJ6aCRQQguVjS3nXZ6nD3FE0rAKBH3L1B9IkeXt0gQg
E28C+v0fp0CualRFYcBQydbpRxkFuLnkVunxfT0E6GEHchGSMXl6QYmSNnnBNkKGdCP0LQgRZvI/
4LHk8DHfyJs0cfZi1Gkyny9+zZjTOmESQQwaSpK3n2wGzV/DkI/vUq4jq/O/PNjNTpLj/13IoWyr
ZgiIi/X16tJJ4gql4GfDln+ujbo6FbvBuLauMc2asPRvS0V1EiIDpgPULrdfEAjegw/Xu+lyUYSR
Sg8Pl31ZW7rqW9hqhH9OPh2ZQEBlwqhWXzV/zyhfUDq/tWvvvIzu5fjml/gbrorgfxNi9yC1mBUG
j2i0kQG2ppOZnG7S6Fy+XFRQVE68yr858KXNKcIvLZuouRmQODeAJHNZjfugcR/+GSgLCEHoijq9
L+xLJReX43shmQ33rZRZq3mugf2bIus/bciKdouZLYXosYHkz+SpaCH03pLp6Vti3iaA/nfifQrF
anZWz8iw0rwj0vPq0js0Jqr3Ky+lk0EtyJe7epVv0rT1U7ugZPENqMRdc425p04ozoedV6/YG715
2BUDVWR8J2r0VjdX36fjS8uvuHO6i3opSyECWV+KHA4Fxjyh2R8CHqxeG2vml9qSevIiKHFXlLGS
Q/4gbsV75k+vFCj9otBworxStkM3LRTJju0pY3lYwwq9WMrjZW4pUi08rw3h7fEwQwxpn+IQiSXp
xzPODGfN9IE5v1vx7ayZHIMGYrnzElkXZ++nGiyx8odreoT3cYzwOFJqmf7V2w0/Qb0BwrPoGXNL
S4PX6y6xMc51ZcM+TblLCHqJw3q8v+8WVX/pgQvJEffJgWXEu0oEqQ5TUNMRnsuDxfCjkQCSVwhl
R6MYkNoBgTARurtVVYAAaxjQjHNfp77a/9MLu/Y0FY9qJmm7x8ZTLvIHT3fbmVTqv6epMPos8nH6
Axmp7NtA3QSPfeKMGUDMtObYNFi61Z5txdWp5CEQl94M2OoL2PpGjx/pdIZkBcc6UemQr+Vi6lpd
B04DUhPfkyUj45MFK5dOS3NL7f+NLtvVJCVpifrYBa3VsbK8tEc5hCCfGvEmPPytRPysLWowTLjh
DaHFyKUfc3QxUantf8FPQj233GJKABMzOMBQQB8q3Hxp+VPnTdwS17aF7UM4TaCvk3IGa8LXUfCe
Dopgi7u8jmH5b1OK+jwx74vlKOqc/A1gCiUioFN56nbPPzc9YuzFKgu7P/DY85d55VcusY7KL6jk
g86S001hV8tj6UpuQY6AomowoZdryYCZrf4bZRXqpioS4fwKUbRID6DDzGgiiJ3SfbTCzTdd5CGW
DsUzN5ALStiLJRyEwgfI7U/kTe/vf99QAk0nBszw6JYEcnbue+hVsaFG0WbGEOqvqsxh70EJjWVe
wVE2z5fy84zSskFsEQyL/rN1tz/w1HnUIaEC1mDoSf6AUJQEPtj60IQwDXbL29mcnAEqTFaLuhkn
ZLaEAgOhrqOw5BY1FHBO6pLJBwVsvM7+fwIf4NIdubkmIMxaIcLf6OSWHv83u6tVthgqKo2X+dRj
Z3+hU4LETBflVNK/Es3vwDQvBD/VqmYY3Eio20t105RLZoB+6CLhFTisUNavCANkOE5SUL7ZZpYd
hz5mIxgA7Aud7p4sv4nXE+WWMC2yDdYI7xHd3KxKQIBTogZ437Q3st400/YN6iwmIj8wBzsn512u
MX4BFU4ltoA8RmWiuLuy5KLaHNouXr/tmbWIHjQgsrILqgWvndr8RkimfZ13hPRC25ohNLLaKfSB
6S5tnunU3p0XxO5PvLp4hSA1kBmas4/GjeAFNnCnhwUGJqG2HfDuaig1YAX6x6tYq/7DsutQ5K6h
rp+qBhIkBgmcHzJOqbMW3rzOgkHRb1TqX2hS7ukY/dg3LqMtJtLRUJUfR9c9MrqNE9TZPGRWGLbU
goTaFspPrTCiL9FOn98mluLx6+Xf7oAkqwT53ESzkBEv6Zc6EK5hfwB4CNtkruY4KvIoa4jyFU49
NlbhId3sVx8cD1kNxSR+POb/oH2zQagmM9ENUc8qwOfnaTuZ5lU1lUHfDpaVLtZ3gXgRzy/vuctm
QnLOWdch3pM3I5WiWR5jnJdJ3/AYMBAQYUQjcTohKna5jm7hxe+4SKuIJQMCMZqm5oqemUwMSn34
uugE1GZ18iJ45qOngQsEMDmQFYyYn59evSHNP41AISflALm0DreJtX2VuLBsHxYrImoP94xYaiRM
PL6PVbeLpoi7yxkDYts33I/SSzmCLFqnV9DkWi6zYnGgF2JtrrJxnrlTv2D9c7n/GUS8qaKPPN6G
DRctQ2M5weNks0gftJxoYtOSnq0pFOSfJfzu03mki1ohfXgnaGk7sLbyGIih7+3xYUqCojRHhkGc
uf34DVso/x8UVM+Xk+YpXL0J+l8ewij/KucMXCNe1Tak2raufmI+niRAIUGZTBOXC07NAky0WeWX
ZaK4XOruorIoz/VZ8F6mVxukL+BbUQZLOgtSNwYzJX+1ZuhjXnAGep3YN/Yg5TgYdtFMZA3su54U
a35y9O9dwXsGTsFIKwUAC0ARAFu8rTFvPOFtsyq+dHGs4sOSi30owPoRVX3eFrGUI/AOyQUBki+N
Tql1tIW37iXWQ1D38TWtyDBIsA9Er1qh529154A+XXhLO4T/Dc+qP1gUaqp2MzGfkjOkLPa2cgNH
whpVi2DTko8hb1KBwgrfcbIsWVHrujcmD6qFHtenLDN+ujeSzuEftJBHwQFodT/sCbHbfuogOBec
pfOHBqXXITMACiSoNb2ZLwyBl5PyEXoE87cGa7oeVFBnNsLt//14+o3Rocnck9BNNcNZMhw+1Akt
EGoiQSGaNPbWDrywVoSLtPT/IOLsp1zRKtj/O8Kh7tQ3zds3PtcSaD1pp004qbyxTx0DtlzaQRnL
8PLAps4T1AmFABUx6ar1AWY2gzHMRV9sZBQDgBMZ8xPHICKQq8ACxZZE4a6lHNdwTZ+4PRJNvqnx
q+7zXh/AxH1OH6cvu/3SR5aW5+Nu1xH3G00+x7teDnBGiTnKsIGOCjyUogJkSvDfe2G/ejCvtivn
HIf0GN/F9dVe8gj0Uzn8fVIez1BGTYCGeduR9mbWXZk0VOp6/OZOvW79s7j0/KlB1p4C5oSPhDfX
lEjRmisuXe9RdNcfHtgWraZmScf5JzWAxEGMp2OyLFquoWfMD8i1JlX3j8tESxNorkEYtNap+O7D
LEHcwoMeG5N7UDuP9oqQlsAzJsNhFOwA5KnqHpJ3Z3IUg62feNZbNzcMsTfAq65lPqjb92eJ/64w
gfh6y/Xc7UIL3yzCYFPrlWUmndbU807IbgR7n0tOnalfK4hUHg5pTbwuw8Vl4lwmCxPZNH9Jkrqp
J2gSsRvCDt7jIQ+khNNVnCbVZMGdxZQu+QCCUby1fYGV+uHtlWfnFYRX07+4P5osvzmvXPv/h0F3
xanCeQjW6W8wi56xg+aiwrTGA+6bZtcfWp4ol1PboBdbBvfnBVz2bixR5U4PVpZWpYEH/5HE0Opo
IFI9uok0rm1FhCIeEhq587mSu1ntAHfRl7yyHhDCoAPDE0cC/0Dut6u61XCmeaZoEydrZfFjgwj2
doiKbqMQx39WNXwv1pugYuEzFKJlQ0JONimRCUUcIQvtCOKTFWDNW3j8TCsoanVfQpotfyf8Bv1e
k/dk1SjMcR88UKvUZSJEClG5xnpFrWFSYCkxg8FlspxI/yrSIb8k0uX/KHsM0wEk5XHNqBlYxSjn
tRiwc9VPKx3RyAqzSy4bDw4E9ypA1+CCrtqotb5xyu4MOGgZSduBT8JXQKnoQSem6PRmo2MzKuCd
7bNr/vl5c6rHSwvf/N32bTIKos8mada07geZdizB3t6vEumn1Ytrjyc/zQlojHSOMbxs/3l0a86C
mXXcVqDxdTgg0KUIhvZ/jZm4wZEvFI5qcC66Gh9CrqPEPIixiYqC4FzqDZMQOEwwxtcc4Au15r6d
YLNgE9MI9n0udA6fw8wQBH1vMMkJZWbQLSNQT/wKYhCMYNMCMRc6jzZ8Tzo3WiQIMyJhSTZ6a8DL
FfAC0QW0rFdfKjStFHz48q8N5fOrDw+Pm4rezRZGNuPO21K2JZpzmEBni2ozxO4j0ehJBvjKK8Fp
sImqnFWHNkZkCOJzxaIrSWpn02pAF/3s9p8E2tDiFj8C7BvorKBTf7LVQoCzCWowy7jDhXnH8H0v
RUjuNmsJtg43Gje2ZMOg7KYmZmyfPFDLzSx1kv/PRTXCW5CjLxLnA4WJNkUGd78cZ19QUPijstW+
97plRTQ9JTMd3v9gkxE5WM5RhkGL61nB/CkcN8qEJmailN71hJ2RLOlu0kJFZHAuudl1+MrLSYSh
+KMEUIyjJMqxBfS9al54sVo/KeJa7ovcG0cLACI+WGC6axxaLUpOAePEKCii7RdvTNTFJpChX55p
KZiWOPROnyRvjP17VqrvKoVyV6i8jADu56RzabDPiV3FujTgw8LyBMA5SM6cI0aJraAM0ENcVWcn
DIcVdZlpKGPaTx91XVsRk3NzKKbKoPGJX8OLyXbrASWyp/pxVIhfH4mdZ8dSczF2z3fSoiQFlSpt
betK6nxpoKTz2WKA8WC9ph9ncGk/2SMWLrDNyLy+ZLQSUCSKGXw5pJVUhn9K3dY5hDOqBv/7J5Ug
vsWy4yW3IJ1+jwlwEiVGyKor61b0VtKmYY0+dQu1cYygWzq+85utSzWdEvv84ofCVq3FkXERTldr
iupLLJkhupVFPnB4sd3JtF1NCu+KGqhp6qN+rrBMy0JR7ss2Q4HZOtCIwIczSa0B4qNs7jHyL6YM
yqP2RHfAaUsD7xwza4+wD5iL8y+i/0/lFlOWSyoQTg8CRuQR7B4BZdsPIR7X4/iFtmk2uO75CU3T
FwbSVNcRnCxkts3R9Nph47jO3ukiMmTITIi4pwZB40ZcngT8sy2omAc6g6P06Ee/qR1z2cFM1OrA
Jysyp8U+dHsoOqNg+YJ758OUnipWFxy5VeWw5UQoX/mZbQ34uJkemraAn+ZgMm3SAcQRUMHbXq6n
nXTVq1Dk8taGV8hg2EaeDXdkKzDbW6B21QTyhTNQk25kWG4ga2fvfq8zQ5oyZz3zQ1A6LAcfDRa1
tCz9R/GgKbJLhkVK721WhjMo+5LcB/Zi+qzo1vK2S80ihBdOmid0lLNLwZcwMtXrZOPUnilSUYUy
H36qcq1Gn3K+MZBX21HHpMhTn3aiKZIwrlnjUlE98EzwqDChgaEyz5YQtXbFaglWm+TeVyVTuIHP
AARd0H5ivsNcPFdKt+D66zTfCXP0vLNKePZ5Qx3zcoQF6Yn81RNNtEC/EtxYcyaSygQ75mB3MKTb
wKct/txVZQ/xUF08K5g1dxwpsSJmhUmcHkqF9Pw2egtO6eQ1K3ClV2v8tcInQ/AZF11BOKFKN0gn
HftFX3m7vA3qwPk4jIrS+BTKIMaGB3Lx245zMW9wBHiYBdpKlJ2zcTYAJ2qW9+YXyE/1g786NZtd
MsY4WPImtdDqgfFLWkS2n9UVG+6jWDZMMlqZG2noZI+GJF3XED0q1StFCzO25eC1PLvO7u9+m/Y6
FBdMXJud4P96AtpaFjkvBDBAiYtSPIOwUg3+wG+JENvrYI0Z+9xmAN7gOhUOXn7WDWSJlnOB63PC
kT/8TknO2VU35Qt1yf5T6gVxgxJ6zTxtf41K48xpmtOjrS4Fx+wX+w1IUgNMWr+HixwfUq6MH4HD
yll/Kw6Zql37ea2/ZW2/dms7ufMdnp2F3BVcahtv91eRVvAyi2DWW3MgRcs/XOtP1iEYUipO7Ppa
VqBB9CXLxEDBxwNHzrfD50DsMyRNWO/j0PWlaBMQ2MahUVICWnQC72/fGM/258D6gp+JifK9h73Q
jx6JSMPnPP7Juf0njExVoYGtcrBs9ack7QZ/jXocyVhWDb9/0s9uXv7f2jWsufckQ1Bqfr9mTnQh
tIx+ZAtuc1IG51z0kXo1uC2By8X3mcCgt+GQv8MsL1KRfYxQBRVXoTjIP2zOIR7r2xNFsSpPRS9q
Li9W0FIiIqW21Dovtn/p2k9brdU98Ci3g2MTIRsSZ5pjCCwWEAPsRwhyucqUyk8Gfgckqy5FF2v1
gLITFPoqU85cW3U8OuvinR1RVXV+hFPLJygPKXwtXH+m4gy+54bBSZS+mQnngYdGVhdPsFWjaklX
44NIx1F7YIKy6bqxf1JSjXel6kn0sM4jnF1tD6bFskRhOYpm9T77eKRU/7XRmArMN7IL917VNY/F
ZUhfo6zZBBR+iIWjjncAVd7CKB3TCf6lKcIFiAMRersJCOAjsn1lHzBhCdcHs2ZJI+ePfcOfDGJR
I2OIKBbq0Yey+n5xXYQEsCPUq15nX33VsgJ865cL6SjBkc9pt90/HLDGssN7yj84MjFjSQizwzMp
rOHjo+VUVBPgOz4L933r5Yx6fLl7BTbjg9m86Uw7lnhY9GnDVrFCieOILE3xLECTQ7jFzwpRiHvx
awchHFnW1dzOuVM6yWsxHHboe+BV/fugVdMbgz8wUKF4gV5XclVJm4LobvDfwY0uC/sKAlqqDzIa
+bNxOetpbA7Kjf7TT/iHueWlmp0ufLBUmDYQlPpfFYtyuYQ03JYQZQgfB3SfZn8yEo4aWpBgKHvm
MLf2hiWYjtDJ351kmu0qteNxzr8iS9ZeUtFYxI8LMVb2121pOccsn6Xr26DQNWaHbBYqy9yN5OWl
ciJ6NviCldjeO+DVlDvTVOvkNyAEhKR/WEyYZkHbFOCNWWApDFp2s6bTpy4p0V9NAlmrfsv+rG9W
14XvkSwiF7Ly64xp0w20kLuf/A6s7h3K4JqnRpkAhGR0XqiVaAHv/kVNMYDe2id2i2wU9x/9lmes
3gRg0KGfefEhUNR4h1uG+/jLan75yNz98aYGHo3kQlW4BTpWHo1J+YiVs1Q8JURwmFnDaz+rRGNG
fgBtB919ij4+fSkzDGzfdKVOqSgXG0o7ZM0aJVzVO3d4vPXBkLLAYV2o1zll/9EEGrziNLhrE07N
HoNZ+OubRpLWMMsKJgUUDqI3cmFFnyXoGhYB0mktFjJIOB19KIt7mngCoWvIAZMMQSYs5VIHW/IH
7mAH3VsbleaFlyx6VGNjaDPTq7cUZCHQ4rA6VOIEG1OeCCdieOrYAzq0/wiUZSqfJetCASdmbEdX
S+kV+Gs2L4Kt4rjxQ/QDmm3d6iimqHFWOp6TLihf9R4HJdg8poNkGDwt5oiJgb8Gub+y9Ce/pfu5
3Ka60PWWED8mPfRTRtsZapCernsU0qMpL1EvqY6FzMQCtTTTVKGEYOTETTmIPJ/b/GCWaIONlOgx
lyJBVr/iI2f/vW/Ff656geiMSXbkxyaLJdwjPCdWHDvcmGfk0gi16ImjoobH/RkblUuDTfnkReic
yi5eNg10LsigAMEYKd4rmlrFvveXRtaYcYEJ4nNyDLGAjbcsZAqqQidoMNjYa31qwdDH3ZejL44J
ihPmHQ80FeyRwjsFe1LOCpYlL5zNzmZAYz342ws5odwh9Gvam7vicBuDa3rUzzBaHeJLvPzt33tQ
P0Z6ayyLOJu/DTKatwZ3OZMV35vtGrXNdVgwHX+aHQe8n8aenXHyN+qNXLp/T2IpYb6PUmmGybdj
QLPHHu/qTwJCg6qvDzY9DmjjCAJqUooe/7dsrEvtnW4NdfaAnwbVxEeUYZxMxHZtxy8rTUWbppw8
/wrfYpBdr8t+IWV+N4LTW6WmfuUm8dDVR68zr2A0+02fqwnbHM5miUUVdVILKAGD/Gyoj/uJZLwD
i4oyvbQRAmhV7YVi7JooYV4uyAdIJ7A4NRIPMLm8YkqqnOzvtd063QzNfyOl81vPwe5qTib5oK83
RTMsSxMYW0w44SzG4hNB/q6lCy63tHOLtp8BAlw5tKbeNN0W+qt588s+1BwJty9Snuo/TOjQZD1P
nNqk7b0iulYk/maqtS7yQCigPKA4v++KIdjka9entYT8M6yN/4eZ6poFd342C6Tv0Cl+3mp/UNYY
bhDLLNsw2ubDH3+w7RNZwG5WxMWPPZUE2ZzbR+bPI3fwtrlG7F6Q3aRtKXYp2ap2yQkpT+RVcW7B
8hErs4DVDr9YaKc2P7IG4fgARz5A5a5xIZQvJip64YlBfJ5Jr3QWw8bmGg5onavdCXUXWvq6REf6
qHbgyBFLizVStL4RtoIxsMrN6XsFGOacEEQ0uawudLcR/dET/YK4ObYlnIOcma7ZdAUNGwewlaCC
3vJA7wuZL7IKrtVtByFZSro8PPIaN4vhVI1TbvDAlzNHqq8c/iK/z7Z9XzQvNyaJOA0ZkpB9GbSI
69zTbRpArOlDsCx1sy5A3rgnMWrbN+Tu7Hpwomd1urIi16dl0jFOzs8ykJnPMNnM4hqxgZLkunIU
5+dU1/vBwYnWyxO1bySVqMytEiZP9Q++thdoGoHYfqXm5i76yL9srtapZaihBSGEc4dOmjF6XObv
mizfmxG28jy2Wj0H8le5pvAGvcSOaY1qXbAc8TobkRpAGJlrIsTB2pPiXI/yvgu2ctBPdlWJAqWk
aA42hwL3ogFK+iRknoW8zz9xYTYHT36yclW2gdXf7XCu4DrYSUM3XKzv01SmfgACOvM7wKa07YLW
VY7kVuNzu69DY/zTaACTAMGJGXBG3fpUxTa0+aa4W456HPd3RqD10S453d2+N8lxjA6qQQcbJrPy
RTJJiGNKLKygz2ySGvfzFxbKoJCw7bSsM8GNAhTNmIhtjwGF5sDdTlQfP8Tnqmd5lVKs0IzRfCuS
wkVm1Sbm7PjXhazNLNbD8YzKHSCEk6ypwEwzNwmk5vDrhwPJfp+nsiay5WFQz5TLAvh5IEovcMmN
V/ay+Kb/f/LKjvAg9ZIjjA74VZucR2PYTtLwinF2QrNcVKCMM7149NGKzBCIZo7pmEMRxHghyUQ1
/DkBz/5/u5Ih3k64xzH1DMw+nU61e5qSZi7zNnzru67MhLK5cl89/aWo/VlnetXQvGjEx9zag5OD
pxOpy4Vlnr4+eIpWcYOfRnGiB7bEh7s4p702iSaaCNj3UoWj08EIf3ijNienA9vqM/bfUJAutHzB
Ear2X1OueG0xj8qHEwIrsMqOPG1TJ6kjKrktsP/t1NjN1wPHAAPhevjxJdjWoqciwThFKHXsgWD0
9nEU3Rtg29zGvUbP5NTvS4Tufb69xVQTj9FQxPN5rpkMIYQCW0QMigBpsYmdGbXhpX+bDfVLoAUF
GDCjD3Ar0Q3ojLT70pjPIJEbxq7nBkaOGSyJCSvd6LT33r43PLsZmOdj7WXUJjlB+6w5fXTkp+Yh
241Mz7EB4S4kMxw/0BGOmy7/2TQxXut/EZd6v36AS+tjcRdfqlhBmgWu4EDX9RiMJ5ZCaZdAPlhx
y2EXfIYkAT13xmVsEjLjhGBklMWnszRTkGeJhAq1YF/US6HmQqFOUNF8xc4KWGPlrx2QBLrSEHQp
SCvKU5nK5E1OSmQ+K/Z4rV1dR1/FpdzwIl5QT2e22Fl9pFiwikjYZlyRRXTCkV2ztK58sguLWzxa
nkaWdI+xPyyAk+c6Mh75/71sFEqrphn2LnTGZzw6nBD1tnSz92x0wEpbuitITK9LzvjcOHmKze5/
m4PgYpLcN8J65yu01yJeG8NmnikuUVI4Gwl5j4zJAoeVixX9VAqXO51l9W/4qtvm48WVgWPqSNwM
XMFn9sb0nJ1/0UMbLqU6IgfW5GTX13sK6EWQ59bVK+0pB9w7d7S3IqlMEAoFb2mNm/RIvzO0wz6y
UqyjtTAb1lqU0OyvAbioKGLv0x0h7AqXYJ63OqcBI2fcKBrgxFvygbpeHp+Um4KXF+KUnXCtqUci
1lMiuBt1yQCkTiT9rgDogHdvX0zR/Q6wwCDS4fD3+GW5D1RI3iMmsJEl+cB0YjvIo40b13hPCqLB
pUWRYLq++PiAWtklV/uMSgbjFfKLEP+GCWXcLG+N0pT3exIIfz7KZvoPWacptSG4WiXM1oJz1P83
X6WfB4AY7eN4053WHlK9UwBmvfg9/1ETLFIyDhI66UNrnWubVL3AQNTte5E+JJBMI6ChozkD5M+l
ctHe98wxiykgyyvUWk3dnx9cFJEEgrvXX4ZDTqGlCAO30s935BeYZJxuzIoB2RPisOztfCP0bvIs
7RvQgUe2I+6C5WuIarzRt1DXxpu2YnkwkYAM+Wn0JigDTx8e9drewx9OUwo9BUuldtnvK29xIxx6
7jCl5lZqWerf4/Uv/aYRmLuWc/kYJStGUg42Pwj8KJ9MvWeNJJc1WZEEOHi9Gsu00hH1YtoX3PRn
1/DXaA3DnPrBmOBYyjVosDqX4SgDZ/a2ZhPB1rNKXhwYOKJBgrEDwfTzmO7/oOosrx6RtVpRpeEp
2Oo0n9IaIgRmpRa3no+7KEg9Md8+xuFoQWJITgNENTK1+uOWzkeCEOrF4FNunePUcb5Rpue0bdj/
ndRxXxNj5p5i5R8+xAOLb/1cybul5S1CihkGnTOTDoYD7wzFop2+nWt5+Dt5eZ/LS2mjqyKWopS8
N6bTs6IWLzBuSxyAvBtUcJjQosrSr1cHHjx0elsxOVen3OxctWXDlUSsTIaI/Zb7O7gq9ja1NHWe
UV32JLISwwrB79Oh1gWh2Q6k3OcybBcvB11BCkh4NgVWVXWX4RdhabtO8oi7sW5NjjQ59l5MoXk6
nR2BknNhVzdflNg+0ou7+RvywIkBRsla1GL0PUHV/VO5ZuQgVT0qm1jYk0QIl5hDqecZDjsguA+v
93zeMNX6AP7P0qfbjbge1WirQpxUh2dNkuugIvE/fPTbkGAdCczM+nmpXDeiLg4QOXqE6Yib5oD7
QlIBmQdJic/bNVHGDtGK3wBmoAfWHSuiQ/LPfsNVoQei9wkPZcLHJXgKF2rj87rOi/5+V/HhA/ZT
rN69iu5kSQtab3NjlNXNE/FQsZCIwlDBCoHfGL12HgcM/4K8q/sEXhfVwGvGwrJUecfLQ87tkD+v
Nuj3G3FTMobVguEjZMs+clLEhDd+mqTLjdB4+dgQWX+shttv93DsTJU9zb3ojSrt0KWUX698h7L2
M3nFGQJRBMdkG2VpBXUC4gJff1zrn/5XcdNhhBsZnhE5ZZgYXuAxMTEa1vXW8BY9abkSR8BnvM1F
ha6zCBNzi8sKWTFFc5Uhdrec4Gt7W7nYle0O2gELAiKMcEMz4PF2/KZ2B8ZIplRhSEseDUMG8qt5
Hq9MistLFXgUTu39c9YLnkQ9Y5EPvhicHfOFxC26IAELC22RdHoDP6HotzLsOQiBXLFdTyYz6QlC
/MsJO4Qu0JuSLP/YYr+kGWcENCOAUh/oGZToX/8JppDgVsY5hNoo2awO7asbJt8B5nHQqE8tFQiJ
prnNyxqJa414/Bt8M3BZIWhWxg+b34n1mp6bKqnmY7WoUEh5RYY6xsGnRb/NoyIGLTsYnDhtEHu7
z+oyIArCn5336klZjvsRX+ygdRPB4ilXwmM71xjw/bobsVKrxRNYeEsyl5FIyNiZLWsLwD2RKwrO
UsHLBp0NhLCO5mesAbazy8FykbSkNfsedQRRUNKTBLwkOeV0Jz1KYzDUeau5TvjbvN4sQtHMAHuH
k7bwJCC+RTnyNuWseQBfHzDx0sO3PPCsSrHWjeM0WqksrjPbu2zlWVWWmC5q95ATwsCIs9TxS1+o
iLZ25bqCRO/V0XeYiMMDv0xcXl0sp9no4Po352IEMMbfmOHdwd854npLYTNOG9tGtD8JnYQLnCSp
zKI3zVVaXuzh7WtOuarM6Y2fGEA/3rvOkhoUhVIxUcsOTRJ1cSatuD6veSIhMvwa8MNrsC+x2Th5
70qOfEjSA3JI4+/Q+M70/69r4ZfIlMvEY1i9NeujlJluZXkhL4EKCdy+5lSgN0/dszL+n6Hxc4Rm
FuFjqvCneHHAusVbNHu2wREWeTpw/PGJk09jIF/8VCZ6q/hv5Gs5u1eUnyTCsl2piKXLx5HVKnYh
3gxx4wtB7UJ+YRtK8HfT6fEQUm1owl3s5I4YRjZR801ungvioXCVulin9+gLY2XK2xse5UEwVHqe
TON6+ZQMfu7tjrSZzWxSsDKxPz+3r/AsTyO+u99kkowXJ68WP3wmo7sVbLPz/kysc/1IYBgR+vSv
QW1dlfuWBsk7QtmViNkDDn5XiB/baqg/dUzgDoOYFbQVQZLiE/Uo/rSB7G4Y5q4OYUlAJV+/qv0q
im3VPnImk9mz40yXULzILI7EjYrrEg8PtP4GTqZfx/6aHO+COEEXiPREP4S19hscGfcVC3jgCDor
yPnZ1io3wo/4OM1cyapk3st01LqIhz1X37AH6rvcZ4zWX1Wkx0QvP4qgFTkVcwoDSk0qeSCaJXAJ
lEbVxp0MGQhPztCHJCMnGaYQ5UBJqlpx7iNEuqyhaY0OPGMxxPDnNvBTGEBtOZTNhfyRpwq4YQrW
1pZxrJ0aF3h6RVNJlQhxjzVEo4zgoCkslWXNzyG9Z5i27fzt7JU18ZSzair9h2q+SZmfdBHCBhw8
Z2EzixeVYkI5zbqkib+ZkOqTbYjDWdiUvAYpmGHOESPwkh240TFNsYJNCC/jTvwYsuXv9q/zQKqU
XM7D+/hBoG+L35+GDwP4Ia3YI9mc5PT70XFMuQiiesEDCkYJaLaDRnmP+VlBFU882Yh9hAxkxGYA
X2lao1iE8AzsCKt9idC088RtJm9VaGzUYZxSk3vTxezoiDNKvXErEPK4LQBJ/dqzbM0JDTh1OeK1
bl9bfxQuBraYCh2SSLiSZxvU2Cuakl6whpZWbhBAYKqwxX1+yN4OjoVmcRxjJoBWhLyk0MrsRt/Z
Eu8wqJY+Pc+uWF9iQsFTm3q3I3BB2IeoDZB8Q3ALnQ6m7QUu4b7WKi91RIVUJaK9404YcTQQIyXB
Qcn9pWOZQZv9a21/PiGGQJB433FCekovZTr5VZV8fZsaUs8FPbC7C0os8TETb+RvtlxbgHOCY9vJ
4tNZufpv+KfxxIsO5+xglRkt0aZHRKU4J/AGTfq/0y2uhWkkfwcPpb37YLy0hhWHPSQ9b6SDc+Ki
BBDDPT+SySzpI4IA9IGsMdVEs5JoS48XyVrmXa0K6gp0g/xuKA/k17JQGilcwv7RZCl/P/nHJ0TJ
UV0oiStOlxWGoAZh2WQYE0CtxscsabVrDcDzLW/LxH+vGs50Znurl6ZadbnTkTt4pcaKpz3ussX4
vjT+kVBzO5kJBjQdBmKRT3UH8odWDVPjAlDMHL5+b6xdp+3ODLeK4awKuqdr+C44EznVP0Jdz3Ma
Uppj7WbokAxwlyzTgzYzY5Q6dWDq4yCTg6Jy5Rx1J7KNs9V+vwBrCKaeoM0Xa4jFwqdAssxhwm8s
q3NGA9bmG5fLklC7jydz78TGrx8ZcuCLhZKsmlDQbWkcmS4mRwiP5dR4MCZBEs0WxPtzmOPey7//
1xZvsycAh6ZpWi+4V/FTaclR8yJZj/SY7BiO2uQOkCdrL5f6z/lJRiGJtEP/2zE8a0s+Nd9Ve6LY
OVn2bO4A7EV5pyUb5RTMnLYNXnqUCxIKY9V+W+Z1G4UFoc4B6B92N1sLKPuuJIEuL3aDWlHUAbuN
XqrXCstnRGiE29k68i5ha61w9QYQ9pZFnzyFqxJencu4+tULQbRG+M/mwnALC8r6RgRIs7ZGTWwA
liKyN/SjKHAkjpdEWN0AjKHDd/+rp1x5rtU7mWNdG/eoqOJx1bs+uDbCF5ai5RZeWJmvBG1H3Y1o
vai3czcXIwP625a7P3DjV3bSogi8y9prCIh9glvB13kmdoqviNXmjyuhinXRkvDEWJi4rBad8nDt
NUTrEJF0Cf8zAIzpsC2adiDHGifP1AcNQuYecfvEnBkg/pjZagP2AgVFv+6RckoSfXnGRfUdrF5u
yaHZnWUcN08pnzFjDdTcPmfiJFF91YFTrga3yb+wnga+4Qy2V5X4jHErOIgqbGqlCnezL1FsaBAL
uTGzTtNOCp/j2UPOCiTpF97khKuox159fw/3RMalHzpv9ccCVSXXBkhq8AWR9fOyp/cMFEhJNSwc
5W8At70UrxeDnDd1Go+ZWJcnwQSAyhdyO62SrLA5TOzg3KU3jIccl3mq2Y7pSSE1/NaEfOU02PtX
TYsAqukjlZfSg1q0rOcBJIw5w5fuPWTAKZv/dlxzMtofBBvibRfbg+TRN7gwKYWRF5XaXP5941IY
/EsWhnW5k+y3qOEoRr8PnsDSHpE9HHrAbB39jWu5wc2GVxRMGnw9cGDBlyCQYBfaOParLPZl/QpB
0x/N9sqkNJGA457M9gfllCojQc67gNVI041Muea6Yviwp5bGONF0QfZMcUHeN6f44Fnb4ce5AJbE
0gW1ZZ/S09LKoUISnrDwNLXZsgPYEFqWWr+ad9wywtWwy6EBr4l22wEauxzpw2vuG3gbmh36hLfi
auwKRnWGIkJXWrjMeJjsXfQLdv5Q1Uai+VKH4GAWtUZLH8Z0l4+DKxFySqLuSEozL2aU4ss9xMmb
7ThjQJ27nchCv5BUzlbdfXR5e1Zlh+WqWZXG6cyhMATVgTo++50IHD8JSIVwiTpnplINXFmqzQvW
ROrp6s65wF6aCbkETk9fZJsKIVU7F5MSWLCySuDPrc0sYFGtE/4Plq0chwWcKm+5Qr7afcsW0eo9
0BCHOEYjXsJSTKrVOtxagLnNxZSi3AUKe5T3QPcsYRWZEQO8KOrfWSi3hyZLczkEsV4YB08UCg9q
RDwEwv/U7AFBNDetL+//0PUAAAVmwYHAGp6bZgIwLw2OFiLGYGHf1oC1Nh1DSqfUN/yZBvYqGTEf
k+s1jD8WU5mHFTK7PdeMz8fwU3zMQ1RLiOvTkbNTFQBIDdk3QH9MlmyO4vJMfpMwI8c/Yr//fzqF
j7a7TGBbMdy4eq6skxiUrboPWDARFUW5BOx2QvAcrITzoP8pY6BoEDBT1yzWaOPPFE7bAW3BVNKm
3PB0/kgu24eBqX5z3CwDoFZsF8bTTdNEAq8sYvwCACFt+vJpqTUKP1ljRUKLwag5U5eShjKLXGSD
ix4cztKzy1p7d4FN+2ZN2pixGzJWUZCTFg1SKuhkphwZGiM/FBORyqkkrPjMXKFBi/zS+K8gwFei
bYvEApCBt0IuctgTo2tOR29tyWRO/aR+cVctAs1bHYyuQppOU6e4ijWJIua1VcvzMFW9HOHoteIq
K74mkCZGVn2cZUl90TU/PSzEsZXrTqciWLOEhVSAlw5iFLKO7qgj65RS8Q8T1cgcfTMhO8l8EDOn
t+zwcav/QYf65nzICY4Sqqz5iWvwpr9PJ4riThFSFQDaS9rxAO/mdJOnO3YsRWCVDYZW4Xi2pC8X
bThLJ/ZJfCFZstr0qrdoT4mz6WSWzcl9oQ+m6rF4qX+TTCPQ7IIKqdU1oVmMI0rf0V88HHm9GmBQ
Ac1RiJ6UFTFgIUPIvXlCpwQFNBuyRkikFt7EfTnFz+NuX1paL6IGMCvoIOa3GgrmQVf+N2qZM2v0
Ahyzy1IMuCFK9Zd0VnVk5RTpq6YVK0obRmDHlW1haZvAwsSpV9NN0Lhlzq07lQpjMldhtppG72Ej
HbC9PycG3edUFTE3nRKLJHIQNgtlcdeeQmtZb+4Uw9fKHP9egzlkgAYjUXTb2kys7R+oV60nikQl
E0GmR2PepwU5yqYA9ji5qhgte1Ohmf3Mk4lqDY+ef8etchJ+fmsbI+BBmfSdG6JuHrwNv2sH6Wmv
Gco0ZD0LcBrlkM1W0r2BbaOAY9hjtYP6hwqA9HDIHDhu9OPSP+G7p7H4gqSlvxeQKM1pIIcc3+bz
ota4NxsyU+wmPheceGKd/Wlwq0xtYNxwHs4bMMhqsTq8itz+N/dhGuCyaAKDzpZriMk3omzAQOzX
eVdSis/JLBKZ7BUxVchqUFvB8gwTPSJpxJYKJN4NlAu4VtUrTussOi2WXnxS/adTENbc0wq2Eyhr
AalOPyLYkiyAQiHBTDpewxJdOoNPNKEkJ/AIuc5HxhxqYQtnVJQrWJX/33jIJoDlyNMRAptYqb+T
/BXBPZXOK4BUsv3/4HaYx7bnsppxcrZCVinOahghTnDIkdA3By2uLi7My0e5rd645ICkdvlxtF7W
rWr0A0zBe/p+Igr//6PbTEZfTYDO72COAt1lx1e30n1cHa1jichHlExCgzpr/2OP5HQGT9xObnLZ
5ki/k/6l414p5hO67He5sS9RKzzoCKBPjkKm1h8FKYYTvcApBzlZx9/lKAZnGm/R5VCcjSGzMRNU
1cQ+2WFvJwcpaFz+yo5mUrYapQpvuN5jC6v9dqN1+UPnjcnNsf7u6BqxpDPffepDC1SpCcyH//+U
cIRlOzzeVAZCynLUqg7EIDzJpXbdLSpmPaRS2FTXbE9FwZHLACGL2lSSuglQOhQMViRb+osovUJJ
pJnPcJ/rFeqV7w3SPULXicreLLKwXzz6oYdkGAwErKJUUfLa9XIN1pRouYHwwDfh5d1HNWFd/cOq
iiTFIoRxWxqC9Q7BN397rlfKJ/bq+GTcS0LaTsThGVhu3K5Dm+DRDULi8Z/7aQRwS3qaYGZy3PmV
UhuFera+ixKMog3Yd3JJGbN48Rjr6SNsqmvP/3Yh+cCGB0HOEUo07TW7L97jFZwV1q2I3mYlbSe2
cztn6VVwFUsOC/M/EAYnG6o8ABC2jvs5ZgR+pJU5sFm0ImGTSSKKFeFHWok9pKTTsVgfplE+jEjw
uUAARVumydOxCI6FUq2duHuI5HJHyScXViXXQUH9xHo67525JHOABeREGcngpAk+4yfzGQsfScES
fgbx5MNAeYid3e55af90RC9PVnHUYcJW41j93yGL8qUz3vhsTAO21eDnGSzw0zg5+gM/YrUTIh9g
tHZ6rTIGgF5RL20vBrjyNYaLfdXAgFy21lnMDD4CRLie9JY65cjJs7yLNq0kUUFa0gimg+8ZN/qD
x+APpyKAf63Xol+NjNEHk7nTG3+w0Ric6vGKwSFm4942CxpwPfkmK7v4lppUvw3UknE0U/nw1JR7
Q4DONfb2Kk/leBbAbagwQwNLxpiyjHd2DySHasz04YPjKPkJry49GnYMu5w9nbxzOYHtlH5+UhfN
Y9hhDnoI/eH8mQedXf4JGOVjw1ZCJNJhVB9ITW2af16SQ+cYssNuu43xJL7/GOrxqEXwF7RcKztk
oZlVvQd4nYBSbesTvae7QYqXiS5cYFj93J2uXQNx2N9cAsN/LV/6VyFJ0xRi52je45H+AIfNmy7U
oJ0SOj/B1Obwsmj/tfA45MmOCkKiyiEYdnk5BeeE8iQc4Qz+phvLfOda2hQ3RLRSJtRGqO5Fiprz
xtQjFI2j9lQvaHsrfz4vrBpYdFyM13bqrBEH2sZ/9C/cUV7lmK44XnLq3xaK8opxpjdsSzkeWYRp
0IKbQGXXIrNB928kkXSBt6cGyyJkUkgvVeqeckQEfcmtyWSTjonB/cNgacXEnMLltS22HDWhAL1g
oQnpa+b0W/wXh5Z41nmvPRfCbfb22Qi6kUkgReukHn1geydfINttbNZE6wVDPnmkW2H8RvqOcD7/
0MrCfqqjq92F22Ns+OL21ShBUja8OWB1mkHzOEiKKmOg9p8BkCRfwQA1ZnVLIGH6sTdRJp1vxGmJ
7Lx5j2eb82oF0EpTW0WdF0dWAHhAZ6uWc1GfCz1RoG6auraioYovwfk/Lytl3eJFzU1obnrslLAP
Y79JfmHC0dRPEwmXgJ7WFdCdJcJ3WHjwOZJJDfnESrG/2J3qd60qSfwhzpQlq6PQBc4Ih8QVu58Y
sWj49rOH5yK+/yzA/QvouPQXdODqBfgENnLGpuMTZbWrpt+KCSAiACMTzVUbr5852D1YbhcgiVcU
M45711clUvb+ufoXH2//sQpatk+8jdBWpAoWoHJg9UHqpH45KBbMKxulV/oU/yYxfDyV2AOIrbMm
2/o7L96fs4yTTcxBbgEp7Uxhb6Nq4MrJtSYubUBES6nOzKECuQYObGRGTgPPstp36BqZbfFbXsKH
lpQwAinniSEOKtHNHho/TSxWURbKdusDdd2JJCWl4y1taNYaePiwbEbYve1oMmvb+oTq0jZktsWn
dG5gH19UDqAX4dF3XGGAW+gHIKHMHYNTlPaSLbBVXBbOG8iHZX6Br/ZFhEbZag7Vq2wxateUXBc/
+3XzlyUQAx/9kFonFVrItV9DUoqO/udszxNnI8wEEkFIWARsIrKr6RM/ieTbXMdWw99azyFSXpMd
gAVTLTVmlnn8v21dZCQtovk4dZdEukUQ9Gd/gG0HKpJv/HjdY4nTccfg5+evna+kFFhByM4Pre7Y
RsggwONQDAQuTEfxllh9FxcSfPvC64t0PBQ7ikDbFeQSR5SsaCpdc9Kyy0yvqbLAsDye4XG62QNq
NLumz6jdx8pm9GG1+PZ/2SR2s6vXTRI9GHONYXMTYD5S4/owQd0209wEH+UwmwwBpbEP3b4AfULU
UeGAWUnWMJk9bcIF6oHrvwRHJXBHaWggdmc/9b7twj60d5abXLW1WQgmi7fOGxFJUt6A0VD993JN
BjrRMrY1i7k34/tfO8A28L6/xYezgDtjlONa0OMtlf8a0oMN1WnGjXYkCD3/SiwcpZzARGLyl5VY
DRM2QbijUbMm3Rnb5IMmeUCkk+VgUagvHa+J2SY+IltcyczVpZxFsJaOln5NQo7CsC4n/tNLta0r
40/XiOJH0hMIFvZTP4omnrsa8IjgjDwnAOU3/vVFBO7Awcm9ibtlvESxX5Khq5HYyVKb/O8Iw8a1
kM7fHkh9CX/5GV4gUFIW01kzjNmPUpfxhz0pQkj9h/10PLNYrkriP7dnlMHikbvcGJ6mG0DTPtEa
n7XKx5YTMgCoTJLTN2aTuCqq8U+xZGj3HdkrFyH5o+tAOHYM7gk2b2v0S2Rup5wr57yGayaAqbJ/
XHTJbGh9zfAU2uCa956UPWyp1gZvG5DcHoHnw3CIa94fNAwvShVBbeKHONVNRdEgRtSvNUT9ZD8Z
smx8bJLpcUDl1OXsK64RCj7adXxABXOTLeboF9e41FETjgid3aLhwIK5VIS/oRF6agjj4deqmprm
YXWITWk6sUqzjNjvPkhDpIePscIigkFTzhYyjuB+i6dqvrvkuLQkBY9uaZ0mH++TYYN2u6jHLjaf
Edz7axLd8YLrd+6+/E6WI8a/TtiX8/P8qc97oBDGTCEGTdrMRFkiETGFiZCQWfOn1QUu38/mVEiI
Ma2+MaZ5VfRoXaNZAjoXNx9/twNiFOe9FRNMZr9J6leWUCeaTxZa494S7pyR0XDlrV23WbgmDyFa
nYlehBFcl/TdC+QIC7O8uejh9o95RUF8Su/pwzk4034INQI6MSz7puAj3nV2EMrPeqG3/jdU/kHX
gWcFshAeKMSLn/aYgAnFtoO2p4blGIWxpPAEkpWcjGFEKOE0HAahVu82RjccJdrimzsTpVt0dapA
RtqSPVsu64mHZN+eiQsMWgfBExXk+buImSGPyHt2NSQN2KkBYeQs4LRsdgiqyrlHZ5i6PWLtn0VC
wYHxg3uLNjO1nCtYOpo7THGN7Pb69kR3oL3cic14IaEALk6Sx56xwdskm/Ta7+2OY4TqXVtwSSOb
6oNtQfy9Tw16CM3NdfNEv3Bow5bW8tp2kXhWbYsibTgnLZaDBEngtDoRy2Xfipw7dgFt0f0Onr6v
1fqo3oIcYBC8tZCKVLOgkp6g+Ds4fshlbVFc232RiVJ2hDvMd7RAjr600qZZuELeD+54IAxTaDhK
JYtHU6qfT0DQl7PfjkYT13YAHS9Y0Vey+XnEycBcBTMoFB98S0KzdpbHeRGefbXq3+IafV0xyDud
h+V3YgWFcPC19yXBZ/R99U2s9P2skuSyNh3TLDCSIZ1222aHfdPYLXWBsLCJOfrBbDecuy3ddGin
gKFeAWN22X53QvbpxRb5KxznEC4ASxVsK2LqO3evL3WHYacQx4a9rwUPJs+RYKXCxVmwDriVuIgE
Au79da2LqEWn6BFKd7gbBEmLpdCrw3DT7kMcgDLLH5Fe/5oZBlRsW2kgUiaCys8jdMlkxuzPyBvA
WbAlezzKZn6xMZPBPkxVYrASq/7TgHQqeMnj8PTEje3UZ8F6g0I7GbzfIJyULU66ij0xES18WWc2
u/rCMD0om+AnZ/l7NbqAxnyHNcCUEKyP6raPo+/oocddLM8sSESXrUzCrrJ9tVgdxkNoISCnHHHu
JqZk6mnvYbPjJW7ilTL/1WkMS+0zDk08YeQvgiHZwjxj/ebv+f8vB5nT9KzPBz4lBrhQ2OEtHcH+
wssEx9jPrb0ge2OTW2+A8SI91UnlHbBYiyGRxds/FFM2FLOjztO5sjlw//DznNtUY2G89I6mXGCv
ThaZXD55YrF7ePBazgJSOMAulpZC+ogztRGsfNmFy/Q4qso/LVFjl4u2VOLYOBdqFOJnIbT8sKJI
YZL+wWp/LeBoQ+IUkwfa6dDGy9Ia0M5Mthi9SKnkRCJ0pF7dx59TplK+7DYzL/Ow5VktHB8RlrB+
zME+csuqUz891GtOogV5MT36tlh5HuUbRyxPeINTjjR3H1KuuGNggDmsUOJwsaZe0UdhR+/hZhzq
zaMckTfZ+fkq24nlnTiLmKHZW37PeHMqR1OEIlvLcDx1FWMi0CtAKl+MTwJSNi1xduc8C2KWBRde
pt//GzzxNg7I3cViPabxeEQSGwL14IHQ/cck3Wtyzst7CLdfYyUaih0DxjwGnP8E8Wci21dKr8gG
eGFebIk4PiDhzXzuHVmcLpCouSJhHqWO7vPaZQW8e3SnzMXFv54JfdCKHZa2Oo2mTWO76xNuBr3r
NuXcTJQ07IsUjr+GjRNAEvL4YMEAFZQM7V/xN45fs4ZdXupi3/T5p0y8Fvg1b01SCAssdgV1t+JH
Y9tt9Ja+uJDXcqQpe3LGaxrOAu+0ydb9v/g4skMU+ronXuQqqC0bQRmLjv3eioruJq5sIWvE5ZZO
zJTSuDeOLaIauknvU4KOsWapOQCMUCqPxldn0S7N53apw/+JdwmG/1sHXMxl5Zf+bwYfyWWLRLz5
+nLw+HL1Kz9ZRvMyOauCDcBU21ASGKvGh/Dd8W9/5LgKaNYUTzxXjjqwFBqTi921wn0VshXo9ygE
ZA77iJxzG9X2Pyt4s3VyhuYGh0soRqeRniIrpuzV2tGtXVoIpmbEuKS+ciOqDFSo3LXmgnItq99X
89IxcdFyALk0gMD35GF0zmv21C9H/Wwbs4tXEFcJliblhG5fXAEpHVyhIaCQ8yp2qXpnFw3QEuML
GS3/8QpqfYO+mUxSIuJ3iqK5etGkixQ2jRuuPVWLtg87+gfJ+K9hwGN8bD91LDmSb81qMZERVtE3
Rct7nMVESSHghENg0+VsdNf+LbZfZOcvApRaNubBylz7UkgenlYvmWM8eUlSsVi32tAW89fjMEIc
G4I3ck3FGLStifETUvQTv6rmZKKIcwwK113bUeWMqrhMuJVZGe7uqf4LCEKigwaJXMPU/u92n8/K
lOB+Wyp4yAfsWZzRKldj6/CpOB1slV8C55FabFBstk+h5/7wHeKm/sT/TAmcCKUrg/cvN5TaN/m8
+VAGA8N1QivsWam+ASMWlU4OqjUiuRRHZLRiGH4e5MJXcbs8Z3bggJ613F+dsEBcHPi2naeQv67Z
fwrxjutYW/CoEu8s1Kb1wGtfC4Xb4dUFSJWPn+dKI3qdHWywt51EBVmfb4oMjYOpE9txfxN31s8i
SWFdgDFG7aOhLkXdBI5FG4mk81XtyTCfLeeQtQxAVgl9ZBrQARJ8OM5REm5oEUub1yvn3b70gSn3
Ki5AQGwqkuy37npqNZNyO7ezGs426E/wHGlR8jN7axajua8pjwjzYVygPAoZmGw9iEsdOcXuxLW0
Mln/7KEKlzn0TfGzXsZWnF1HeyQASvBGTHfBV6r4p3kKPR5GLg5RbjIwpo6d1aYF+ARUQbnibH9k
ZVtd0ekokuS9csmKmUxEAtI7SL8Mfwjx4/K8UewpFX3UeRncthQxicQ6PNwfNURgVjsO0DIFQzcd
GgO3CiOBwBk3yXikLqf/A1ji2zHgZw9SAeugpb8mJ7m8D6qCNsHYQdkWzljjsF3rrGa/+ux71JFi
LpHna6H+rGudk8QZc6A9XOKFyGXjV+RM2OHtAU24ctk4v2TCKWGnPJrKQSquhrlsqSs8WyRq6rBa
9e1RruSMWPOX9BtzHGvjF39xTGlEjW493Rr1VxJcUyzsQUvG9TUK02a/sA+g06zdrEMULoleXklk
dtHgpTb0Zqm2NFhm9aad6Xa6VToitO3txIkDcwkIFDVZF0oBDP5Pjo9oFD7/rdJxb9zmRf8cBfhy
sDiVGb5hvipd1AfKj7Z6BZI41Fb7I6bfTLv788isjhcI/cx0U48BgCB6JCC6mtzmXP8Xdnl2IElX
jrGaPZ7gFgrdZsLCFQMQoC6Y/e2sNCLs487Vlyjm7MFFFq2YojYZAcFKQlW05iBU3kKAW0UIIqdW
NpatjPwaHeakVOEcK79jiHZsg2Q+pUpCNGg4HFWFbXJD+YynTA14ugC0haYYAaZGszYwAMebypVc
1cR8/mEm5i/jhfY+rcXfAYMlJPi0XgoTlRNQ8af8ePzHf0qdMpLushArYwT9vhdNgj56Qx2NJa+P
grCE2F3B0vH3xuUlqEc1Cdc3pz8woFbEvSo7jjg0iifmRNnm5yTGaKonuPfdOzEAa30Rd7TUDDTr
Vmd4WjfXkASN2z0Yj01GKQ9RYIpI7tBjYDU8JOu5Kuli2aCFSn8GJcWMuIG1oBABbaqM4Vs1rXjn
F0cqIUe9Bip2O8jyhCOK/Gpqp6uCCe7m9jzWqlnj4PUfwHhzgEPqLNeO2E4gzFigS3IRTrPH5yt+
FIRXR557RYoFNyLVj8K0u980fx/iy1BjXVZOOj4x7+OsUm1w5VQcJdN7epb/kNTcVFGIW72rZ8ML
Qm1uCO4NAF1LRlW/seFVxsBXzS+tLyGBhsdqip2HivVloLfZUDCN57DiaYOpGq5jyqAiaLvOxZiZ
HGLyY+HFr4N3/iy6NZ6TRiMoqT33Y8N5/1S1UVS3z+xEfctyEWStkw8HM58losvhQMCcagq+AkUe
CDODJ67+9+65W9zGFL5NUvmoolEl3QkwJgpO8kLmADS0kBW2SUTDM6luElgk8IwtzYh/exWMRmY3
sIYMel6vTxtBUyew+dYjP8cUuiTxyaDyfYUes3EDyQGbFp9DFbHGDoLQDZItKTPpB+uGJnMriF1i
GEPQ9lv0nAjX4+K++5j6LeUUgg0wMD/j+qKQSLixQZ0PPua1HzTE2NDPGusRLhu5DUAJSFN0aYwY
3Y2wYiez4mBSTWi2bY+iVSrnAitlCjs3lA2xCozDAeehW1hmTENI9q1ajxLOYorrzL6oOJ1YCpMX
kKGO2x9j7MPg5UvErVx4Aw6YlBZtRUJt/p2bGfsB+tXVQZ6rRjyf8fcj7SM0PyAtFHv9Rjjp52S7
R+qgjAXHISTj8pwye42IoWrsqmMiH4kkD8aCNaScgjI1CD+x4bG9gLjxOcSm+MoIB3/1t9hb2+Rl
dVEs+MDtMBJEp6vDmy49F3WfrAFiyWqBcYv9LYrdT+0VUz0A3EkEaI0PY+rKX/qqekAmKHqMfzQg
e9P+Y2h90gKKAgTJ4XyGiqyrWkFdsxIVbCa9UdsS8d9TE5f9spdgXbifHwwo+600SDebQnCsBh1f
21970kX/271+FYmx4M7Au5dwg4dxclnxZJVY1W59VOQYgT68FtscM2HKKyaQzicynl6YcaBGcciG
ts1mmktgM4S0AkCYjblmAtrt9pGaLWudzEIkNAIamXguSrkvoTHr2XJfjquIevUKqK0afxufOQSJ
nXey/OM5BRAZDlWe0v/5JnGJHBjLfqiHTmnBNGouimqj6joGw4+pgAA4BPVx6wzoDhVCZ98JYgwF
dXzbcfJTpojaaC6ZklUfC8c7UNjR2ZSqeqtpKs04cNpQv26jK67ZsouHORX3iWuZztlq/dmRfd8c
IyWrFAJmWBSTwD9tfxoRWZN17xUZ216WEUGofoyuqMKHSzeT2xnF65hkJGUPZdI2RStplq8qY2mg
Pg69xquSueUzux/Bh+TGeacc3KbMPty4XnwnTCZx0TPt8MMZd/3/XZGFct6GKugjcRs8uVD5MgUp
JOjfPQVd5MUet53yOOOnamxB6FBODTJ7hT1J7BBqjVdGrBMPwTbfzFzMe+1Qvzw09A4Qqy0D9uHl
gfLQ5E/Noz4+mQT56vLMvqcRFZL4BicNE58pX84Xg9XtF4fP/41PrTa8BVcgUIrK6pjAHblPTmUi
vt35OsVE2BG3uNUnE2OpXGZFjHh/8aSNk4S9+vBh/LdN5e9mgi3UCKvFfaNy6EUx9QXVXHvraTUq
e+Hde2/8kHyPoi6wPiyQmTx6S+eD3a+9YpHPBZZtHU36XebSW4UwAVHsBriLkp/w19Tq4iS8EmRZ
UjThhFvs5W7IvLw7aNoxszzmV3L5t0FGQBfmdSf+nDLM8VbRVGE8Gr5xnEcR53dVf+MmuYWkqlyN
zWllvqioDmUOi0ZISvFUhOJjU0J6dqHMamqnLZjud9JFDrpDIQaQ8oZBpTLp+BF+WTrvw//CBVbp
BPtk+sWVWCEGh3p30i+tT4MRveCTE/AulugbHyad8maKPX77tsycIVjQp/nBuWonmSVhQsELxf9E
BJAcSQ/G4NR3rzfjjgcnqEvINCY3AZQv8go6tfA+u26g1sTGlwwQTd5ueKAaTsvY/Fd7qfC7yai5
m+Zwr068N1ZT7u1AKBdtQIL5GRH8iNUI/JjZDmMkYQEn7njWwx9hCsElfCp9GYgzyIzJ3yrP8fpW
bnt9Pk/Ox895PVLh1aEY7MOKY/T6vdR0/Ag1xXmR3EMAF6GV1kblLv9abyY5e65YytjA55LCF6BZ
jxDZd5uTk03ajjdSqSgLvyiev7jG2ZB37PGt/Scp1/XkLL8VQ2NdnsQ5fgua8j4MU90pYqK7hWGE
OvrIRXXKmnrTPnxsAai+911uSW/WH4lPSI5DaWki9NwAS916stQMrbeCqg/jjyJMmGNuTiiYbvW8
gtMTuzT2K/35aJ+obO9gYi/ktahM22WswjaPqbNd5sriD0vtyMPTkUI9DlgJDf++BO8Xdu/nbRcG
iVmVHZV35OKutnwIm2nk6e5Q/LHTMgKZETvcNdTNqu9uf7s2BQn5ihBdhwDi2M/FqVmN8eVXiE9X
+qLx2z+fmtma67ZKnaPc486AVSfq74QxDT+PogdFddg9mnuOcAAQutSJSQ6bXG9MtbZJRlPmb0cj
a5D3EidOMvyXV9gmpAi9Nm6hlrrUzgY2L8sdxB0BOhrtlXn1T6R8EiuykCEmHrk5TQkKe6hiM3x3
0RQugJco9iOR/lB8/YcjtCYtiN4qTsPbhLL14Ahp8q3Nn5EXKnnBiBTPVOlIplrFja/C0hsDqWnE
KWMdQEh7Oi8Serh3fFrScEOQ18OEV52Hki+3ZasrEVPqzfd36VzZTR+N3m2kNvbUs4abPfPlTe4p
M5y1r9hwGD8PNNamQiY3PnZbAytuYwfIeUlApbr4DAO18btIWXkuVbfZ9Ucq3w4JkswlLLAiJWLf
oEyHMBtE8bqSNUYlHwrb3HTsoEntk2xGNNZziS4Kw/qMsDa/eLpSgJZ3cjlieR9WBtcgdTBOsSNO
Ywt0jlNlZlfPRFbQOTCNCwZU4jXu5gfxd0opZ6zRfeVdK1smJi3hXr3c2LPkvsmPCSvJ2mKxJkIT
WPwQThOoYOMhYK60yiAhALXqxWiPlMkRw/k0TTYxp9tbaGBl/gk+lShI1CfXkisOv4yiBoiewm8j
c8USh6ZLU3Jfi+J07vxrLealRvax5TR2h4sKgX4RFoEa3nol/Bwd6LYAras7MynP+8ykusVTHi3e
wHmJdxELky5qRwtA6stvwBBYwz1z/fprnKWoY9NN2l6H2N6gYNl9A0WhNedSbszyjSsK+3bAWNum
JpSDcUgR9Xob4z2oEhKgxzRfUxnr8yxeW9YfkCoE/ZJWNEdk6XIH58TTgyHxSfexTBkYpq5N6f4t
iKeHz1lUCr5N+tly1muKupdqaLuceQaLlD9KlL777m1enb+YVKJI5vXcWczekLFFxiL1aqzx5Kly
slAjyBTpwb7RK/Oc33rZH3fTw7IB7tvz/PUnE8LahbiGptdudaSUfES81hX5hiNqc8gvrtFFltI6
cv5f+5OAxkTM/RkIJQNiHvqpWVTvZQsA4zEt0/kwPbyZoC8WG9HywjDh7flAqZB5jYWadXQqggaF
1L2RTFqkznowhyAggmhVOLKO2qKJOCImBJnukNM206lbTmF0gBbWgtWUf2uQTTH2gI9ftzJ5Fogv
kqlrUj1fsfxHfXrf/UbwMLlBHBg8JS/TqWykd5ts/hp3yWd20b0DNXQmqh9JNDoK61YeA4/fLUXX
KlaRbjofXZTU0/1ciUM/jE9u6QwwVsns3XJR12w0c47AZy6L4ok9pWQrqHegDUZgZVocrqGuZYOV
usnaN7ySLLAl5ARJdSz1en7jJpg7PBc9flBR0jaNetAhDr50kjS1ClxASfxhyeJpsm+xb4uenwBS
BvjLW2TAdFZwKaQ+WuRR6W1F3SIbnN02lbxAqNRIOaCrwxn/7cshSM0puQODDY+tQilD9wO2+wK+
RekxAUoHgwR2xoxYJYtCqRz8+AwMduvqgnYtUb44dyjwcjqzj8ZBU6KEdwoisK7ONqnA4GenMZQB
kIj5Kdik0p1+8bLhypLpug47TxiWVHxlwZ9iRMCkz7h0GTUOodb/RxqKhu12KcdadvAm4ffsewVx
5vyjCyn5SMOnwGVKWhZ34v35qiw63V9OJwVfaPxSS6zNWJeMt9louoHlKRWgmcV14tTOm53MyJBp
TVRNAxDeouwFU0Mhn+9lqFV8wzQpTAlw+fPAjt3PYPjymqjeYvHup6G8rK0c2VkOKFO6WL1eYJBe
3VQaYJWPd2KDIoK1iF9R6uheFViMPpzjaPLImUr9EKbbEOESPWYzNOQLMpXA36uQI+JjTNCl/nP9
zQwL2S0w52II9oaU+KfvaQ6aRySlVkBM7Gis0/8uKz0zZikucdKm8kic61PqrDRxzM65PrNtQan9
BEhzkwoetX6hwXEK2xGZLeXMoAexDaz8o1RZk/UXzMWG1mScVdEtu8I95rdHyCwGkoALdP/TTA+l
7St8pM3yfjOGRvk2DYs7Mr/E8vDZVTXyS9c4rji7AEeZ5CLSni+gV3dPLZWvAP9FPWqxk3pfSyUi
HhiOfMlyu+xMiCK899CfX4gp3DEnuE5Mmu0GMRIpsIK9mzT9MpUIwONN8+sYWU1YiJG871M9n7NU
pnTl6ENJcIO5/lCJt4LCLqnhn+oYhtLQfdA1US+1i/86Nfo7yXIu0iUn61GV9SJ8a4+BW/RR5ciA
0gzgsRalcI7inB8Rl6qSoIX2O8JALatm3pCS58cVeHqhp+jkYPS3Wk2dufW6NArgde8eXG2VUJ8N
vh1jsi5Xh8rCaq73INPo4rBafu96q92fsp76aH1HD18YZpQj8AoIj74697TeidkaoFkM4vlO2025
/8h+uKc/2jtcyT17OLNu33/lw4mujUYa3GdYxgbkswDlS1yZOcg2yDqUJqez6qIpea0BmTAxOdLl
kRFOrenxv3PLy/znrXLnH5buEXjq0Y3Li8JHamrbcoaR/0BHAC6q5NwRFQxwu3czE/OwoRZbkeOD
xXgNU+Ob20ZwEtHVmtc1jJMSCQc4OYkXZ0KrnaKFaVGFi0ng0BxgfAHn3pZIhETV2CzPZufdwvsl
exYegora713/4auxhCsmT/94bnW+a4McU8D8UFIRYvz6qB+vjqXsjOX4n+G79gPrnUDk/hkr5JYt
cnOzVjGBOZxPKH6Ymo3cgJnLBxKxWBAavaAQXTGjpd01M0UE+1ie5xWC6bkFbw10/dU1NzFJYUZR
esB4wmMw3XBE3jZVpNRY2DbflgVGD8JeTOOrS6COQF4lw7s2cEwJIpR75q+zZwxfkvZDirtFjA8L
PsQncVcdctEFtfDOfQTuxzj/SLU4c6byG6E+ve1YgbhPUiJ88yaLY8exxdVPipik03C9vRHgnjob
0OTq4e7/D7aSCnUfWfN/QmaW5WsGNxHcLW6iAk4M2dvWKZtUN+8TIwtbI8hA8t8clS754GrGj9tj
XfjSPagi2z6/tHMghd6UPvR8QPrkUo9iZrVsaQ1SNlY8L8ju5MoN6u2QPDvATIN+O3KYraS41iNT
ssBOpFRX8sxZKVTqu4AVxf7jlMH6U6aTIMm4vR8clHDfP+x/xIEiiWQnlPdrwOVqH2xvbwj7uORw
dcZA4zmHNHdjlYmeanObsAkKUSOAHzpvUgUiE//5N+33qCj8ThZwEbD4s+2P6efhhKNtL0X8wdMU
DgsS6QBWgGrTz8DZHexIndtkFvPiyJNDT5H0FYIQXz0pF+dcD544Qbw7gp+pRsHgPNbJ1byB6SCD
1m+bhFFF8CnNb1HmqZ1y5Y6L+kWh32AhGX2MtInjFdyfqiGTnnfE/zjlNZu7STrN/wfOxJB3dhP1
3BNdYU9qzd3jFSyFd4sVgI/rqmvvcjQIVCpeRR3cIjt5Ws+hDsZyVSLVYtda/zfHF9wg/JDMXqIh
CqeK217WWHx4puSEUnqUtJpDQql0+0V2QTOvvPT5Uiu+IVJXOWBVngFKfgKcEX3RV2Rhjxam8TEl
DJHj1fmMUXO71zpXwLJ9z6VHvg4GI4APT6lUxT5dG0nLgfYSRPqkp4qY9A08wCZRmr6pgm1AFA0Y
+Tzm6wiT8aFJavXHDo0BwzGNieyshehTtsxhPv38fTwEOW5Rat9oMP1JpH0eDa8tWLOU4VKCBwLd
vKlCugABk7N/mYkgCzgAJeNHdOXk9K/3yTq4/oWtLzgnNTbrsBEmws2UokCLzCqsTjnNz3CMim4M
hbcw9h54KcXeRAm+LS1HZpaxtHmn/ynELYLMo0VASzdgr3Arsp0U3zxuq9UJGOXtmkbFSHIGEFMO
gx8bH2BTE9FxiZuOnqCcrrMB/btzt9JM3fwe5Zpx76R4ypHLuYybAlvtVoqwSvkMQbafUgdULDFK
3oGvHK6VrsAZHRIvAb+PSLZ/Ajr07W2lTHWo3NM8Nudo+cSwAxiUqVsVSZ9mDff5xV1LPF5Jowmj
18j7fmi/PpSvig/ie9bKdFhS4Hm+gjjnzv7nSQOYDbh8rHkGgTx2/0jR3YDvjIwPXq0eV56SBKcZ
2CAYdZG4VgcngMuEKQuFHQt1AcEG34KMqgddCspxJOJwYdtOSXAGd4Dy2SS7RI5IUG+Yk/kcjlbZ
JRf5upE9XgFXGskd0I5tuCMULy5xKONtS5geh5fY1hSNcO7vD7YUnh7F7OcnyY1GU9YY4PDjJq/0
SrdSJXu3xxQ+M9smGxOxo1luH/ICClMMMKTl/VHUb+vsHyLwWqNOTA9URIqaBZ1QR1zpDOcBCEpm
gkuOaLka160VgUF5LQjFki5kabQagQznULWp9mRIpZ4J/8GHx9Ov0Xhe18ADnNJQO4jtP3brPL3k
iDtfOHMRs42TD1p/dJMNGOB6LfHEQuj/UEJ3PX0O11nfir8S98aw/LcJwLs0USzblrMFCxc7mtrE
b6ETt608WCFC5tHHgATwwswpNLH7+71IO2lVJ7YfmWCugzRFw9zOqxUgZhZqvaimZaoh6ylsPmjP
2Yb400o6BZLL7rQQm/enCQc1PjOgJEQDz5krrF3IEFtlm8r7h+U71mK+CzHrfYAwwwajgbo/aGLD
0yGIB25641NLdR82WSY/eQBWQUkHr9TgQ/sqUVyfNms9JdfXrlk0TMDsgYEjEXMcHqcsZEa+QFIa
r0R/4Zrb2NAoLA87TEkC6DHlQzphFOk7iSmzvhJYTyRhU+fMQpfgEWvSzLZnCJIhC3Yz/s4Ny60G
W/RxCsGHhdzqYD+ZW1E3gi3c+4w1x+88NrAmwrNqbBH9p2vMAUKrYIpAJkpjB4ipLjBMid7hqVZb
Rkk/KMVMh20xNc/KeM7A0RWzAy3OvMIk0Xaiqv9ypopVtAKWHQVDYgYzRO0ppTzo0Los+gEG2T1C
VsplRbhf0vwlgi+dPqjwjGx6Nqid5D081+V+7dSLCTrT9rbLozt5ilMY+xTW4RT/HJTxoIYdMhk/
xvPqSiqyl5poQRZtHBNnTnSeDJf6M+i9EMI31qjZLY9jnIzQurjM8BohG6eKTnSeGISDtCW0VoAK
pa36hD6H1znFM/lzjSryw0dThi0cO4rQ61jberztebAzD/JeoswZfWIlLxPvd4FbGo0TWonn51uo
kArRcXwtHCRQYIe92C4YIFBJvbSN6zVDbMB3NiwoRZISUKKbROl6iIIU8WwHB0kz+o71doCoPRiy
d7vAoh6I2FrOhFjbqJqNOWjKZ78iumRLNPG0RFJ1BgUuq5BNFZDpPN+egpQZYL3C0h6aC6Jta19V
zKgUo+f7VkJty+jM40mMRwaj+jGB7uDjF0tTkTDbUGvFTrG87OAXsBwksUvsf05kPovWJ3U/pJ3A
eeSg/hDCv5mGFy/01EaXb7G60hF7vIdoYOWjMsFoZBcdB66Q4Z9D0hYxW1jwerdQW0n3/qWPAVWm
3GFBdm3O4eGnug5efRHRMFwQP/TFCzUkj6iAXO8eU7pdB2PDkgzqZ1hSv8Bq3lf9pDeRCDYX+qw6
7z6vLGak57p+8IC4hZALU/Id+WM8XvztEbqBDMD3SREESlgQUaYu50u3xnTixh70FfGxUFvkctAE
kWMe8NfoGKSWY++jIudyV9wiiLwaLN84xxglSIvFv+ISAL1xbn2WUjnTAsfqJgcmasjxOd7DrWFo
YKZ91ci2KO9lzUXYf+JSDpZndiAK+YN+nshi55OsHdaBWmHGwVAC/GUgA7hIBOmOMMWGzwCe13pj
G/7nVZkUinBIJbr6I84PykiQDG9pYjm36X52b1T5uoRTAkTlMaxGWVdvnGbX+Ucme9vN9Dhs1anE
B4NUuIT+KhfILh0IFSm7DXJFmP49+hWHCHWZqIqVxxh+Qjr74E0Tt6KPkn14c1PBsqfNAdc743vI
IPFoCtMoBJTuyBK5VxRKw4s/SytNhNWAJaBKdsxnQUt0nkPLkMheZWn0d3OyElAwXEwB2oGyJdDb
skQIQPEXgLXGjF6+8fP5+EJHMflSmiFDD0dzMPr9qmWEEXVKiCIggqrZVNkIA8qcFyG7R6RDmoWd
NG4Zb56Tw29meaoYS+UJ19D0srx6+oMaLKyopwDwojNvRcrA+EWVS8TGyABtRS3GTH9kUYjlDQIv
8YMwndOsBoB4aa50KAj/HUFQ5y+V5Trh9OCEAQo8lEA+onDDo0f9RIpqX82IiydZ/iUljjU329CR
M/s6PSHT2jQPJeh0m3AgXHUtC5orFQK8TtN8vReePmGwBZjz9sv3VxhrGNS0Ps8IY614Go/3xn4v
WJgF+K15N1pUUZSCwAQC2PmFzXnxjJ5G2VNIQcOUCovQLFyBry00XCkuFiZRatm/Ik7wLJN5Tyhz
1zW2rj5X0l1ByiNWHoQ9iz35lrL17bkTBWagMjcisgmWYMK4OMLmfCltgQz0jOkzCMmLU7StTfVT
2JXJ7OMemJyU98+33J0FAADnF7IcidSpxKxG0c5xvnII0Wqor+c6WRDe4djOTxmGTEncVCzfTx+V
S6EXW0h1d44n3gkh4jl76tEYRZUUENASys9ak3CxBrrjk+h014gvx9F9JV1vXZbLEoLZkCWbyeRH
QfS/7/ioUqJsJp3zaZqnSRzQejrMfiYhpyFL0/jkKY8JOrjbeJ/vzKK0qvww2HVxTCc+MHA7Lydq
D3d495sAg5UXjaF+gNCHMGpInlhDxRa3gnFhvokUQ7LOX3K8z2CU7Q9vUDjVgi7GyExUHtnRjgdv
DHBXSnI9ttqHSxrQTOzhWQR5HPYAYoPsdsyHSyLvUknuXF26xNklhFrRae/43lBIalzQebSCL+2p
XfTfz0unyTzMDmkD6ObpFjeGg6j0+gmZ0FSGRPi/ZSAghPO8TCG6H/FgyjjrDDmukJM8GGq4EkeI
ivtap9Yqkv3Gbr67JAqe0crmW70SIpSpGu1Uve64g7O4/a9smOarBbJc4eVMoAuWcoLGTB3H+GUi
KS3kE4j/4Gf3Nu2hODHi7oI/nYgaBUzkjoePgrYCFZ4PsUyRlk1D2hWlH7XbeJM6LZhquiWVL4CY
DbqM+sOMd1pFw4EdFezNUX/7wF4NqHsSmvUcQPdB9v4/r2RGUaSNV+DvXgjSy+y3gTA8OXh0eZZg
0tfsSDbIIz3YHcrSvpt9TAYh+S6YTK1U+IOs7O736YVJYDlLwSjJM/HpZqJYSxyp6DJmgbAKKihc
2pDPmAX7Ll2iTQQxZV5JSOst4Fw0oR5mxzGhyVNZ6z7pmm60eYkkyG/T0NwqpvhQjFbrufEhsWN8
KxFnieNH91YHxq6+0gR3SZtZ8O/Ec/ogAFfBTxkLHcrbCad5V006tz1I4lbLoTaWY3hDRgeHUc9y
hJWZ4zwQ4ZACOSL2BtSdeV4qp8SDWfY1eJT7mpsWZCEG9eB0dSQR2u5raSWlnO3FTdWpTfyBPPnQ
SU73HxlSMIIidBOYp4QSGOICBGIHiEm41iVlTXWfuat7cZS+/rtXqtHJDodME8DaJjRziXLSojLY
wxEDbcfItdMXxlz6MWw96anesYF5PYR+jlHCOm7Y1c1nFlxtX0D0e+morvupyT/wKxN7eFbt6Bcu
YFJiUv5la4Iif6O6ixxlwR/4RYtsU9Fqt/H1e2xmw0fqKwD1tibVLCQmu3p+pdnaIH8XTVVP7xb+
t0TPRM02+klpFrCFEe9DlOg8H4SbL52u1O52n6e5O7ymPyzFVJN6Rs5LSxgFTZ3nLwrrQ5aUP3fZ
jTQnQ68YdLFFBIB0O9y2p0lY4+MkIOrBWmYIo0JuuZlhVzQAbu9RYD6TehBvvit21+OwRTegb/nb
Ot6oL13HfBW2tNX6RITs4gEEz+r4IHqJgJFWKIXTu3t0gel+X7UXYkZ55UNIRdTrsyDUy971pYgc
P+x2y+5SciWoNcusg7/vB/ASMLWJB7hW1hwAr//14ZQajvl1gX8d16OZRIfpYwIUiOEWJay6Eqn9
coNksxElrYvfGsUFWAU2nfUmXOSR5jBNMWBkBarEQ73Dcwy9kfC+8Md6tqO1ivBfYlgwslXBSzr0
TEYVDTb8GDW7HTOy7p0CwF8v5Fl+ZrlLKUXRUGSNG5AMrBb+1U5YsMojsGbJVz95wHrTgocch4Ab
bSAcbgV25KCLPobdCNBwnos6WXSVet/GfwTaMAovRaLEdih2DozlYb3WZ4wFanDkdItq18qnCpg4
mXthle6JjR+d2a6KcNqP2Mc+r1TIQaLThgkwwdlg4F8Su6cFEdspMHuuFG7X19MgN34EFg7Mmn1k
bQ3DKH37aHjWHR4Skk3vyfS8ajpyRynmpstwe0J8DzXv9ABLvCmJWj/Y0rw0zc3mIMpS7mBskBI0
8l+cN00+jqu20yENd4NA7H+SG1Q4osKd3bPpH7bO/3j4+y35Ejtl457hhvS0eADSxF4n02vbt3DH
EyKH7H7TgHBCuaLxp5liTFz7w9Tlg6PGLnVN6inzgBrBgN+bAM/PzPRGMTtOi2qkcL/t2TTyzNRJ
OSUKbeut+tbBmV95uBXurw1lYPxpLco+YNYj9ktr4U86mxj2uMM1OtrmZInx2pchmlSSmIUH5Ogl
RKsczi0mJhJNDWRekj7BXhcez8dIEmkjJ2X56gV2Xh7NvGbvz9tqXYPSXeiVgbwSEG27WjUmJ/uD
X0eJKUrWcwxFOsNvCHq6OZo+NbpoNx8CeYwXjP/hueWzlCo21UeEZu13GH6KNBjqzdejyQAMpJtQ
eDoUXbAPNN/Yim3XL/eNDH4UPBssLQZ63N0CWuDv8Qq9bJMrHBBqNVVudk9ohRedvmb5Tae/HwPb
3q74d/MookS7Io3rtJg/wrFTrAQw2Py3QZ0GbVn+0is8hrz1IVJRhnFgG8AZ7ICnhiKb0bBwdnxP
+1LjVZ0BUEBc7xW1/0jlnkNXSOugJHNDrLQFC31jBHlAGFHckz9hNlHxTitOHiFh3uQNSF2dAnwv
aFRnz6QOgXbhSBmmmxvbVKtLduwrkoqK09WiTdCf6luUEKA223VErIuvH7Hk9KvR1f8KOo/lCGdE
X9JrzJGSVhPCr9LgW1z7hx5v1UCWL0zHGwKKVufGcijE8HAGwyAouDqT7JzR2Q5wezsWpTeZ8Nnv
JpPnsuIjpeHEPzJsd+JdGq83HVbVO6rJbBmC31/k4HmwBS0CVPlVRPGVo9+5IA924fH21uQIocgp
wImU4VyMp7gGuyqZbite1x6uZcGtIfjueimhQE6MpZJcBVpz3N6II01iXlg6dt5ZQihMCevoQcaF
38ihHwurFampEsTp/b/kIIRGnw4HSk+WJ4VCZ1ZJxygp/iyU2nnukejEbuE2MRYrqNGUuOauOjgo
KB5ikTDZ54/0cL9szPsdECAdKZDwenvIPBPVXD0T9nMRlzEXWFmFQB4A4BkAa155JduyrcBE0BQF
zB8PIYJRWjRfSsQKmd27L0rQLPCFghtcTuZQGpLBbqXUY11DxbVlplLXk2v8m7sdxRVXx6v3zcPl
Ns0/NtJ4cacD8ZY9Q8gxwlscvUT16FQRQg3kMwIqUPGuUzeoHSaAaGTtS1bHZ5GLqNEZHf6XJWMK
gKjI/NY3TAd4LmfwCxajEzHHNu+hzvNepopGg0MGElyJFo7J9plf5LsqHY1A9z0MGm1oT9VIacUN
imT6DW1BnxhK2lXbQLyYa831fkq1ZWGS6QZJ2XMmV4ZOkGsmDtdZeIAY76CkYtCzIcBLEAqi39c9
FyYDiZc02tb1jw5xoNKag/T+PknCPUwurryUR8EnnH2Gej2N7tV4S0L6Z7T/y0J3V6t8ow7q4OtN
v9id3HW1DcMfHLiXAwPnEmQ+wPVJIaXNnx9OrTJk/wxTvM//3B/0HM1W4X7u4wDf0bIMrBrHS9th
yDwIJzFCAzIcgCO2GWOoNhsHsebQtEtiLf0yNE6ULQKgpU+QrfuZoLn2tTmsnkLsAwsPtp2vZO9a
6dPKGO+JKqBhrPHxja0WLuTGrIvy4wgaY+LFM2h0dv43SYPSw/A7/EI9HWfzTb/zTJpQRZ+IRrTM
KGBqFNc+6MONlI6epx9sjYU0ZA1iaQsPAbhqUp1PAnwtbIjDev5hnptPasUZBHHUQ1j+CcwdbNfr
TFAC33azkpoAR9GGPj6bhwel0QvAdiN+VhbmhrZTRfnt+8TxBzEco6an2dhJoA1u/FavFTh+/YoC
j+VbFtJJDXIIq73g0SyScz7W1qo9OiDQ0b85pEzoaJZuPNta6iaXssoymPvSFABHHlQ+E2MkpiK3
5L16NcUaFX/wbvzug/BUHLIB1YBGKyXFb1k4nJb2M6qWrHAwWxosssYdvYPwVXTD5JW+NPkmcwZC
2adly+07LAbEvfIGHuAPf4eLGN/aSTneIvEdZWm1R4iUb2JBmRqC1PvNILCVqwNcsJiLq7+zO2K/
Gzf/+0Uj9ny3aFG4PHjTjMLss0x4xa/3gSNVGqHZfs0Wb4ui+UAIA6u8PUkiz8k4+hCBK0LKN01s
SJNMgblXdMItrJNO5BsBu+NErEyuGhyLxLg7t+OFpjXnrOVn7I1k3yczhuYukT/v3ygHGzl9u3dO
ly9nFnL6HL5ixPKfHLX8H5+K/ELhoqfLlBFBNMRyluWslgu3lweM0cQ/lEE0WpsuVVlJpI6GAbzo
KlfeJE47IjigZb/yLmB/jWk90GxhMmM9Vx0aXAnH+7r9R4er8xb5AlNI8XBqaGu5PM0u9kVYhZaf
B1ltc54eT1xrFXMPZ+6Lqj3nrr+8M9q351Yw9yYz3jq9wt03DOsCeD5HQVjLmJFke/FsAfkayTsw
skXIOgxuRE1nRK8EUvQd63HJ6Hyd0inISLGvfYeS6NuLyufzlo8t/BcqtWrXWxTIWfCq/zMDq0ar
tKcMql7+vwcicEaq/YOxIsGKrxMrZkMQmnRZJF9PiIuy9p7HTZDkk61q+17huKRjFEpKUnzePO7Z
F5fRC4gg6Bow9alhYN/LTHglWLDC4fCxRYxmP3EKl+VC/t4UXf+yh12zDFjniutwXnsRYFFgU+wz
HabQHLtsVh/NmUUk/MvDytUBYd2F/BvxD1cY8RcxZpIXm66Sj3poHAfz8AS5Ybxbro1j7MKSsjH3
Q1vfcPkiJwfN4Bi14kVgkXmkz2DtOapS13iOQ4ey6cD3XZdGq8/rdu+JYLXCipthaC2l6+CpZolH
qhbcuc+GSZRs4S7SiBlnmIYH2DrJbYOooXBSaPKvtZqatPuuoTC1JJAtySqaM+tidpcRRNaK368A
hFi86pPQTZBTd/2MSWDd+Ut23C+91eE9uJJPOpLlLqz8F5/F185kEiFDNcr/+ncaMug0Z/0ZwxBD
uMCeqiGRQieH5NOSWFQFgFCUo4A9fkdOlUoPe9M7JxPwBiJbDEFo+9YIIdUaQGghbNoHI3ic6qAO
GmSdx7hSXrH3HYwruC4VzkfsEbUFdE6NdJbmfbbUUy91ng5/Tw1KwTyFRIqHxkcpNo5ZhZpC54YR
0e8YMC4myv1sb+MTwHPNxIJ0ByDEDtI5ECTOjZaHW/t0PfFH//+fLttqB+BV8NHl0AUgVd8hEp93
D3tLnncNF79KAu91YO1qhK914WC5Oh/d2c1RMOkwncpU1JZSf8EVKJKylFcd4x2gm3s4Cv/yltF9
Z4fRRK3IZohghtT2kW7K2HOEi7s1dmH1U+7qxSD1j20zgfoM2nUr4oMU9Z9K5BYJNIfVYGMMcAv3
NCjxQ5Bit0L1JO23S+QIhMCQwnDa8+k7qj6GWkMtESPQ0njciJHnbbNwSm/UtG/i3Btk7JNCoYSQ
DfuUqB4KasFQAO8BLMdU9DWgaxcUAaYmwrnroqek59NIPEwWgspZmJ2XGP9+HJU5O/udti+5Iwo1
+HfIT88Z+PTkQ9bIK9Kv2cHBR2mlOk0wb3Bwkh2kLM/2A2HsCS5mJhFlYIoU6J0r5m1KV4ogb6YQ
eSEf8i3oozYVaNZPKCiXYqtDP+EhLIPAyrmM8c9pGJyppRdgx3uxsHq8p9Yd7iddusNTRukLLC1f
RctexNs1oiELPj1mPVSVe+itMwvtk1dwrqqJfxMc+HaJ+DgFeFksgIp4pV76WYddkchjnUeToHWu
eOlghAf6DZ4yyxrUeMZNBC4oJ0i/I582vtCNv/exVmSNHNcAZzmJcEU/VXoh+Boy8tJDH6PSLlxh
CobmjRX7/v0EDZVNlB8qfgaJRoQi9l0HQ0xqz2LVt9PsiXs8u0PX9qoH8NfINwfbsPjIzXw2iZ5L
KGowy3gG9sa5dQDl1tZq5M8LmjN4R5ytYe4hWewk36cFbOHLdauM3p/g9ReZ5s+aiKmu8xKWA7eN
E/dSP+3SdC9Z7VRW+ar5CKgFhqIqBzjowv1/Q3bcs4rW4DgUfAfDPJ+SWuSMgzoByS+0wlNcBEK3
nbfNE/GS69QctnazvO2k8fR/t+WO9RLnHlrCEBlRxKIOk8a9lXbfCwvzKvNf6hawHAsYlgF+/JQ/
uR43drLJ0MgQNB055QIspPHlpKb6nMCwo35jmru+HOEhV9r2c6NchLDrgOdIWq21dUcgCseui4bc
uqJHGgFeTvv3FRGuQ9ClPhfOOMaqH2H64Gj6VH+PLXOJQ4KlNSoJ2z0zYA8xNiuK4h6qYqYuckhb
NUKY9mSquu1AILSHlIxqEDiN1to/yVuM0LLOOEr2CZfY1DwzF7fQsz3lXXh9Qid0PKi/QDq70ad9
0z1s3aAxh2GWSNBC2H7BCLYKkAebwusHhPy8HG+7Vw2nZTQDoZoHUQ9xaZgPBj/wFQ/mzqAb2AKb
WK4xIOnONfNXMbYXVRNVQidOvpfuwcSVvk1TpLjU+idXK/Wv4BilFRVTg2bC2o8L2vWPQNROcemV
6AmQYPdbaFbVftLzuaHBxD/Y9Ni4SRIM+9UKDpcjJ6sv8f7ivIX3nAPXs3C03rMmyOqtASfXLTEY
hf2+J8pt2o2TwUKpZWnXeFNEICIX3R5SpvwkTBSeAE5yNJFwuuTmRRRVMeux4W7fnCV4xnAgmyLW
4S/kEIxHDRw3StnGBzyylHlPyL5E7vgog6y69/Hg0nktr2b+ItODcBrz4k91CeYxJ5Atx7+AFNRm
FYgHdsZtmF4Y3kRw2RlsoT+esQPPh6w0w2KZ4GcrLsPlllHjwMWB77BVgwJuBHKaFtRaXCAC9/hU
YGWmPe3Nman9bw84yj+YD6g7FGURF/lArVOhrFe6d16fUTnnfsoOmyDf2Xkn0+UCNFI8Ra4C4ib5
tDgD+1h3eh0AFfWalYf3DjQCuQD+K19c37f06vqFKNad2X4tzWBya+/1ZPjjSucJ3sxvbRu22K/F
72VhCpVrssr0x9w+8iu13XbdOguxgRq5b0QTGesfyZcelcScnTNYCSkEofk6kdUE1pfRV4Qx6MNf
Tv3VqC/31T7KMaKHvzv3X0MG3uyvCJd2erR+E1cU1xRcq9crhJP5Bu6qKIcyVgXA7yXq/hIvodeC
of1j8bhRv30ApzLMJ8xnfxRgOzXSnDCpeZm1V0i7U1x34VwR+9Ca4YfiyfwOPwACQXr0ByOSgqFH
AOnyRdMNkxjHZyFNx4bVQbks1ntwdNATuuE0MLM0Ca/SxPxw5d6Kug3TKa2MI1rX4pMFA5ust+mC
49mBGOUdcbWE4Bxh84ZvpvysDuf2sQYC4cabYepoNVQxxb/P7dISvUlBwqEl9ts14RyBWpC9in0C
I+hG1UuUZlfLGCjbaN2PVcGN5g/R7PwJ1jQbbJ7ifw0VU3jx9zi/uIGP5/wrC6WdFEaj/vpk/RwF
KV4eqCei2cxUjFiO4SYN8Wmi2QVmYWsBpQhA5a/AZelg4aGVMQlE4o8ZM3315WpLdtDV7D8KhH9N
45DLubG+8rbNR7RBTpcRS8TkQAVy0Pmld+Ysf0Pi2+wmgP/vlqymmK7oW02Ry1gEzG1aiA+zLmrt
VqaMQh1gjsBsJfmsgaHRTUtX3VkqGTctsbca3wNhEs348HZilT3rf0kW8lSXWAVE4RqY+dMdolMo
i3C0Ctr+B4zGLdTAqTjh7hpw9i0jMEr7uVEv9cs7+WmASp2o6ZtuCyGVrhCFwlZlbmC6bu0Eh136
QQct9qPiNWbOAa3BI4Zu//b+/c84GqADBXZDGFaM7HfYwK1sO1x88EtkFNORHFtggvCXD7Gt/8Sq
yRcoRgj3pynOTVUlAStnBvKMLpov5uvJAHcpKN4hXHindboVjLVycOyRta0c9WS0CeDaCAMygL+v
XzNpeDzPv9AslmlphNTik43FX5OttGtbuX/KF+UMAcYiJnjvXkW/cSJyuAIiQEhqcHDpC7yTLoUX
8Yh336fyalcUibfHjP+LVuSBjMM5p7TGRvyWnVANOL9pCmzsrHZKMZl4p5qLLstt7Vr6InYn4X0J
YyrIH1K7uIEgvJJRh9f5TWs2LDW0gVjZN38uJ36ONvW6p5heOk4R6kgKZRCXrajoFZ9tjnprUI+E
1u4GQbnA+mR5czUTEiVT/9gwJ2vYq3F66jhWm75hTHh0ZVfT86d9/hA+crZkoYKJCiXQgVqjTsHE
gayiLyBMHhJh+HInkLPoev8oerI0t7tK100IPg7EF95rAWPT6uOspCX9Kdu9kUUoBB8U1QHpYeKm
ZPbRN4BZhg6eZ1gLGA0XFYE8BHlk0UW7XEFnGLeAgpf6eFxLRZJDtRaS2gPwRS24xQzlusMdiwLP
+viZ+BY5oW91N+6ZugfWDwhF3rwGxIIRTVKF25HzrUbeCCt323Yy++0GAcCjgKRH2lMUPkHkvyay
O9SYzf3OIK5ke27zzMPvWQdp2prb/BnF/E616dIKiCpBx9fPzH4AIEoyU6iBrI7GQchg91LLBOyM
LnDX+S+b+bjY8f0elSBn92stPc/hpdsef2yR1zL5U6xwLb+071M5/Bk0MnwitmP579n90wR/fgwX
YnJhywO+UADURqLlIKRkdfdDzLGF66lkvuTV8M/RSoH6XZQxZOoH9ZBgmnb0+lSMwcAvrBfAWxnt
NVm27eDTE/WfggJO6xnTjMQMFJ3gF8OnK8ywMihoBcCFJG5acrldEAJ8fcezUXdx+r2c7J9ONcOs
ezxFt7LLr8N9RPvVZXgrpbgHDPBmZI0KSwEzO7r4aPkJaExhYNzx25sqr481Cam1LxajWeKxUG4Q
3qBnCSOorzrA1B5w9QMgv9gHX3Vg6Dw/tkh8Xgwe50LDMTdu0zyDUPFQZ7VdWXXkZ+kz9hFCVotv
6pvAakX5i61iyDfKRQPpIL8UGdhOm29GXKEYRsMBihex1kGji26fzQuT6JDTQeEFum01KmJHNWfh
WBMlqyqFQcdvQ/Z9KWgDFyZ0SsS9cympm/5twsIcCOmQXAQc/7edyYpZ9hQ+WxzcOeN4tfiYV+Tz
aFBz8QhcRvSalI3W8Par1mWr9IeXHhl1/LXuRVR7+isAaQR0NQELljdBlK1Mywfc2iCAJfiPIhkC
JbWoZjgLgBijQiui2UCDnbcVt4uqZTOHoI1cxdwsTIX/HQyRL3/yhoW8HfH5yEgn+geP9/SkGRnq
UEjz2BQyon20VPElX5Eku1Drnn26DxLzMVZCK0gdS/PZ0YFh6lQuD/vgnyGVs+uZEnU90ogkbM//
QfnOKjT0sJpsZ8x7VPWHnraFIp/4940i57hEZTt73bt9Vh0b0WUSrEz9b8EfcuJmJgRGQklV5KqN
2zkfDi3VFbCSj0oep4CZg7kB9IZ/LUM6/DsRlMOTaHF5x8VRnRxw7wt8yT2x/wwBQkCmkmzlNDdt
vTuTK2DtBBgmOhPgnhUwY+chp21RAgg4Twgf8R+3lA1nMYhWDJM8UqLNmYCqKChO0MBpQu9WTu24
XtPwV/uq+1eNhzgo/RdSfNmxbvoWC1i5N8wxfYV65QgaEV5+VjjKO6zIbYZ0nRzKW4OpHQgJ0FIf
/gKtmIOEE03bfNGidwADdgBQAjaOQwTw6U7MmiQcHuh6vfcCeTV710Rt2ibsAdmi15A7pDRjKIFQ
VuISS7BCK2cVrig/7zgp/hmCq+EFpUEpJKfVx/GmrSCuhQKFTh0MIM5FdrxsdF09Nkun5OWJ+y5g
Ps0M0njjU2QxUY8ETwHsQ173MHQXOxOqr7OSnkcw2IVpFQjTMlU19uM84r8SpW+YpVl/r8QEHz0L
IwBogLF1Vq229thrKW0QKLg+eNjSAHSdLUy0+4S9l3YxMncXkXITVD4uCO1qviJALHwkgVPP569v
aMCpo9d97UTtxjnUfT7RK5VvH1cq5IKRfKFh7k/Dnz6eY3afJvEgPfutNUU0Bkdu9gYA7VYYTMv+
EQWwNtVWdbwAC+qBww4rIEhOgZpoh59URZOl2k/rV7yOxgVNVHeNI3Dh8Y1MX4C4QmzEjExB0Ri3
p1V5/FMlQSNZbwhOSok3lVzpL7ufV7i4TV+TZ72/VS7wuGijqUkOFSJXVxFjpk8rrQ8kH+JjfSKs
sAyNprz+MdFa0QcZ531XWZxyfybzhwlGvWOpUZfMfW0T58f8Ngyidyc1ZjMhb4DG9qOe+Oe7ef/S
5P60x0b4idfluyLpBYfFyqphuTOTc3QRVKGLTBoTrTs3UoQpxDkQ3qj/zb/H49b5krbzF8K0eDJT
5a6NbWdrxXBCFUaGgclBnsz23YhOKstjMQIjiVZam8Xr2xRdI/Z4NS24pZF1K+h4v+8W0xPji52c
ck5SZ9KVpJI+ivIwyRd+pOc5yHS5LV6ablZmyL6PYmaqNHqlyRZ6JEeaURIwM7ewqenjPRC1frGh
XPlbJSaB8mlGPyC7A/4R2cndylB3t3OACLkrSUEN3wxjOPD7BNNrKtUmFjMPnmFWaO/2FQQ10cP7
dZRe16+fuw7N4ycFmzzRKtQTHjEjReTZlewjvr0gn0qWDqqeOCp+vmmrIfH3Al3LPxOC76lLtH3g
+FccjiV9YVyPSUUM5O5wvQiqxTgj0j5ATVXD41uCUQXUKay+aj+G2mtGI5UItVkPc/9bwr75Xae6
9fpsUN/Yt6Lvf4vvFzYdd4Qx6UePUdInDhNqujbPcXrZ82YuK375qpepvW/85Qh48RqSwkE6xA3b
f4Bn+kg/x2Ntk0nIRtgcKCXNnpo42JqTJneTxDkX1MR/vQKiMiXdqlJeYTYBw0dqG9qXPb2sGwOg
TxKYJN7htOfnXi5LyUrC3QYH9hm3z1jebtYWSsy5o00BOSBARP86NDYeFtaTckT5kDoEtmZdbGY9
zeevfaF6xqsVsA7ZUlWxk4Vw+Z1tyK5KTdkop+RQoLHiRbBtUVfdb4HutglB0heczckTv6VlvYnj
da62Ovm1oZW+uU6iA6iJj9tXOctb5D3ofNQqr3dKkQw1AFZLGniNYybFDrSoUHoe6AZCqf1dQQrE
CPxTsS1RNWXpTCTyg2rN6JWn79RnrV3Yc8pRvduM4EmXy50s2JbIg+GGYyEQkXl397uDxZCjzzqN
CLs7WFGvdZqK4oduFdAUK7ivrfJhyct6ne1LPLUDRo/pCYSNkb/gbKmEYjzIU3wGSvuiPEZwqtB+
AzLlgulsABWBW9BIL1ozGXuuITRgssTSot3mOEzUdTpVAW3kSb0lGlnAhBfX1DwTPZXH7DdnbCbT
1kq2tRfaTO3/VvpVEBZ6PbayYuB3HTvaHiwdBEy9UpHuCd36x40zIuD5tKToH6WCzaELaCjpQXxk
eqTyNXy73p8FnIWKr0VCe2g+k6LombNs7b427gGnqUyknHY9qLmqG2xU9mngE6Aw+qv0B6I8wLE1
vfGPcAdxVP574JtzjtebcgEE/6o4xoS/KpRSJgjJzojsFjG93eEav7+M8s5WsQrNTLdv5NO2adfe
GHAizYr3UQx2agB9xd58HXZjyLBQGHAJg1GdIcW+Bfe9tjzqOKXGmnxDo7TtvzujUfxtJnCCYEbD
AoNw8vT3qIKnRKAP7/L+1ODNL/e0HJiF4Wc1HWkEhYSniD6XIfwCzI+JUD4B3cGqLMlWRPr7qpR5
Ypje5jihq5sZICa1GqyT37l27jEkwqLahTI/TJRj+0IQ0PSkdfL/U2VECoc8VgsnFmplnms/M4G2
RIe2gp+rlLU22I/s4YhHUwhWZdhJl9fFDahNA/A/ly31OhZ5h6xavAxp2Sm4Xjdfow4ZWgmKfRUC
Z6WXiqdFIdf92HqFHhw+OCMronxI0iVQJB5hjAv6Y3ugJgd4NOgidzdgrNlUQPizg0NmkxCpVlYA
5FJLJZgVvQstTEnBlMhFHp/bT9OwUdVpNzMLTBrG37l939JaZ8gFM+aO6mUJjZHHufH2tI5v5FKA
VykgDTq7Bo5FWCpXTc1EXpvBC0plsvaah+Fvg4D3StxqdagyO/9a74Elt8ol9WYY7hlttuBwJat0
0W8hsmVAMtlBV6fuWkKwljosVcOyKEX5C5AenPxfI9EbL3qhc3PfYtbKi68Mw8PXSvxvL0VZjO1t
zJsMT4pDTK3lWg8Mh7T9fHhUc9HkJKUP+4Axu5dl603FguBkCO0r5+2pIAIwbwynjBm1mDP3zjCY
ZJjs/otHuoRfDCEuR6Aju1X4dtqE2tintVcNseyN5lvO6dl+8fMFdsLZVJryKJz7yZFI9TkkMG5p
Ecq8qgDJb55p1q6+Bl0gSx3hDc2ytIa79pioF9TldL4a5L2d53t0iuj1+HaNi05cNsDblsq7FeOZ
88MeyRRIPOtbe7BxdSzsanQs6/vkPjXS+XOsz0g2I7Xt0K+eNfhHO2iYUQS17WhlVsKMDBL0e8g2
r8eL/kgwqG9XYzqr3JMqtiLBEUpHVcr4/ireHJYluy88hQapb2EI0Bdh/3sOBqIs62g3u+/ApBqO
uWFvKFwcgOmuznpdMc6/O5SbYwghUTRPfUTTr/1fZ3xi9n1FmDtu+vQP1eumujeYP2QemPQ+IVES
sHAUG2lVA0oVeA/9yxfAp1IHJEXDDUjQ8akcVKCBwO4IQJzGPAZycpgoVjvXXzLWF+V6g2MgbaTO
Z+gAx71MkCHu1tAyafTlZZk/mDvKfT2D5rGuwF9bbKhhebildM/Dy+NHYEyOULhD8a2cOgfUOaed
3uW8llDtn6jDb67SsGj/3G93c6DQ7k22KzKPlzHVJFDePll1uKawmHB9hh7Qrt+cz8pSsP9fc9tl
oyW1sRVQKL3K0+UYQwmFHqZj+P39GmRAXEMjDd2xQfB/Eb4bpN9Q2OIr0cH8wfuNGBM3ELiH7sC+
ko2j+xalSZ5vctrMfzpJwHKcNKX8jQkIbbqM2CMbH8wDNW6CFGVjZh8Rq7W2hLace/2DOa4Suzbe
Z28sSUM/OXUeqZxE/f0/rJjC1f9WzVejgyjXk7NNFoqMV/HWACDRZuKxGbP12sstItWTfiki7IEw
qjrm7gA2ThFgR81M54VFaiU75qkXgtGFW5a9YY/PmlErlVEIaHJQS773MOqHavDkIo8K4A6i9O6x
xNqRmtlhChPBiPSjUJQVxTnDPdP0Z/UY4cpsDW5Tz/a1S2uQjZnvwfCPUvtoDZVlwhhxrLxdujtG
kYq7/JYNeHYmu6SZX791GNR6N5GKkuLhR0Ygt5kdVVtMaU9ecczSGOE70a75OQynKd1KPDYBMj/2
F6WFC+y5t33qfJmLYOcb08XB5c9T6Q9mvdxun5ot2/TNDK/giQDydh1cBt72jaO3Wulgtfj5Yr2v
JDXn/qN5moHYd3FJc3hFb/Dqa475eFwXk3EPdT26Mt/p16AP72oejS16PNodCKMgBmiBNbKlnrA2
2XweoAJUkS+0OrB1Agjo9CJNegVUbEAJ1Ir9SOa5UjWTxyjgABb6q8CgqofC8J0PrUTxUoZHljYu
IDuNcY0onyBhJyEPKT7dDp1kcyZefAy6xJ7iJv1kdd7D58U21o2krhnKvhHMBLD+xoBVvB0XwJ8E
zXfM7SYbIp2JMw4lag+kwQmpsBkqC7ew4cLwju0yMOXu+xHZXxgfHo0N1gdU9zzKeuml2+PXji5J
d+Yky8nrnEnD2Cav99WAo4gCBdvRYMPAxwSqWrVZ4qB4avRLr5lh4gVxnxAw1y91Jigop3zf2V4g
I0KmyHrJLxp45KzMTiK45lswp0L5DnPI7+PHT/TcEv2TkjGBIrGT0Nf35yopqIJnupt01MAW6WiV
Kn5oAH4uEYO7snXTP3/dtJubOa/vQXTGRhugR/R3s2fafY0JVdsD4+XxQGTsjsjcBE2Y1vIJkj7j
gNcLVio+yioCCwqRFFsV7EdaFIPcNAHpCxarbaflK9lFVCm6n7X9KvyjWFAVx9Ljp1FL9ngIedPP
qp70kYIBLG73wpfWDyN2hht5PfMFJHDcCKtyHUPTO4eNe+6MD1ClLA22V8pNr+he3n1O+B9/oBbn
Cd0HOauRGnabLWA9hCF3qmVmDmfL/9BLbQ+u9HN7ZmdURBPK/F56XKGUFn6n0TXXJq7k/qnLMUXL
u0lwV1Woy+cGjtrupVarwGsG2COetKc1De3g35N+FBofB6ro9O7rfIL6lyZbA0XgZWU/wLH7YvC/
zdAQCwAf4heeGCyn5lO1XNsmXhvoYIM7E7sUNEcojwAKvD2c7rJ5GPJqUN0QSHIBml7nZnOrp/Q9
Bo3dKkkEENdjk8uf3FHXrsjNnisSh0+WMlcCb7cGSuhY7uE3bhIvn/vzvGYt1Iw9vASc4cAawDv6
FiyUlqsbJAGvwTIn2ogjv439GK6PKGU6s50l1eDfk+SnzJUnUqTuPBNdbc59uhWdMqgHsm21vSt+
zoj6VO/tzF1ITFL4MwfxGw5UWUgzleLu3XMbZIi1gBZp06DzTtZkYzKws/GSgFRsr18faEV+tuNW
Rspltz1M2GwsPqi45+GS/lAwO0MDIJ5EXI09bxF/oJZwmjtTJTdXLt/QFTDFptcZi1B67D0ISj19
ZbPB6r702dVdhromG58hn82vcc7MPwxz0LAt1C5ZKhlL1q+zjv5gbBvYu70Ny4mZNvCpe8MuSXwq
VpKnnydHB+32xPCHXr+huTtIMmBH/nrMkSJ5FFB4tdDWj36toKXM+XLQaZnFgjvAQRKl+vsVZ/Um
jDmy57qNVPQcxjARpp+SB/qJJJU6DJIg9XgulJ31ok8de1ZpqEn1VPZj9sxATIdMIE0tpkLRsPId
wVszCT8Bytrg7kSCPlC6J41KVvfdKRbKmfcl/j7gEcBM2aCRfsfwIE1W74IOIwM5SCL4EQRVM+Wo
N7ffBOP09azGRPgyvd+n+eF0Exs6hLbrzdWsJn2PrVSZOt7SZx7O9i3S2AvBNQZ1VHFWg8u9ltGN
T4Tb7j3pDmXTrFTs45mdGVJxCDTNCl0n4TWol4yE6GI2qJJ6CtlCYSV6nl9VdGCqO6gSREctwVCZ
CI8lsYa9Ev0tmvxwTU+jZPXragc+N4TvlstIqcVYcgJx85mhhxhkq4YrWPlq8vC1CMm48V4LGlZW
ZGE95V732Ke+4UZyOeA+kcsJt2ZPE7UNv6DSmKB8M6kbQdDecwTP8Zbi1qnwyrUcUMyjppOWgliN
iHq2GgFYzwgiAg2pNVuJuNWRR/0KWhlFUYa8NFwaFj0rIzQVVFIdkpYyM1/EzyLF0mzUHrPGgRyl
ykMjITczgkzMz1yHmd6n7/+2qvuX94d5Pzi/7euwdm/1ze3A6U963GULuwOFHsh7nx3q5jWlR7h4
qIxEEKGlGKNouAMtDNl2zhxTlp2NxgmrgTB7fubXKd5SNDd9owl27PoHgr9p9ykGpkJQcPIfZ5SY
VknvNOUJ666bE+4cfXLSFuk94oiJeijm3jTx2uwdvNkzLkOF+73Sza/CpLlgAcQRGKFjd+cBLBy9
S4cARehO8NRyNeGcXfZyLfu0TBOA9kK7LiRAVcwwjvdZtdsmdn45x6qUYd49n2RAIE+raBU9BF1X
IMojfjWJ9YochbdRQOXZ5jWap5KmxIaF7Hzs3hBph6jaLJbDFkq37LqnrTF+x+7ZxasBaERHnIM4
zTbpqTfEia/pEoeBdKM2R3NiZrgYHX+18eIwf+tuCWwH42v2fRGpeJeJIiUSML8Ie4/Nh4KGIV9f
VvDdjJ7b0bm+CRAro2MLmaCnM6kypBDySLe/bOL3Hef/CEnVBSzb5LockcgRnRZbjMu77AOXREu2
k4pIxiBYd39pXJhCukew0R8J8nFteis+gH1q643/Souuhlwj8nEr/YNUHMIwHwqfcaqM2+jeocDY
X9DTOmifb1yhlpQ3QH8FhK3FjsEaEeQbP4YxSb+lTa5jT4APgpVP3bSz9cUs5Ri/FUW/PiKchrg0
wnv+axw6EfMIQUw4lxdGfARobSMKdrb509QXmYDJr76uudmWC3puO+BX+pTmbTwxXoVJGv0EdJdL
5jTaH/vcAVdzOy1uxTR2RYTaTJ7vn8ibOKEwdX5aPjYW30LbL0itlnaSiOpYUHMjaayA4YfdiqKg
VV3U5Dh84EfUXVj8068qxnfKr1y6kVB4hu/emLb7L5GBUmFovXTifIviFMDSGsOC7QH3G4mS5ePE
ZOxaGwgmD9QXq3Zpg+DWeNwFgoh/s7Ng53MoDp07XtyXPkZRAntb3qG7AhS9ioh9AlDAIzkpbL4D
k+aAn/clU5ySiuOOcRklH1Lui+rV+4S8z+O7mUH8GwktwO7qW7vo4RpOYj9aFTgZ7TATfvSLgswK
7xFaiqMuLhP12Pc3cAwNM/oqZ4ontcSoL04lW637JimQotPQMq+ima/6vFlCZwIJZ7H20LDgNMBD
rRX/CgvivHLQob+KUwroRpgea67YotY3fdPLIUdoRo8E7VsQ/9m68TWwxfr4qYrxYHvCx7nb+2AU
iTnPs5DfeBLU9x2HeXB9T98RRbRiuFJxoBwCV9frMXaFIThch7J6MocUr+E44to1s5lRvgZDMTuh
ScOlSHn9fI+mNmuvpjv4p51cp2l+f/KC+egV+MzHG0O9lgTXeUkm71vuHQP90Gi+4IzGBA/vxLHl
7AO1N0NBnSskakm4augVHloZFddvSNfpC71G2BPMEMAb+U2h4X6vyjgBWMH+cq51GcryFO043NHZ
6fo93xbX/5hAvxqFahYFHarZiSJN6POkXmgFrJJxGtgNXgAjhlDn8A9n852PTkfzxMKrX7YltP7I
myK9XQ2Ku2YURY6jhuVs7xr2k16zXCs1Qq+6Q6qRWPWmethmkJZqDHWpaB8lF7Juz9altEVTyeOA
9ZSr4MhnakN/jctJ36rkoAhmBzZg31lLbFJvu2RKSfR7hekl8yJYm0+D/qGr6Kmj7HNXaJ5V769t
b6Ip6lvDWMPTTQvJerZiunWHtxBTlnkkc7WQDYdAoVdvdCKRCglpHl1Ok0f8qWcYao+/yhX9Z67b
Z2/V+2jqjS1lFZpc2o76l0l+XZk4AFy02PknnT3m1iqmu4EWIq8sW/LlvklNveIEIYhst95yE6Pm
71JY5TpMy8Lg/DdQ3GG7OlzBzwqaiszL1z0jeL9CRry50akQClV7We3msN1c15jZDcteREL3n32H
+t9KVm5Wl8NlMDY2cDPN0MYb3LoHOb6MwQTZBxFPhtoeB/qxERoDJ7IsdnNqM5xRuBMueWxcFyVp
bFWcG0E6I6ZsJJyHKCXQMtsm1yIPjkn6J2Lsi759ThOsLmhUhQKpQF/K+6hi+gR8JrZbJ92YEQpu
rCEK8aHPSxpUJbh0MdiyyE2/wUUdMio0LmKSvVH+TRzqcI6OPj1xVFd1uobi4Fpj6WoOOi6KV4LM
MwWrCA7j7B0Fm4HRSiW/3W8K2Bgck5Re8hi6x/PETvZAsq2hJUWWPwATgoPVyNHkd55fQI5gnre7
Cm9zbwL4rmKkyvWFhPhIzrborZP5O8GmpmsJxVI5avHHy0ZDuTn5xBGDiHVz98xplDn/ykxvPUxD
fLX5b5epWHYUcWqS0ozz7AEYJVI5CVJB4s3vFT5+JkYmsVhWihDyKz4zHP8yBwAGhVQ2HDjm5Zre
L3J/Caz9L2detq35/BpetnxbKrZmmzpKYaHNbxpml7TnjvPOHq7i5k7/GNPtoWEtQc1JcgWqVWTh
hrDh9m0QeBdyLk02fpzq3mDcdWerpJzlD1zOG+hnGQJ/6QharWx+SGkbP2WdZf4EeNcfxziu2KBQ
Uy6nkG1TvJ7y3VsiCZjOKe0GYFa3eq/oTl7YcgtKGka8yNjmI5Xt+u7YQCzEeFPXyQg93SRqFh0v
UTwwTUgEodkwR8LaN31K8OcgPEbnfarum8IhK/DmSkyT97/wWYW5lGMlFI5sm5OpxXicd/XseS3q
0awVHdaSFu6W8yl5/YJjqjJl+wXwvVLGS2oGkYENR5/FudJGt/I0JPhXzkycJZBibgXXBmlpxvqS
ASw8N+4HwkO1/+5OLTtyF/FQdtT7FljFEr9wx7gaP3VeL0fEqkGfeWBjwuFyo67vcLPHcWefrTc4
VdTfXFkZSfyt++cNembVyEUlHoliDQYdx2v+B0tw0Ty0zxfjSI0J/MOu7FodXBcGgLGrdGb3Vzkm
YYpjUBZpWJd5f6ks0GtY8IUWaGjCBxdKoHVgWoyBjb6LCPqdiD0OQCxuvpJqO2CG6ykvJo7fQX2X
NRuyGIVHxo5rWITnMvq33/vBgat7l9eDhFsQNGchTeu5Vy/z3DzZO8f+Ix+tyRpMsaAGCgPv1XM2
zYfE8msr4f9Pfq1t8YfwXVmW5bfTSHojhO5T+adhJrvwu0byaEPrg1A89hlEmUx48ktv6j9mJpGq
FlOq/jlAcVDB1mKbx+WTHPI101Ot2Oo3BFm3Yub9rz9dJMi9RRyxz/xQv/qQ5UguRBj4mS976BOI
XcRuHMFCs9x3+SneGBrkIgqReQL5vn31ffqZidC6hRiW5/G6LrgsvsrhufVVjdxCrrYJw7ZHlcuZ
MXuK6rQIHRzf9Kh40lJjqfiQdnKMDErFSg4V/XQfIolZjkRB74OwHSklVMw0C5TBjNbmR0aoMN15
ULgCskY7oH8ffGrqgDc2+OOU01LuD/Naz9f+hUby2BFZ1A+Z0K3tzyD+oeh97ali/6ptggtxWzs3
U6LPdaUUpGB9EBwdVZ/aqqde7urekfSpuXSmfLXWsaNqIOt8PPMFCiI+OV/DScv7ROfZqnPXAj6B
Bh1PmQhUkBMUzhKAm7gkwCrHCQRHGRn5pPp9HbxRsFJeybgFVc0mwcFsIpHGWxFIV9MNIDg79NyI
NZRR39GJMp28fyYHJucUsB9EHUUe9d7zHrgFnZgPtAV/nEHuHUC88xpdcUIZ5LNkZ+Gy/5rDYhV8
Zh0OwFmhYBpSoigXSMGGmyG9zfZMFEqCFybmIoocI96Po/IUaN6Xhmq52UyCK1B4RaHjwZugF2wv
v2Wvt9CH/3up1zBsmBNlYaNPA8fOsRkDGeWOmBZbofiXwgVnEk35dgWggVxx4tgqdwcNUBqai5hi
JVdQXh+w6b5/R1whC5IwtZSWJV2Ta6Hj24ZwqqqRi8ZecF5v2q18v8eHbQzwdiDii9V8CcIkKeqO
eFRUp2GVPp05hiQoWQyxKzysPjnJsMWcMKDtPs829pOh9ARfCIUrt5YDieBZPAuWBULpl4cMm8iz
+wE5czEeH8vJlqmGGyV3x/3fqI2rL3tmjzmrNTiXoU1trf9ywHa4NrU89I+OceIM7TRnCjKCYYBQ
Ab1vL+LMCoIfyL5yQ95OL4REQcSucbnSe0x6MUdsDX0SSRvWfvJKY4TRfXT+tCrVM61NJOSUmg8Z
gz0DlkQ7W4YCdY6xViwKVgR75czaB2v7GkdEPoUfGqj2mAT7OgAs4vs+590dH926bbacUS70xlPv
LEBf+6jdoaW8bS1XA1iYoPuBVZmFg1hp+hDHXP2mghP5R90nFaq5EG+3GY3xHs6oPluB83A8XpqE
cHivDSwi4K+jTLWMPtCKGnjpjc9kE3xrM1nVpzD0svltvAOyFp/rfOmJJGVeBTabhwc7erwAH8eo
q9Za1mWUDg1yeuT5z9Kvn1bsJhzb2DNtfxTI8wFrpG/WLwNsQkCf8WvH2Tc8ACpgLbIs9JypsBoM
C5D08hrBCSxuaNmrq8esR7Z4WAiU2NjWWtLvSa1KX7Jdx7uulrV0OLEYZkFznQKWYn26j3mdnPRo
3KPvsN6KB3f7Hl7zGlh0WScwlq7dwZr5OXgdQ/WAlxQyVKrVYsyjCXjN9Pb3yPzkjHfX17UyZXhH
tRsMxzjPhcBaoExfxG8yqOT6CYJSZ/bZJCckHfDKMiJHro8mh9YbT9YybC6YifGnlGBvlQA9bnw9
jz9WvWqyXad0pLTQvai+It1dMvgEC0uYuPL6T7PTuVYDkiSYUW7vcaur7U3jq5I0hSgQC1IPEbl6
K9/bhQ+BhR3OBGant/QH//bhejbklFVn7uO9Wjt2QY6+QoBDQro1wOP8qKmZgKOeQH3clCIqdLjc
2NoZCRVYh3tMgV8HJkCWPXokHClavSE++a2TMszL0NGcm4HbaXZQjbgRkaQcR/c5goYVSnD+N7n6
t9r8byHbeLU833alXs7x5ugaDy+w7X0/Rs8cRQe8j2d6Iz7XEwoAoq8YKSyqXNH0xv+qUWC0vAb/
63UrZ+M6L1ZnHysWWWvrtOc6t66JPpch1i5hQ04GvcpHU22tgyaia2Pt5wd0tuGVtlMpZ6hLDbB3
G1kWOZNXmmHzkHh414LqS38G3uVJOtpKiz90/5ri+w6N8M7b4rrISlGSi1yavT+VxRZAuxNWwfiO
ohZpCf5ze1UbXAgF2usJ32IMVaQlbim8AMglwzmUWJXVEOT5CpSu/gTq0+6t/GhmebJICtSbdINf
LUF+ub4VuSgsI7YUk+Z1pxtXxuaivEt4HwKPpNWXHU9Ou2Ki9hfCFZ1s576sJB3+5ERB76LSqAGw
xi5sHt6gtvy9IZbV9OaGFw3rk+kQIGb0uuv3H9YiAIX9nUp6QV9zUxTarj9K6U//nFK7ty8Qlo5t
Ifl3xijPECu+vmQlgHI7DFc3mvxaV35NokEpiCd8DkIz2lmpQF8SR27iYjrd9mBpyIoL6PQnLIa9
fmOGKdtro11Zp1Y9REbKAZk2bEzhmn+7gA+LHKMWWtRERQBfer66kq6K5zgfdSPP2MD39CFT7Wxg
gc6DXMBRRS8AwYgT8f+LYHzOmtOFWxOe5//in0W3rWPmN00CWdOv/oFsVbseNoEOBqoR8uVwIRPd
cBNRWhIffUITBCt/B/2fXLZq6rk4SFBlXyWD9il1UbXVE1ylHciDeXfA/39EYs9d/Bf2ehM89o50
k9wbNsUAre/v8MKlJilmssCRKcL+PsiKeolmwPA4K10VCW+dYv/54VlDFFoVdjectBmv13JhGTkR
Oazp8H4igu1njYrkcdXpseH1AbjB/I8AbVgz5YTlxM3Lj4DpJFFePHewlU8hUDOhgn66gcpoUGqj
dofLgNqUe2UWySaRalk+yspRGTgGb30tvtnM1ZifpW1uZNyTD1KlcKt2Royttg5A0NxYCnljg01l
cQaS9dSXCqVgXgHHBHXXg7lrJQpzlWzGCvsFRCwWzzX+T0mk+LHNKPNATthqO0nNzrHwmuuxzYQf
TvrqMSe6kTWsTpW7hBs+uNfdRmtoIiVN1mB+IJrkYRtD6xVCXHVz4boX8YvclSgA6v4Ef7PMRf2W
UMlpsnzdhap1yrBCKDpPgC904XZxg614BU/VPDE7rwsaigfD/FWtT/Ax83fr6nrT5Eq94KnpveIy
mX/D414ihDRL5Xf0OtWLlDZbIV9zvkzqtpw9Ky5BbWDIwQZRY+t56Lmpo93zra2D2R4x0IgP0B1m
0nU7WbFfY5gDiB4C9fkB03GgY1fDsAERMxxYskO3ElLKCP1L1zXi3WLH96C1VbLRdr+Jaczx0U/N
SnZGc057HNQB07TRc98x+lQcEgO2ajrih9FK1/a34rtZNCb42f7Arhj1G9ln8bCLRH3/AWaWrwfn
f/63sPbTIs33c2Rno55U28xIBk6wEuKaX5A/GZ5FFoznne8g870YRHga1IL0HDNfjRdxYsDF937M
juw2FDhBSuIWQJkcdZfrwknwjm2z0LbI3r98Gfh6Ynuxmh0mTKZjKY+cQLciu8Sd1XVytt2iWJ7J
WCEHafvsQv1/RYpa2Lfs41YaoSuwZISnzVsvyne2rq4DXIQk6JwLXqFOXH/7BzWversNBAP6HFtY
VmIhbfQedlyoiU6409z6au08AlpYArIzNQYSP1nA2l3ohc5cqsZ1XuNRADPccrgE+VEnjXoRcz6J
GbXqunqzTCg6zWAihU2qvb81xglzCY0UAMpaw5P2Ki2ES9QkUQkROYVecxGcRetbNDfxJyNvejs+
ZYsktElzB8qzQ67wU2Fv3cd3pPTV5rtB++xdHqvIS0oyN/PTaVRXwSgTIvzabw0iZeREInQ1qT8W
iTybmmWR6Vn1HdXQ68+3jozTtazlJKcCBrg4awWbi7ushOGyXlrbO9G7AoYbMMRcjO9hfWJaZKnq
i5pBPrHJsZEUr6zqxt8CPRvRSZ2HbAg+9MeTXvOioZQv+nSJEo8Czp2ydZW9fkpKu4+bkGh4p6d7
hzk/rZ/wtxx9EQYcpCkiZ/KsPDt/cgUqg/v/uePBQ3c6m1ejTGEZu1Mtv8z70OSCIkF5rVyWWaE8
uHPFoYH5eY4Wg9NYHeA4zN2IanJG9YKwULGm2xOJT7qtLGcxpbliVjBWrTgmHYvj051mmZGf+hiO
/swNh8vTkUtoBnPmnhIS3hP0loT0gBlKJ7K4Tx6neyvxiGz6Rn/p3y3S+Kzu7KJsrUCP3OyTtf8W
5g3HvieFPOD2O0Ze9NUsncI8TXW13floedC4iCHYDYpCLCWxvpvjgdAVvn+vkkEVXHIPtZZ9YGRH
XjnIpJaar9zNwTBZj8KIsqwP9XF1ahKmHAvkqf0o3EsO9Ef6jf9N4vyX3ZB3jnJfkJrlr6FnuFsZ
+0eoPyFykcG4bQ2Tq1bs1JMvsL+osCIXkBUmKMjp5WqsCbMhgqZ7RG2DtiOGN+lhQTnDy2ExT7Cu
DILp/sqgSXfVvypaAIzkFxC27EjGDQXRZk+5ujohuk/t4eq6kVOXZbG4d1u8JzWb8XKFeH6nqrOb
8XZB+kAa0eIqKcvMnOGqZzpp8M7s85cgOMuvQgb+uH115u2E40Ha9Cz+3IIFCabDXkTmU0PZw7Km
xKhUi3J3f54c/Balun9DQBOERtmAMWFQs984etVGeJhJFoLhAd2BXzp8GD31zMxDimdbryQXINMR
xjPd08FvAK140o4+8UaD66JdFY28v/dxhOPsDbhaJHdYPX2/cBZdwTHQUnpVMY5b7uqJPeUv22iQ
ZBcjX8j+Y/M1zHMJu+zseKfBDWhB5YP7IERjKP+Kj/U2nNd+a1rUhJFXszm0JfhrGrJqjIMhfkw7
OFwRqBD5vcY+0CPFgTUg/y+UwckMAoqun2SAz+ry9aq0olH9YQ+EKH258Jeke3dm0WunAcvCu5AY
mlCEBarbehChnYth4BGjpmMpXyse1Iy3xVe9T9AATnTxsjlnUX1XL31WfdIFGj/cd8BRQlxUfy2m
n3+BPKAagWcTWY+n0BDf0JjR4mRN+9sl2lTpzaEkqWelkG0ZDv2XfhRYCoLMg9C2t8Oj3hDwaLoi
0q33GnbPOz8v3bPirZPqHLqP8Ydg9o9Pj2S3QyCihy3r516SyFaCkXKwfq2D2CUiKddUhdRQUiZM
VMJ1r1vsybl1zjOZeEd6HqTkI9x2YMXvCZqQ1GCXzBGNFvFDxJHHGUKcMVVXGVdFjIrLVUJsYEjs
Ui9dDG51rw1SF308NXVDgfEV181U2sn3d0OVuTQ/NGZyM7uyUzSau9JE7bxfCwl2bbE41tBYBOAq
IL+92H+ZlMVa1UPIEpCrVJdAGcRKhsE85XcbtA+iMSghDENzSmXPz1OoA27H64D0L4jnW96XNapM
Yp4x3a7cjr9c3D2SVlaBIy56uzBJDxI7jyIBSwjwPUqa8KWYVGvqwPuaCknfg06RHynUCacm8nW0
SEzeG8x9ROKqGhn4C9TteM8jfl3LTopd6m3nk5SiJG7l5s0jq/Rhmy0djvweXLO/Oy5SRgg0B59N
CVk2QHXj04SuLVZVI6kMKZKm4Pv/WrnciAIsKPFhVymvb0fNqBRos3Zpi8OAGGgOUNN2lCZMVAZ9
cHzzyhwJMQ+kMJ5XauWdAuAeobLPu2YT1ConJjW+NPAySZ6T3Nw4qv8+ubEFSqhCL2bOy2Tb1/7k
RWfvIX5VFeil/ohdRL4zaF+4t9Uvm491poHyi4cfi2QZX6qUcrMRVsHbBJCZrXdCmuNJFO9Aolqv
ZKaJdoXPojcFDhwhsevVADooBrQqQhXSZx9Aoj3+BYB+7eQnJSB8kglRSOK4qko9fdY25cxEuuES
DFSbmN4cSKFd7h23E/u+KJaDuBwRLjm12EOqOXpXBu+gylhMKgMJGd1bY4brvJ0ESyLyai4FQQAf
qWEac1lcAkCUq9Z+vRVFVtzrFf85d0DvD7TkKsDjv9hFYZ3m32itHGg2njwNK9uFvJRGPFNqrBsV
HDisNcPmgFxANqXc3Uuso3acXgTpJqGdbmHMgFl06qc3ONmOvgPRTh6CgiCnG31INhvGDkBvqQT1
e1m3ZutxoCFWI/vsB/b6dOLjvOtmWTM6dVggWlvbKUiHPTzOu00RyYVpmauqZq2QeIpMqoWeVnPV
KkTAct3dlxPNWBx9W19M467YYyPmoZbzQ6/0Llq+Hb2dDlTpkOmUxNWI2oZwziLF+hrpCZS+U9DE
eN5VifO3XUUX5m+9UAZvihWNw2sRkFA4WyurA14lbjTmY+mIaUFyOL9zfCzx0/B14GCO9L4/rAB2
U1WaW4jnQ5L2Bj3G/l/0th9v7oRA6rKTdwj0YUJDwVMWf82+82Y9lgj/r/1j9S1LY7cAGjQ+BdAd
gk37kCfEnfLGBphFClk/6+XjIJVjdgpd7k6BNmsok480k6O1HewNZoDEj5W6bR1AAg5gCHgR4nkg
KLkEN6nTlZ2vUPXNiSsZWUtgv+6ONWtdOPx36lWa9kmaA6Hhr/uuYShgeipEvT26eWQR87VVyC5J
+AB13lMb/3oa8mblW0Em4NBex0H2nEMTYLWBdmMK2/JYPW+8zTbzS/IWgq+2mI5CWcIOeI8+pN9Z
9sTJz7fmgWPjKe+uYaiX4uzrC01ytNAZnMJipcwZMp30Xzc75ZLp0MZBcufxJdENClEFTDH+kJcy
rdBKJFF2goWOttCZgcm8VMUXFZQcGh/IlfPp0hrZCJydsTcNoY9U/vVbEg/LyWYWw17hTUspowBF
H/iHoUmyw6TxhrZNJ7Diazb9eFfNJdWHgiCGcyBZrstlOJglxo+ASUVypZCVqf8pUmSHpvgMekmp
+iEiBXwVV974m/A4wz1ehjuJW7xO37//ylFOgx5aUhv64Vtp/aFyXCVxbTt4ZIiCnHQ+HdQZzPEh
6GtgeFRUs5vGcGgmplhsU9rbY/NCXW7gEAGm8WkJ+5JgVQatEeTDdxHJjFt/Ud4b8Fej+iLAv21I
k78j7MOOPNT+1+Q08Ff+b+Q9NhvFEy7VyhyMiIQAvgtVpppTzqRjJJKxwKwv9uKaN4V939nI/hgP
1wpPGXT6fTl2Is08NGUUearVj7LYzAJNClgr1BfR9gKNs8dh3AWi7FfwLgYmLnHCsiXefKH015ru
39gixLzy7/ybrCGQpc0Wn7Dd3/i9zfE1Fx69KoV5X9mPX+vxJ6rEcwBo6CBWWi2YMG3/Lx+gXl/Z
2QFGLksVLl6v9U37Ju9dPoRtsg6WYhKyit1XupUCmeLRixkb4frXlfpyafZrA814mXpL1xjoQruG
EGnB7xTgA2XVeifWzNX0qg51ZEqQyrscw750PhwrRImK1JjzV0eXWefVQjsDF2LPRMtBO0hUHVpP
L7lROO94ranl+phi8+20NrW1UkdGf5tC/O2B39ewmaCkCIuAC5dPslPGYJCbxARfjRUBFQQRV+2J
XIkKN79fR93bwbaA038RcTLJa7pT3QoFqD7zVKTCXWROP40CbLleWVY2o3l9yZwqxDy2IunSV5U5
xT/QVt5WRkJgjWkv3PeuZzSQ/KcRr8xdcZve6YF/+JIuTgTfjpW7UIWvkr7eHT4Mn9Zpq4Lo2qIm
lCCFAozYWvavUZ8p/VBM/gkWWHBHt/ukhrRoIegdtQYQxY+j/RZumze4zujgjTsmcf0HV1Kx1M0f
+kk92oYNm0WrEkup4O+f5u7rnCCoROTICqvUHqg8nSwmFQ6iw0xcPK4ART46KMlB78mHw34qAJTk
LNbDPQgKXYaMwr/aCmix9Oj3iAOXskKbPSCRaSOM8StQsOtN61mlH+KokG6jAdiIRlBOyh99oHHT
DgtU1Jl4nyVxb9RcHheE5R+zne0+MO9YaGLWg29gzxaPljQc5Ep9B3hMeVSQaHoAhXB/ivBqeOnc
/W5EOqIb7JpXzZbqoq402rBC9JOgxYm2toe54cCg3+ZOkt4tVYQV4YF/+AsrVSGVlFJTuW0OdlcG
RwNYPYXEHOhJMw0wMUTL5q7JXfteaJUmL+Dh7zFwyGZzO3TQFxSuRcNtKMfevt720oaAzFgpAeZZ
O9QtXoLcRPo8UzMmRyOWQYbMzC532psvat7S0b4nUgSHjWQDdzG8RNGlpt8/WPIaMgHQAlPniVmt
+6wldfP3bQvh4wfvYePHGSdbHGRQGVRff9D57qTlt7aBv+EBFAk+xKNtZGuDCIFUG5K8EC027i0W
9z6k2sxOeMXDXsK/lAdAkvpgxRmCh2CfEUvyCmWIegN7YFPIZLaS58dX8a4j7F4lrrFBcYQt3Uen
iKnMOAxMWRcR3iWlEb6rgbkMIs/s+09BuQKFYPxXPurrGKMhwKhvOfrJBAjSNRI0V5o2QbUr/Q6I
+mJPx7rcZzp+bUCu3xy2oGaHUWP/HSIwDtIX04pQSaQrxHYspSOWOmKhwWXzTVW9u/5NChlI3Gq0
JB+JL9vB1C39JbipFTnT1pPb4BG6astSAUAVyaMf3C1QqYe2NcWODGSamK/V3jumlbDy1cs7WKaV
IueYhRJ72x7g/Id52Ybdjbn1STj6Ghr9q5IqV30DoJadqtLxiSsDdS9N5q5222XZwslimc1iRkbT
xgd6TFtxb2FvxBPWDARJ5ius1xR9Mx8vgiS97/wH84yOk0J7qF0fS/0trI9GpNsLfpIKVZHCg6AK
nBmQP+hZ2dMNjPXtNqykDeMW2ut5nNbfJF8mlFt7lKBmkuGrM7qhUjZd1O7GE1jkdgHpqEMJRFD6
MQcGe4xXbIrqjk1l4aOsqJVBkH3OdcVGkAYrCjjKJhFT90QW9Ob4W668Y3vWK7LNaVBsYJJwSF2G
wR+Lx/neVZAVOLQhYmlqfYii3b+RTppP5GgV2Xa6732COXekKQfs+oSqLZ8rlSAfUJw/tx/Z1rM4
Uu3CrdLthE2qSAxpomsf2iDs5QTbA4HIK/hrM0EVJh3eIhCBM4+Y0jkJl5OD9pn/NBL3lwrLBGO0
Z0jIOCZ885ukrmM3++KdSZ6nq8/NwCHqBStf202IRZdfYTs5u/r4yRN2fJWqMowdIeMX7evJqim8
u3fnGpMf7bsK+MONnhIFA/sfmzOdrsUc+nfkMzh3N+gAAsl9lvxoHosM6hlTRySXhU2YyEqn7X6Y
85hG9adsaw+KwpOTeSTDnKu6zIRW7T2cOlkY7SxghP5tGrTZ5cKPGhdjBC7JppUpOwXuhT8E6Auk
6RnsrPQYOX1gbW5V7KCtw71r0ZicyXzolQ/imlekj3X0owiOoIfeuR3C/4BfTqB3AVrwk5HUvfRe
3CgGzz+bfplCwL4OUKuek+HYht1acZr9Ol4eh982yFQ7ybDG5fx9HavvTktSMPNeGf6hNQWpGt0A
ptPGHv9CIb8wP9/I0U6dn8NLgoAYoXgqTnBquoEtmF5CoRkMR4hQs1Pz0OsrWYZaGVyC78x6FQOo
lDWByAjaSAgTA2h89pzs3pOxjicJvj9r11jac7juRmixNmmTW1NcseDavxsWama4QGrSk3Yp5B1B
5Otr8mralQQyGcwQE3+J+HYlIBdEihex6d+HK7JBnEuBeP1derRD8BuuZf3oY9/SkK+N/Pc0aVhD
mYd7GqMiN3g4Y/82tMLif0kEPmagdCIMKTVhPTxje1I7c3s5pWXswamsFAtEKmp3QQVC5rnr6Vxu
BokNKUP2QpquGdHdCVznsnldZKfWucgZc1na0shrLuloi3oqjw+/yslUJA5x0kK9TOpDsnMZA9Ar
j7BtMDngVO/VZH+6FRqnWXXoS4JKmNpepEz8M66SnDcfn8fO2AoMZYeygP2S3xrEPZcZKhjC+/Xk
/XHzwELe/kRkk6VO74mBTmSBOIK9dms/vePW6xSkuKd3Szl6tUI4xP819wFRTLiaGXh87Yspnd13
BE3bzv7TSjOJf5daNUNSQvRp9X8QD1ERhK/e7i3qjG4pscReyjUmzIgxNOQS4eh364cgq9PXP4nS
/pR8KInDRD5w3F1BfuPiR1FWWC0KwpSo5motuyazwSAbWCafBycgKrhKhO+P8GuINpC1xmHhIbrB
Efbtk4cSlFspRdxNkt8rLEiXSKFrg7hG70sgx1Bkzvs9LAH1ivTLyL/5uX1YJgFs4igqiSrVXUyr
YC3Ihtyl6xb/hjCsKrMCStbX5lhfG/xZunMGKj1Ra7na9yT0//9S0nFc9kZ/1GmHVptPFyp0lkjk
u/GgI7Ywb9bWOywObEaviNqRDdSpTPuPJlDzQAeMrCrJ/SHF5jD2qXi6ectrdhFzjrEapGpglFHU
4zcblCd9UrtCTLC3FoIYsppsMJvNbLiQJ3vewirPifnb4js6k2eqosCNP9EhRjCZdoy/tYwe0gld
7st0Fl3nhxbEbLuP33VamZpRQMar3Nk9PbPTOvWPTYehGmx760aZD+jHPIw+BRPVK+B46roff8LW
vXD0oKMHMIl2xlNLQwcQXkDfkIdYwVgm2SEXWAkJvpIu4+Y3sPn2/hHJdwe0RTK1G569ehXKmL+5
Z9H0keaC9gN14oT4xdGJn2URlRI659ud1LWVtwJEeGwfI44i+H4WGK+XJadgw+ztY+D0C6o/te1j
iYi0j7CICXX+LCYAWIh5bkztwSUlhKdnwXn18ElYcTbZN2UY67ng81+9S+6avpakT/J6SzvJr/C4
UEklKVCSb+3ZIRs4xWvxYHvzalTNLJbQTe2+8ruVU9j7G/k0JqNKbqYO81Do4VtBltbtLtz0Ow3A
zNNiXZQz0bYAKdmvzDXUMDbMWX0FTeRgAs+GX+3R4NJa2EzPDl3oHXg3btlHVeJTfhCmVXiI/cAR
fR2G/8q5vW2033dMDA3WER2mFFyrejpVPVq+Bwyuel0iQYeFePj7LFdiArNS4NwUGvQhlFPX3Uo6
lmM6rAj8WIWHg12n8LLYxj+v9bPAQszeoVRAxEKtjJOdMi/z3yzWRqD06ZgqIybaLIONLNzHgRWF
nWD5PWx4UKhSzUD2/3aetL+yGhDcIuqVjbZ4V0rD0XUAFaLGIy9CYz0h1/npdSx3XBQ97sGSG9lE
KSnnv08bjKSGjvUwnNiIQ3wLdLrM1kcCA0iusLnH6ClP1/2RhvtNkoJGsfkfHAsrWhB/gzFYV/X0
uZAwpw9FZmKwgGcwPo8fJjogxfNwAi9bss9/ikSI+HoJyqxkS14Hg/E9PKOgjD9yafIDZuILT/Ut
lRU207O1HLB0y64g9I/d63Tw2ARK/dx8fI+Kr/3CqzFUb9ocMTEKLdZuRbV+B1Gp6tSiZ0QYddO0
uvJsxbGTS9XKXFrFCtkKJmG/W8YqQ+ZgGq5Ry4MzsLkSI0DUFUGwxgy/Bsn3K/8RmaeF4ryO+hOj
o4FTbIryt15FQnAI+n4NiiWt3q3dtaPqH2/hBGpNhNK76fb4Mm2p+Ws6GBRobJOjqxDyphEW50Q/
T7xEDctPjRCogfegyqQaVVrXxdoVmtRLglZV0/iiKoSWa8Ihy0IMl5aQM64yDecZeNzCWLpcOgMp
jCRlXklgZuUlLxWZGo6PiOxhA564CsGV+CY/A2lDrwYvKudkzstQixAu8WGSGO763JSn5uQJFKUU
BX5Jd6Cri2nMbi/pGGYj+5j5/26aWxboptm/CwftQCb6MycRU6ddDC2ehD2nr8x7Zucl+PbTIVxv
CazHmOgb4heeNKMk4G6kzPie6ZCiGGou4S3mi+HsiTr9md9PoQWHxSu75AOZvMtWYI8I+TPS/NIa
sqrVaDN7lg5xKGzCOb5EltxwCLuWbNFA5r/TKYPa4TspQxpAYm8fpF4Gl5Mb5mqpZf44w/ADX+jB
hgQLLZpkrTD9YEck9XZegFPpuALfl1OGIeg1ecwzR2cbPX8d+AglKVtLrmOm97IRIUL8jyjhTciD
L73I/BI3JJD7d2MInk4Phjb9PMkdohwCfzs6Vh12KhV6spRYhzVDgtGLZZpdDg80ehwoBcA167c3
+eEend0XuPF8mSXj0r05OeLFrPxsiVevqVO3XLka1OoSVy3+K6k8fWle2aLiyou3CxHQ0BU0eHWq
wvf5lZMf1ok+eE+Jy5y+ujc8+5nCY5UYQHrJPgiltsVeEH6usvVqI8knsbjUITkkmP2lms1mrL3J
avlpJP7UzZTnYzlcLBhnqHXRIXWlV36MRBgh0a0sCcEClEjZWCHzCw2H7O8CUnMdSbweAgC8mq9x
ezyVRhRDffG4l76u6gdvY2iffW+CEwtwVPjDSU18CJR/upZ52EhmEraDZMxeQJcJxUT9CLQzN1ms
/ev+Wh//QBm8o/uqeljFlkrjRu8P+9V69Z3MD+VLtl07ZyuqkUEQdU4twMz9CW40KbeGhM5Two7P
5Kd3JsRchL4Go+te5g2AJ1Fjq+gS8AeIcfb0xNZAeoZ8OnG/bHIPTLQqKbHJds+liYE7iJQiayhV
MzW67c+8MgP0kEryB5TlfMfih3tTikTSGDjSkNFAI88uZ3Z1HilYf87sAC5lt4AIblRpsuUYUgY8
QZscz4qVmDxWrCTj4bgU9RIK3xmlcJ3c3j9ha0d46V3GvY5nRPA4QEctFAulX+WOWBL5O8HWiDxw
eECF2rjtL6MSb1d1PeAhCb/ybo7Y2qMohnDKADyM2oaXHikRyD2aeKiQetnw60Lq45UOUzVa5NbD
THpFA+d9Wn8SDTSNlfxp1/MOfQXmAryKOE33bAWZdvRSsUUflfHz8vd3RxJlD6Jzrum5E+sRigQZ
+XROfKI1wzuuQNaXX3h9VPWkseDrfOVGuYRjt5pORRDuGXC5IOJ3OMWPX2Kml653fDARexixZ0Aq
mMH/yzi7zTqBsLyXtn5GZYsb6KE0KyvXLWQn5SiMKpFXr4yUUYz+5Y4Clyuyco+MEznijpkvwkec
lEi/GZpYjXcYELQyODwAKUpycXw6C5p6Zg71D6vgMnFyiUhrX2fLqPLc+OR0Aj+cJ/d6k8MWdEc2
PhmnPFnxMmVwRMUQVKolH7FdnOBRR+sTLR39CE2K3FI9tlDhfnUkWo/ZJ2+w0GTYMdtak/9KYzDA
PwoXvCdvNK9SuE+vxBWD5oBomKA1QRSohNL1BX0MRyVL+3RKolfG4HylKO4J1qHbiMKGlQhyNE5H
q+mjZo0FtGeC1ev+n51t+AOwX9BlCQJlYtoZ8Sl9LF3OUGIBqcdnMOWJxrJSl21dpN6wu4vuHVUh
KnfauQDvBKI8s+5guwanvwRpzAnGlBfZO3WYJNbzeyPuoy9Mrz5UvK5Kkgap/8UFoWGevMFP9aTS
yzDB78427DC1p7Dc1aptz+WTvC7zysKaH1mwYaO6lh0OXeBo6PI+pezuopLajmB93Te7Zpic7cF5
7O+MYwdBAOM98j2xeZbyuDgWnSo8roaoEANdfPUEWm9rJDxzVEyHefqDLcvwBokPy7gn9uyjnY0B
d26Kz+wEhUrZA1ZzaYRWZWtD9N3W0Azz+SBCvgG1bcXRivRmx1QNRWrEoXp4DnsQd2ORovJT7OhG
xr+GnX2+YGpI8OH3v0/cIxnv8QbJQDLxn0N2TLvCCjuyniAyqJ6EAiXi0/wIDaLuPm1MKptlIC9S
qxIJ7lDFu5H53b7xVfsSc2EKoPk8HvwpEptcCFq6aX0GHaz83S9JJ4J9MxpC7dzxE8uHgCwN+0Qe
m02FpYXcWIRSUtR5e1xOO/Xy+GXt6BrEGhmmSb2lNpS7/2EpwXYxw4dsVCwUOrDLOhuIndM2hhqF
8vh+ZvT5dT17UmwTeGbEKdtqWgsT8LsJvKw9UC4yFPY0ad08syiqZ2Rv/n50Ho8AeVbaV+uJsTui
uyoXAIm15dcNXsQcIGGJYawtAwNOAULKxk0WRCvmr7IYXSMdhsAdFtu15yeUbUzmoGRZ9H592yfD
ZM3oNeUf/VctrexQeLFgzCnIXEPcJG57JHqLe+VODPyDfos6rpKDa1I5prIF/tPTN9/H/0lNg+07
DWC/BFqRlRBWXgB+qmdxQoWgHwzqzn8sW/EbZk+O92Z1RoQffWKz2eUN9+eyQc8Qh3/2W9ndRXC9
plaTrGi1nSwhh+/lRB/Ic4eKu8q8XWsFBUWcMt7Af8OoMLig2nH3TIRuuJ3/QmbDaYCBf18gAkUT
Hrrjgg6k8UlDHiAV2nzQ859aXCEKgbJ37eYDGuOXtdp1B9PSpC+oucDItRJdRpHpNe8Sf7FygeRb
FZBRBO+nmkg4Wc5LhKpA5wGpQbqlaVUM1Kho6Ln1vgaHSQ90gKALw0yE0O6dmV1ENW6WfM6/pYaD
jcxqFuAN6FxXTXd1oKgXsJh3/ku40HEdsuyIpI7sI4z9mvvGkM+hPMZjwY2AbooxWLpzpI6As/zn
rGfZ0CTCIunLQtI4ZGhi4KVM3zPV5Yxe2qgcSVxVPjc6t//E4AtMVazEPB+W/Su3WRINqhu3jC10
KwWMnVR1GuD45rUUGprPUmRpsX1VUkwoHvIHh1CGnGtVc/L+FE9kabbClFiGHsZHSlIT2CXk+hUS
nlR+uvCBp8cfO7wm9WACwf3OcrTTCP1eNEvtfip+LFX8nzKPR420N/p5oLnCz7CEBC3svifXZTRG
g6HG2GIw5389mIv8/3QM9TA8SzfBrYBcC8UoIU4wZNpNvRxQg3qLgpekRlObQz/I2ErptVsAYwF/
BqqEgWtDDXGFY7xmJidYyyDKOfFDvpj75J9Dt+GMkeOILGP8V8ZsXqD/U2JsJzsmAkN6mPvbuGVU
DeLma2tu6zvHJryIUf3U8YZ9L3wODjW6hYCSMLAHIN0txmy46G8bFGLLKyMZw2ub1pe6i96EvIPz
nsUy+0u2iIH8kS62lHxqSWQu6EJEDvxBV654Mmk+VK5wvs/+8/RYnV3eGEqPgpyB/9UfXBhYTF5X
53+sFY4CgrFBfkNn2ZC7mTcxUhFWVSCtwcP4z0HtqWqD4Ux9YJUWIK1CotiBLrcOAqHzeFSapm1+
DzCOdkRCXsR4chmiXfqeExvjZTXHkXrcftE/fUlrNLuQO/DzSNNRSinnAOv8UBnay3lYWXax6kI1
LoE4yrcHYJBs75V0c25ki24FzhRjZKPS4KImuiR5DyRfihsWtdUlgwKDxsvfzlZ4IrFn7riH+ES/
bE8/HZRbqjaUSD/gtrB+LDR3YzllgZSEhaMCc5nWPVUSNUCpImcXx223PdajjtAXSK7pNFV++5H2
k28Vy6tI0OKCDvAJVM9eKMApbLi9fTvaiLI/fXDkY4+krwt7u5VeDJpUarzF773fOX9sNR93fVu7
EWAXRnsWRUyE5JUXjqTJTmmIx4SHxlQ87s2+b3AMLn/wT3XljOiLr8BzOz7XgIKpIUb6Epq32hwr
h/fdiSm+4OQ1lvoXeXifMzzuFWcJWjjG99hZTWNCRAp/j4G+26JVhgQVdDDidBHfKLP5MBoVx28U
5+grXXO+PBZRTrtv7VArR5qYCnuz4Dc9/FB8U9iFCgEKW6binuIQraLbsGbvylkocPzHiN3FWQBH
Yi/1Q+vp6y2UXx0SPbCy1EP1kP8PA66+K4TX2dq8uWtH8F+W1xV50bJr9uUB6uBzWvA6TKdZBmnW
A+MNjD9+8hfqdslKcy9ZH+bq5697PgszW+ASxQdPGXY+xUiGs3zVXLpf27MrKcx5NMVsd0H6ifTw
kgVhe6j4nj8tmkRers3v2X7e/QAeHA7rjMZV4gC4xUsjkpuVJ/DFk+xbgRW/p/L3MQ0pUvZ8wvZF
QXenyxPaswoHFZ13sTIwChkt+7mZENRDXKT1QHyCQQzKYPjfcfqtf/vJGXCRLAUytnSVdD6OmDqn
488jAESlOFXP6/FjseD3GHVlM2ltX0ESLoPGNDquWlyGvfh7EXSq1QCldPvw9Xr+1JHKp+SLSpHV
YsIAYy9VoKW+8ETdwZ98G8+BK+TtdUd0sRAAU5B+6V6zhRt8+LMVeMRR2QsD9XInOGwg2T50ss7c
oT84wK1vK/3GSBd+ruX3AmVNmApjqsIZsAn8nv5//XFsVJsiGme4okF2JO/CVJrpFOF7Q5kkXYXm
ywJNG/8SNZl10yYb7vaCd2b4q5uCVv+hDANUQLQSytfwL6MWair4xEIGHRwWCmXVBA1DhAua/nI6
Jc1R6F9VQognlqvGuoW7XEpynW1ksK0dP9+x7TqrHaoZfQbv8oXIktd8iLAHG/W0+4lt5uqIQmLk
IJJuoC19iwmJR48oEfVdFL+h/navtnLFgMlHniOe08Ax1anRpHKZcZcB2545iO9MZscXwRL4sa+7
3YB5IbXho+LpfKLUrhsLfaxh2147IfZ+ZiCGZnYdRhl4ymtcKflXLo+3bhwZHjmhDCIposDxLjR5
ZsEcfpEjF+QXxdniZZbmP4MTHsAGjgFFK1sX7K/PfZ5RgljmWChPUd1MAa4aXK3pB1TA8dzuNXQS
/ltut6HLmnDNSBj9ebtiP20bc9Ycd6bvq+6U9Lh+4SQZleWTQWFYSudtzbt+NW4q6VwjVoZ8vViN
T4CwHzkSS+eIpNiKy1ZHaygCX4bep6uHIMEb7YSBdr/kPEZjKorRmz5FU/VzpEB7vHVwuRurqtLU
s7TiyVX+3fPpKOPo3hoq16EqvdwXQ4sJftsqtKFg8kO9Zw71ftaXgKtYtYah4N5cND1EepxzZ4dn
XSf0WhnFArCRqp6uRJy8arW659H/W0Adtd3pD/3YHF6tyV9R6KweNlbpmsGWKFEO+vyexHhnx1UB
oDOn5uzr9V1EoCZqZKn7uDrEM37H6SYvrzlo07Np3SL1nUvGYARIlZXJCCvbjtiO1VLTrTCi3fk0
lknIUkfd0MxESc2jHqUmuE87kTdpI0TJ4Nv3KKz3tA4jrrfg7GjlnQjfJNH90jCgR5u8gdbWIMi1
kXLQhhnkdfKk56i8tw4mzX1/16IXtfbylKgKjpFltX01Viv+6ekU6KyQYaxSdINkcm4T11c823rP
3PojdAFIoS0unSjzFs2OlfNnQ1JUy5297/iTzHjENcyOrwehQ6qbSMJNeYqATyWsgFMLtiywFtJ7
IeNsilNmp+LptiaU3eUWtlEuS7QtsLMMG9UzyvyT8NLXkn4s2+7CP/qdHHabB0XCrgSOfvdUSbJc
iEG3Xs1QogUE3GKFi/7wJqBcO0QJG0Mwwie1CdD1cdpc5C1xJ6zenRKxJ7KVUQDmqwBYW38Db+Qm
ARvY3pJGlxtJuIQbl9zFI9/NBREoeepFtnmdcj9MxZwz7Se8up0CHWvzsbzdBc/z/iKPRQWeS6ta
R7OKeiX84LqY+7BNxHqX2peEJXbgTmE5j9GPrIHkPniBM+kGrNxrK1uYS2ea+Jvz5gUl0mXtCa36
Q2/zCpXqvpgRkizcwIBh50x37jn+kjB2qO2eeO+4L3u1ID2qc1LTQWV+TKtnxa8L9gQOlqfA2Y93
U8h9PPaQKCCFweHM6ZIaZ5U+0hvrn9AK8Q7J8Xf+OVuJmNt99w97ytYmBYRtU82JOs8pUdFt+iXw
NGD6LCxum0zB0ii+9kByVYpaNR2hMr7lvexJ3tOWmWsumMrZyKioxuuUCSpLmFyO0dWbnTLw7g57
/Mk9kq2rUZbajyeMJxRHVlZThnb/gL/q6Vr2mo3qcwtQJYXqwu3eX8r9FgHUKpYmd6/fuO0g5HhH
EUFX232qzUDUpaZdXVljgSYTwW7ndlTLNiV46cFUVOzGCqcDCqbBDIbSv/IvNVT6LuPdmqe7TiSN
2BmXG6TDDhGAl/a3JKnIbSNXa6vK4a485YfCLV+VVorF6Oe/i7QeXuEZcr+7omNbfoGwT28fA5F+
w9TwnRPJPU+o5ccwQNRDuM6EJyBd8LmAx8+WZPn5EoOVD74wBVHePjruZ2cairtz11WUOfpFKQ+W
CHXFzmCdrMB61GFcPagrW9o9vDW8RW1BWZSas4q9fysQLp5YIc6MvRpvhD/D44zGw7ZCTJjt7S5d
1SS/wvA8P4CFRycHs9RJcfdPgVfQyGjXneDcPDch20lA9oAJy7uhulbkp+o/QCoK+6p/BPVSzcAF
e9uQbcuoF6BmMC1wk0Oix5hZdqNWlZ6uLkxIxzZjtAGAGSW4aEfRV8cZlrtJKuGAEh01niYSELKV
4XKpmmwd8WmuRThC58UW3qkiUF+aHcO84g4cP8W4Vdmkktnu6XZ1vxysMjtq5YGo0JnW0KBW8VOl
BhdjgeZe6U3/1T8/GagSHYvSscfyaEqcbjVrPyvPvsPJFkzb3yH+roGyrA6+uVNw81W6h2XT/QCp
LGZIa6VH+DpOYzGDhYccTaerASDkWQIMItyRuEx+8Z82eEastzdiJlZgWJQcRcdAGqEcj2eNoq4e
qPp3fwF1gcoQtQGFPCMQ91qld2fLN5dRxgcOfWuybikYilj2a0E+WWQJzyHu65/yqUGpAgn4iX1c
sxrfF9WRwHFNje8yRHBiY/PUkTmkLePjlYDYMSAI4VDdyfy2QIq8gzZDnVo/ESMCDbLeTxn+x7CX
lVu1IGgF7lPTLCvWL1eV4cPjz+Qyo6tcmClNmxuku/7J0qUiYMB5WwB13g5fPT4xsOvZIciVGKhg
78Q9Krk36oNe8o5A+KT8YqcxR914cLvWXfVhtCiPaEdqPMelyTT932xTW267N83SlsC6fZaDQkxB
kWHP0zLNiEzw+dkCaWKhwskoSCesyZT1j9VnkVVqQFOb35w2VmE0QbsQzBinNbAkwds3RU6A7j0N
joK61VmOoeSofhIjvoDS/+NulOq8yjkRKhvppQUC6fhNFukAC23GoucxDXR6HoNigVFObmQ0ME6M
Szms5KkEc/4ZetmSvD75eX9lOusU01h3rpYzjD0FE1n6LvzigDB9aXJ4pbvqDNV1r3RKFi93GTa+
bqRTN0v6G0zO1hoYKzDxi1qZgb434Jc3Q08Ib18vnajAu37c7mFSeGMpG84bYH7N98b5ySF2dddB
/H52Vfus3Syv9pGYGPVSGWqzysRUvgKEso0TfVbr5wuRcJyM53PLwANKTiytvm4f9Sy1D0WGU/Zn
15VZkAgqGJL57S0GodJ+//lE+A370TPoltkHeVMKwQEQiv6pQKG9BcaQhRW3ULps0UtDv42h0ZH6
6V4QzRhwLIZjvOBlQLgMAwwYoFe2Rt9kzi8hBzt82k9WYpe4cL76Wje0s+IIzv69L3/bR3z/ux9a
31GWHi+17Tjphhc1jRS8jJrHjTm9wi0vjYXQLUtie4dSHxCH9+skvRcsbIivbmElHAjRcvAiAwZ/
B8luuLiDvVFoQshXNjVfrIMGLe1atCJWj0gXlICHurRdx894zAtRHgoCOyT8fwYIEMci11E4vuqp
P9Yh0LUYSnQ5QAXdwKOmWR0CVi9Weloq5COfwtmEvQ4oVoBFCSuDhe5Aq2PaAUFLwArxcf76z5kf
9H4E3xITZrm8cUSEGC1VaqaCaxhXjExUj+TWlGp3Jk7n9yo4Rim8xVF4cSBLwbkhq9QVdA9yWKEm
AdjkjRDqYMCSvxgcv7L7Gf6W1p0vsAmSCWk0FVpsZp3xad6+UTja3lLpXXjSiM753zHtEpMyxlnK
1rX4l8aPlP1y33mIDE0uAW9hF/iz5fsTLzBkWP1rYBzE4nV4O9iDGvUUgAnlkiIfE1yYgRjiIFnU
KkttL42YO1nSNJZsRSj7gKxM3RS44uAp9mgN4kPzwur/yW/QTHNeYc/Cy+o1b7d02fhNfgEvITa8
VLYW8Pe74LUvhAWUsqdv/NJQNpKBP6aEY3trPZlwRSlPrgFkzajEqplmEvlCa1VkYitRaYub9jlJ
SJDl30B4rh7KV7lNrdysPyewRTH3WVVhObva5QK2upjn9V+ShsohCoOhQTen3mcm4aJX8ugbzkxL
5dr3b/MOvlTn/oTAsS69bOHgRtrXrmeyGuoYH+97C8k7YnUmUl2Q5g/yb82G57urckII49XYXVzL
9Qw3OI4Lg7lkHtr7VJxAVMjEL01aYPg1EkqhBq4TGGxqIt5um4iAkiXFl26fvZzExyc05s+GcTem
j+4ETOD6VEII/XHnnYAR4ln0YyxlFyM7JEQnGB4PVUEMRczV4vm992fyc+VqhF8OXJhdGEXMitEX
IDojkeGx8AVgp9yivsgG2LIvM/ri017a6a66bIMf24DAvbqKX1u8eMjr/VkqwbjZfrN3za8QZwL7
57sVFOVOxY5h9tYu6MD5MTuZufmCrtmn839owFZXWGowSOWNHbbrjLH3Pa4ohbQheud2rmPR4i6n
uZI7Rx57MXrI3jwevOnKsn3nXKIRW6JDrv+aIrzK0mHkSGdon4FM6E4n3saaQFpY0egj6G848sIg
2TsYozPonowhvl3xiPfntzKiwkjDMR0sb6K+RFHQ3Q9M8euyGpoMuHSte4vg7uerTtZ7LSOl9Vco
enEveaoZUdkuBMM3lJYvG5jXQe87FsROpiDNhonJspZa5R9+Jq8fcM7Jd+sAte/FO73klA5FNnHr
PQI00QSGcFg4sM3gFdumNEavE2iC1pMjbHp2bAbldbGrkxZkcJA10KEtmWPbgqQmSzp5fEKDNXi5
QTna/JwjOGcKErQIco1CZ11+Xk9ZUW4ywd4983YHYDSbg2DSXheimcMv8/k4RofuYCGK1ZrUHR+I
41WF8N0QQgX9hct0JWckD1NSQvUJPpeFvXhCnaIys4ZXaRV7+5jacTfM9lgjmUUb7Qs7KkpJF7pR
PhOE7FY9pfWRfuBe2PJ6NZQjTZc9mt2l4DJiiAEbRsn1Ml5G2kH+z7DKnANLnLW/Mz994DjTJJN/
hSGZLqdMEVWdUpng5LizRR0DwfPJc9zfwDm5BjH2l14SyfydAtWZwSXIsjZXcqr8qVSP/ruG/Z7L
p0HQOUq9q/3e2SxumMJLg8W15KtzjNy9zJSBypww+6qJmS5j33ZIx9Igq+mXpESf+Oq+a0sh71ag
rwrP5KslAG4nlpff324vVqjjwpTix9xSN62ahmCaEPE3NJuS0HCstEvycxk7nC9GquTndA2tQKyO
VXflONBHfOjF/9QLlFGcfJycDC6kJpr5egEDEPC102l/BfzHZRiKGHzGO2eHUOOicPEXcPEBKlPV
wUnx7XZ0Rc8DjPPYdYm5p7adV9MAWu+r9boWgWEWdf7stHEqj1SrGdO8OmccK5rdeW5e8iRzWndl
qzuhpjTVA/69vQzNLOhHHqlOuBtBdlQLtsFC43LGnmFZ+h/AJnw0b8S+A8ROapISW9p1tfIwPSjC
shpT1Z/4Spiq9MSZJ7irokHF2pjmxNG+cSt5BjTVvKqoWazql/Yk7y3HhRc619jtN1SSXzBCg5ZI
6Qs2syg39xHTPVYXQgBAEg1E9fSkDWv5itOPRSe1sd87KBTB5eq82xIvrRPYVmQIp9oydtM5i0c+
zFFnqu6D5WFm4ZzOXHSzkXMuowC0fXfzYkAkiOt6CU+ElibYUUH+jgKifwt8bAZP/9K/1t9gAimA
W8Ltv8Z1uTBYvzcs716Hjeq+TyzIG2JRtS/NatbjgAgFukFpimQDkO2n392bKZ9s03TOQNu+RaUB
Ope9gVY1zRPVHil5s0ZUdtNpXZ/s2EBK0ja5jt8tqabhEe3RC5KBfl0tctGkbj81bAvNAXZ5oG4V
lt+IIBf9FgZf6FIgDZnFnLKv/y2pkYcJGnzumJRxYZTDam8uCf1f6apwPscM11geNORp6snkRMRS
u8anaA8uDM1pbkUGtrdgdvvvRxKwQ8UwVSSeqyppYcQXPih/pQSZyXAyWLICuUC0v2fc0cWhnpx+
W0JO6QNE50s+zTNH4tdOa9RAgNmuLyCKP+3wwUu8OebHBgtPSgdfHJSV9VBwjhXNNTG7cv996D1Y
Nc/ejojXOT2qhH6FrcIkkkUcAh6UGEUhfZ8mMtpsrG3YdZAC3ZVoAUhl4+TWkyYZRVpcknlHQp3a
PwMj/4az+LinPEYc3rOmnkCMGRckhLXYVEmD4P8YuvW44QwO6y2mcH8qBvT4njTeNmBbImlMOEW0
gF/EgXM82cpAxA92C/FVOWNIIOQ45OKHyRIaDpTd54r/wwdfBUTuEJzt3m2qfYk7SyX/LA0aJOud
ZS3DltDkvrPvRaijyjf0Q+Auyj5K4NqNYqKVOm82+CM5b5JA8ouacESgXEOxyYCp7YRbE6KXdfVE
dsWrygpPQyYrA4RE+znFqqV6CyypnfWLwDbtRlLJi35K4EZbXnhR1yf1qyXOCporYaEdPQ9bvek5
oSQc7hQDHJfZyjsizC1OCGgZP3P2rmXsztw7/0+s1xBeAVE4RXMwDqFR4PBM9TohjDI7kgA+gQJl
3/nMaUJfPZvo4UnBnHDA7opKXmQFeQ/HdfJHeaGxskliF+DbK9Oqvj1P3CtSqHepJRO0E/cz5pzM
SHpGSpZzr0HHp4OcmiXDAbHi16D/4TKKq9zGegDhoLmdYl1w6YzyB8HFPandWf4Drru3NVsulzbi
HmhBoeGaS+3JjsDyOCNiPuWsp6n6996eWa/coOiGFWrv/xV2cBAn0LNCufXV9zhJ8FaWiABnL0VS
1zBXFLJgF23Orbu0dJkAiWuXe8yfYA0uCuCMBesRgyGs1+MDA546I+wA1r/b4ieG4i6J0fKSE46l
Ehr22HQbpOdJZC9LhxbjjLgK7Eetsh3k1/+NBjrsknI/Noye+msbs+1nOpZ4VZk5jFxkcTIomgPq
cyYZNqHH5U56lYfQpM7Mf940FEa6IdxO5ERM3hjB45s9iiCXrSnncc0n4Rd9lAPgtm1Q91ad6A0v
liOSZOWldQU/h/6joSlDF/o4uUdxNnSk50JJ3OoyR0/PCZ3z0WnI6PO+BFuwQH4312sXC1zug+LO
iOB31cxoAmbk+kYUL1ryfvXDkDf1SwfrjKaORowLsr8lmVLUvP04tHTex7zM2YSQCs9d4RjHToj5
j2lDUztBSDK4bnW+21G+T0h+m66mnW54xjB864dmQee1YYn1mj5A2UmPwKaq2hmd//5vZv/qSdBb
Lb9P+MtuDcg08BtwcSe20jiXfpjQZMnqy63yAVlAcvUFY5UDF20yAgIHUs1YSclXwun3+Q7C6/0Q
3TNNnwXTcTrrZyLdQXMY6QQmanZL5u8cEv2kQqoWMvsEwEd2c9Bvw5gbf8Ei3I96F6r9t0QRBzNH
J+9xiZK2gTjN0bUNoxIE7gOoiAws0SJgzY8qj+pP96oqj70sK2IVkoFmkHN08xkCERfiUO8sAVW5
f6UppMbvzPMzy/vd52KkuIPqKiBcP0fpJLnEhUFtnhql6/6hKV8z2DdAiFWrm2R8JR/4OjcvePgA
dZmHnC9TJJXwkA5kZ3PmsOZ8lijkdIb49cerdyHL3yHSfuWG6j7IK5dxcwpE3D4yJ5LYQ2WF/ezo
vhfI+zr6he2LZkzwv1jlNbECqTiTSFSJpp47olVFF0LJGUcg6LTwIIxSXXr81LWdmPJqbnuraMex
LGjuOkVLAEg5xnqCYEZayljm8P6NASAMJsQfn9wYs6BYKq/PJ1wk381psZbhJSJwwTamOr3P/u9M
REXsyGRF1DiTYvvkGuWZ6O17iDV9sGPasnQuCkxJpgoPoumKi3fWbzNpCka1730lNLjtUnJR0J/b
nvXvdgs4ypShy4bxeKTS2vsSqeBISxZIH01EZodd3D002mshQaO1ltKCFUW9lqfHyf/QljLqcJI6
tE9LlA9rTub2jHY9fcI3msIL89xSD+X7qH/ulISuQnIReOXqBop9RVLxTJnLqAH25TYGt1xvOMwj
KiKpm7yRG3jJWBRLMa3kuSkv1DEQa3KBmbNi64MMe8pUx29up7OsDYQzIAyEWFokGSEXtH/Toxe1
nxm41D2Jvd1z22GphL6qe5pqvhUxZmeB9zzWhNnZtgozNgGUnOuW2w4nvOF6SAz+CpV50BcWEmGG
2f/eXJ7kPuWeQV9OA8tp4An9yQnqUuudz0L1pSkQB46Mycf/lD5u295+1H9kH3s4MiB1FYwTbLUT
4VtLpP2/EXZmFPfV6qnYc64WryxJADLMesCYjEPyUKC2Oh6TKgCcimnnsCiTB/fN/7ITG8uKsbOB
+wlkEP2fq39UYun9xc9d0JvhEcyJw6FACcb2Pi19il0ad8Ceb8JUcu/px37KWKLpRKqMf48yGqg6
sIWhdXDuy5e9GPK+GWUUlnu8giGUb285RwbtcnLBXpFdeHL1YHIUfjzGpdL/sh4yKRWGkFgDQw95
HbJHREZBvYv5IbzkRkGWBjMpsPvSgXxF3T90bo3Qu77x7npbcFSOHGQZSw0S/akIAQbCkSj2cz9h
6N+M9zTs6Le8aB0WNvBCwmTapmczfbU5oiqkItQpsng3wmr0hiKNPfq7sZoz2Y9oye5pq1GZFrxW
AC1pCoHsU260EGMISITUcqG8ZBumYv9SzOt2i0JKnO8DHSQJaI7oSKo4GRG5DfiY+zXtMHpbdY/s
ndTqtJSNEAIgrhwiwmZPHdECTS/qz+OdFC9g8VUQbAo6RPxQLfW3YEt3MVClF1/wPif45NIJ3cxP
UqhUTlxzaD0hgoU3wFskD5DoezvO0yPabWjYmVN89QkKgOVC0NY+ARPSrB4CE4699b8BVYjSLLEG
bWlDa/v8dof8ude8DWR4Q8ooQi034Ig08gk0FoUWz82lG/nweyb8j1RSIag75gUEEIHh7YUOB6Jy
tTdR/wiw7kdiuVdJCBqnFwf6HTRHBt5Dgdh+PjoMD1X/c0NvqR+a6krteOatgLxDV9Yuet73wAVg
BG/GX9tMCVE8GEnpROQ4P99hCk7YvwQGUkMSxXW6HiKo57etcbyGbKZAKWCiWA2sOjbK/rNAboAy
v5u4uoKBTDYIuETz5KDpyF/bWo7Sc4PJulOeyjwstW9NDoK13G3Nt9yoVvgKMRRzFbj4/C/rkaX+
GWbzMoiY0AqV3AYBWHkrqk/ou56g3yHruJBipDQ5XaI6d8OzksAmZgC8xO8wknINvlbXGmgv75h+
MyMvSi70lioXQtwaz7Wgf3SPiHBsNjviySl7E0BUoTzhu23t9j0X55EfeeBhqCmgemqFM+J/LEvb
tE3+5CBp1vFpi5PiryHYpbraiD/7/QbXeBWTxW0UEkYMVD0jOPrdvy6/7N25bw4Kbrr7OYmeVJT3
3KCQPrjh3Xu2RBH+r0Z8sQrz0zlkv+m7WWjIOMWZD/gNNkHrcALpGj7TVlHrqz7ueFkr6RGCOq6r
Y4YsnxXXgcO2uTE7QJ6PtaaFo2AnjnzcSkxEgRYM/a4rrxAUVdMJy/NUoWkXDhpA1EqL4SK0TzMU
liHw2Grz+aAMeaOIx6xIpnMJ06M+sZu/eSjD7ZuDj8ZkobIeAiXV5zCi8zCfARCVTdU1Wu8gQFlh
/dR0gxiD+JVJzgHxKULXLll9mM9w5lX9KPtO/T3eyN233mUXzXnF2Zb2Xguk0x+5fWFaqyMtYj4v
CYPu33qSkwd+pvK6DSm4pxMP35SPdYl1ve9qza6+lPatTOP4IGrl4s7nq46zL1PI9Jvkhb8PZ6YA
2Lwf/Cq3+dVlKMLXOrKLiaeO+8kcb/xwF/NozSmJTB9Nh+rlKe8IgbIFf+TDHbAe2kzLMSL1PyOx
31A47Ns2d4Bttr+OBEfwRMXTBOHTv9l0LhjL+BZ59evHERLyZQeqY7nd+bjmeljYGSbbsHaBcPf0
0Uov/qv9T1JFz9gR9+Yifzt7sFF5CjruV96knMC1mWWklBs2gD9GImllJijJBc7iLJFSlvIuR9Ei
IksgUGJAYFeIlrPTVGQQBpD/KVkUc7YscoLSW0v1P3KXduSZwCCubfj3ZqgoluCGxHZiEMnl1u3B
j1XMdHkYifdO5cdzzmOc7LLmV994eK8zYiMTxIfKRbaNYiEq8ifaQiCIYqPzjtCUHWxnnP5iQpJa
6oZUEnTMKvL0EhFM8wJutyDuBgugnqmkPQXFaupMCq+qEBXdK0wZIZow6cJX2JXY+CtbHjbVLJOF
/Xp7SvPY2QKBqTbIukW3wIIvsYwY9wpJIxQp2sOaOSwqcweS1holS3hZSWZcAyTX/k2xfNUDKPbE
XNRqhcaZn++1JNgysN6WZXWXLW9ySQsrVxTV7hemFwOnqpf6kFwnDx94RFPPEan0juY1mM9PY/Vx
fh/y9ndU7c2lXhKOoSGYWBzb6YAmLeUqGuy3kNRrnyE1CpT5hzx2Bi17zHYf7+Tnc+07tMpUxntu
Co8UNycnHkosEhOayuf+/K/ZbzEh7YuftD33xQJ+5GzbBsSWjQDqQOMG8o+gJQ7LQmdw4QzYunON
2wQO7TDTSG3RLSeMCHQ+Kz4Dox+7Ug0LlI/rNsjxxcrsHGfiOGqEc1VdwG6m1CQ4ABAQ6tZ1cn+J
aoDLJ49bZ592sO7hP+z+XpAa7TKh/VMYSXvut/6Yn19xgm83LsXdRoPon1finbVs0D5X1GimyKUx
Fb95Q79oJW199EYuN/eoavfuBFpr4qunJ7KjfgIDRWlW9ft7az7Go8PWDcns2oirnoAQVH2Jjkqg
iFKJPZ2MleKHCmJqGkT/LUcdwgWnCjLe+axoJJFKaRTT5i0btzTKzYAQ755Xs4cWq/jOpoQsmoUb
fCS2aNAWRJwYjcIsuOsqQlHIMPjlSfTlCp43WUQh49TI92Jmj2CubgaBGkkmQ3P1FdyejpXAUWBJ
Wekt0cwbfxZMy7M6R4qqYc4ppKVSm/KyeYZVZ147G8lBkC0CpBQXRcIhOaHJuxSCA4KPudC5cU44
PcvqEbz3WUnvLY9xW+AHQ9TECDSg+7Pmf/Y3FwgoAB99Eq6arREr/S2FgV2N+5lHfjfbXefGwpbo
vqsDvyB8DcAaqhk0qpqd2tml/09FFPo1VOukxl0BxyqcZ+Mxsi+0KyGGy5FLsCVPVVrAbImyb0Xb
Am+U+PhfBsnmwQW7EzLklGIuRBy+EQiddOuTp0R0DdfWEoRAC4Qt9kjYOSqVwNurfHhERMdzwIoX
SSo2uXt8KrSdegzouBYq9dFY1jdk3XOgkodgXVuHr792uCnv4YV2B7mKfX8mMkLcoxZ3+D9XR9Qn
nCP3IoXdLYWYTdeUSEBDj4ai7FdXgILufGDqoNAoDOKJ9+q1nS+uG0YRBo3fF6rGiZ/jmUP+qntM
AaArvcwJKNU3oxtVBQZR4wQF7085UUOplamPBEz348THbw6NhxUVjyHIiGV5OTeDVF1iLEmFU3VO
wFUvKCkTJb3cCMUS0xFGfyPzFie2Y9nVLzvmplrNQ0WNOZz70Edswr5VuT2YIq8iVN8mS1gKbiCi
JtDzflAf62967IQGzdB6ME+eeI2OcPfws253l822EC5UpMoXgmFp1PcRX9sifslBUX1EJ6ltygH0
ZBs+ZKGel69hSF5pg1n4Rb3AiLKE3SNIqDxFTFrCpePuICB2nj03tF8IDIpRffE5VU+Reo6fDei8
BcaK8hghcIxpmTXAa39nQJDGpr6mQSULNN6JBNcSkAZlm5YRjWzdOuj0MUxTTSduqHfDIqBwMK8w
s/Agq65fpXHBoAt8hMbSby0swMAgwz08uW3ImoU/mklMZWseKSKDqSiqAQ56X57uUzShwRReaLrQ
owLkk1pjs8J4esongCnCcPC8viRRPIGXd7I0QSHi/zz0NS0t5X7z3e8OfleHd2r9mYomlGa8OI8m
I98jXDq4NRMV6IqtupTAQ9e9KxGJMAkW7LlDivh6bEXweU0YgeIgDnanyBpmrCx3TcBDpejV4gR/
cAl0wAmdjdH5B1Io8/qGyuWogcI4Y2JYiYkKTa0wkAjG94uFpTxsiopOEcbTCUgpPvFIcWKfBmbM
qzQM8x/l5oVWVra8/S7vC9hevYWtkwlIvIOrn+t5vmNrmAfCd0nmZUuAT8LE8Ff/asRzLqI5pBJp
0wmHjBSaFemYxqPy+XWdkGc0udGXVEU0kTREL1Ugeb1kr4EOqfIQg5gZ3TjEFYBSr6n3jecJ1/Xy
hKDWwcxIQPUr0e+Xs+YDDsAoC28z+vOnpgpcD06C41Djm7P/h+aBCxDNeaQw/XKNR5uvwVORjsrd
SppDHXxHdLfBF3j+bGxufuymvm9YRJF0fofPClkkfrv4LbN8axAlHDJG3g4C6R0Fb78LU0K/VCvX
KLecNglaPVQmMU7/2RMD6xhQx5/5wJSECDYKhjbuYFDSADoz6VwGtgZertA4bl844Aqj0mJ8rC7t
hw68KLu/WEHB0/Y7e0hXmOI2Lf2E2nTSnHoyCpRPk35zUJvg6emTQviUJgo02SSywMevZZibU9z8
JZrnT+eA1ol1aJJEHuq7F49MJpS+hKsx5OPKb7rsryHR+0lmhogbLAe+sO9bzb/02xdqC7prMCXF
5TvW8POkNw3+iTWU3MOl/HNNhnfMHe+FKeiFPlWLb/kCqt1Y6q1svG7GJGg/6b59Ly+yuwmwh+Tc
u4DJR9T9UTUwfFF+n/dlFwQEr4S0uOTVWm/dlXvHlHFCXcU+SqATi1bA0X7xQ8MgSAwzJdoWw8QS
7eXrKdpsMqrsP0+40VU8mjCX779WwWyHTdiBDSaYPMogVEvXjVvhIy7sBnnAvqtzI7mdTkEyWMTL
W8BhgRZiLO5wagMhb5BR0ekr5qVVgoxIO0TReeb7cdPTyuxAVgoBEVILRr8+spkUYnyX+9CmSlV5
APJLxl7O/U0Bx50pjVr4tqmrMJmZRHqgfI/qj+rtqxBMKjAZ8rChfXw5wDnelTZIUt90Zh23nZj+
Qu8fma8vA9vivKn8h/kbwX/NQ6MXy0cbyZGIjQ9uLbcEh83QDoLbBFwYDuv04juBfBsZgsLDmAxz
Pbw3juwBirnGbNwkw2Sx1EVA3T9tRB7wT2g9DyZLOeu3LzIsu/N7pzOOnW+fkqgL8ZSKhsvTjBXL
byutKO+9XoQbzxpakVAVEhu9Rxtkw7OpR0Nh9ken9kklR/Qm2AybIvZYtY4XsOoWwYGWO4yy31zI
Pxf2x7ZC4yGyhWKiWJILjJ34L6kZ+StYwbYJlD2oULCoQUikEGQKfnX6d1Bt1zDajctD9Qmog9HS
+6A2v2PKup0tw1/7IsdDLx2UXUmM1zjCNdqSvFXM5RBB63K+RIZUizsHxo/lcWYz61OHM1KqCuL+
08Qzdez3VDbMEWO6Q3GPCrB8gmbaVZsEAgNIAhM21+XwFqX/80W+eKMN6fw80R1fd9/BJIR7bxVw
WtPVYzNgkaOW+DFlPl/AjFfjtFsN529im/lSLtwvafGP+2M4BP09M9U+g4UvCvsFWwvyTyRmzpaj
V4hH9Vac4Mjb49/5XeDBHzvekSGSkDNR04xWIjx4v3H6PmocDZoAoMv5J3fQizPsKTniyyX3FExN
yweL29Y+us7XMu8VOP6i7hvxVSr/cQ3SkVyB1hp/7cJtF1CNWMVFvSW/m7V1mS08OfaDAbw1ave/
AN4pLGSVcDrKxQQJoy2paKzVqYkbCA5YwIS4cmS423kIPGFfg1g1fQIajXECyUKxmp2Rma/qzzEE
g6cNWwA8GJR5hCVCz/nW6UVOvVpbWH+T9mXyH0K5YIZ0oW7ZeLI0Dc8U0LEmX725drOWPpc0EJa6
nr0T7nKMrTsd/0oHIxxSHWsFgO1i5OXA9GT6/l5ffDwpgicni28N+lSrnDRl1c5bUUIG7TisgZwO
g6kumKMIkWhhq2EDGU9RwpQFKQ3my3+04AqkTgpYazyIw1e7kz2YxJ05EHrcK7ygyL7nYYv5Jrgv
MdN2TrjfNjYwXitDE9dIjixza9/lCSqx28mwRSHq7tHZQMTe9CAp7cw0daH9C9HhUJkHK8iOFRJo
hlovO4xoM1mfhAeS8AXKCzJq0L17R1swOr7byzFba3mMp943HL1tnZG0C4ihWfUwgJ/3hbimfeUn
H3Y7muWvYzUs3X7nwauHHMjxIo7iVv6RvDEl0pjgfZ6k7ycBnOhbIkCI5t6ZmhZ4GMjrxqsvEPBE
2H/Gy3anlH8rQFCvAJvzEJlSkAU4AbpTEWEnkqQPRNEF192OWy412RWT8o6DUk1iQLPxMLTtBzbi
QWW19lJeUp7/XvWF/Bt/fES1KbDZIAcc7ibvFWYlM4woMbnO5ta/yg/2Exzv/9HkyUW+z0YYWMbR
+7cOWRYJqZdPkINOG8kmB1hqISfArEDE3IGFLe8AY9KdodYjtClp/+kJ3zbR6RuJxXaKxBrYGV5k
J37m57P4Mm1tgtXxl/FjVc+4IsDva+BaWkyzHRSw92I4l4eyNIoimfCWYjjHEhefcHFzZZLpuAHV
wSWPtpZ+wvwhEIAk6WZ2hyI5dl1OV6MCfBk8MiDhMtBN1eE2CB4e1DNQRpzz7ILECWAU4hv5dgZ1
z4yxrQ58+KgsMxuRYEKjHkyH9uLQHVY5AoPSpQt5W0vv8Ixz+5sDFpFOCRIM5BzKSFF6+0EhmwIp
0rvhgeSXgcL+dPNBHgPPMjsfrrF8GapZA66fqC6Pr4ETwVzsUjvtVOBcH/mKZJXfbOmWEpZl99qr
NLd/dhStdZoJf5VtozU+zvIHF2i1h+MQAo0Z05Eu26wIWeQm55Lj/hgnj1NjZoZhFj/gjQoNf8tY
8u2PkGGjCE2bGkxhjXAqK95C3PZZ8I1SdVrUJJ3Oqv9RGTv4M2/rKG47GSedfa1Fj4YjkRjQ4dTU
Yx1lAwHKVKTXZEqM92L/qxjEr3UMhgmaPal0RsOLHEqskaJuAryD5/dO5j2WA29RJkaur6WXnyEb
Bl47meANw6G2DuSoEgcTuaCdq+IuVoZ0mNLw0X6W8gSWWivUGpRMqT+yPC/qLdjRJJiQwDyGIH9r
q6aL1QPP+JqF+XcHDc914SlPcYrzdaQQCweVLK3Tflah7TPd1jdvx/m26SNKJMIWiECKRk4BPLNk
RY7z5FWDMnlQp2z54ztBUzLkzO/UwLYjEav2DW3bMiVkgwC3DD7nZOFqXCJFSK3/u9jPVWe15LZH
OLybBTqJCdqQWfQp+Q8osB7+4XAxueeFkEGytGcsDRW7gBmWIuSRpeAnoIvUARJl8K/+ElecppMU
YSXA5h+9/C1iDYx9kv1fS24fGyXu9RMU8iAft8G6J/w/Al79Q8ZP0fICKAm/k6/ubjTdg5vCfvEp
DaXEMozNlSXtvBPD/6j7icMv9dZ0ZZbSLein6d1NNcREDSsJVUB/5KPhRCfxCotHJmcwbjgTexhC
Ik27zLEiDHm0lc1h3tj3voo/T4i4GUsLxRUknlT91EihIG8lS8xOVTPS4vwH6I+deE6BByozSUi3
85XqTKf8ina9cPKkk26E/XRQKhIOpYT07PIlZlgl1CAj0wTu5cecPbE5LY5goO0wvK3IfnQqFrYF
0sMnVFyx8apv5RbzKiT+1IaIY1JLHmM5ZBsll/U9K2bwX8LpV9pjsNq4g7z3l9EZsP/2/otUkaxt
ULVTxdei8HHuXFv4vnrvG4cxYVq0AP8VXckNtGXEYd5BL6yBrrG5KflQ4rKX+LatyQE400z7ANOe
kcykGy5OSsj3G2ZeAugFqkIgFYvaCmdpJe3aqC5bdt2TgekUoodpWcME8b8BbrCc2U1rHP6QQYXR
OdDAZP8Oh/vHDZfKqXS4fRSD5T7VLJyoE6Z2a9q+9IAR1Y0upWVSfrv9rl5wLfQ43/GErG1GEi49
UvQFudCMQ4Y2pYDoAZKCk1gGQnsU66/Vee0Y0x1rKv3LxD9OUj+nFIsa3RpXtFOEs4zhwU+aVPfg
gjBawpkdPzbN2ICISSURdBNZt810aJ1wj/3QPjiskxJ+eQxGIWYmQvzQMUC83T4X1F8A+na/eBe7
d4tiCEA5zaAhyAnW50KCr1uq6moarzXsbA6bdm7Q7oniCeA50ajvrAj2lhuL8A5kUjKbbNuBE+pg
w3NNWGOPD83eALkRm46PPvBjlZ/e5rRj8h0GQIpOb+lNFpoPspYJXE/iO5SUktWdNsf3nGQFo3gV
2xHBR38pz6jJv75q04wytJ7QfDsvcsD7/NkfSkx97VINYulx3oKWUUN6D3pToPpd/g9DD0aDwjyZ
i+9W3HbzBYaqwPA071wxkgvq81AYW7wRaZ0ah1QZqlSetxAELY783Pv4EvGPbUyrwMYUdmF1ulFu
WD5F48/iA51cu6BjUSEMJtCzunZXmsIWdonUx2QJ7vSd3hR7DRmI2k24UO7/RdFYm5PDe/h77CIh
eyqonz8TxvOrls4P587He3xsAke4mYrDzVDGhCfibfOmUtyGQPMkLVh/tGHcsH+5IwIZ/9mpfz+u
GM4UBCz4xoyCDgTfaRnm75hR5RrBipWDP3ShxmJkqgzk+lzuYp54fj9rjHuYuTALrazn6RLpUNd/
KzkkQwttXNrXJULcsr4iEzWc9XjcvJixL48SpMrh4VYuse3n79pLryVLt3oLn0XJOuiY6hyrY3cj
xMe4VQb4DWpwiCk3qVcaO1q8fBlsTVS9klwXaZGOwKc68jMXxCOvkB60Ep5ss35n3rd1HTmKnwiJ
VABU9gpoFTJw7PgZFfBgSZH1V/3EG+cr298IuwLIkv8USZK3PSvzrgazAGe+VR1EmmNcVhaeqNpD
tMdARRo+hL+mZEPKCSlZtVZRbW7j8Mg2mpFTKD02lczmxTq4LRH/F0n/ah/1BEMLGVqtV1PDFzQ5
ogx/vay/jlKI0THHvEA0hWBn9i4Az5pTjfkav4UI1grffpnkzGXH38cmNglAigZlUyPsGH7vHWUl
jOb5ENdRS8YLS3utUwEpjnbaMqi86WJEFmi2Ly5tx+w1iqJsU3Zu7hSGhgQMwjYu9P4qx5zCOIae
jxqXr0Wy4nmoVEYBG6tZ5o/jq4rwGAYDuu2mTuEG9vUBIEqQrFbdLK307Uws8xN3zBsRnytIwVNy
ro9H4vNf22WWz5cR1hUc19N5LU8qggF3XEwqkC4/wHnRaiyOm/gDZi3sArJutfZz5ARInx/b81Az
7ObjDoJWlfzp8UlsXBmsJKHWeqpg0vRAdB+0hCNU6hBWajBk/Q/qrDHhggzuAkk9kJPIjDzrkJWf
qE3Dqv8Fl33MmmDeTK5yhfw5vv/EgXEq3YCVNzNuIgN7obQhxPRdwa5bWDgYs0fcqrAyEarR9sDy
Q2qDmyYQULajuTt2lr8fHu3mnxj1N/69JXbpbN1zonL1uQO98UmcFj2zf5MYj5kx3UslS11SaiDo
8A0C4ehPffikomomBPYNHPTsmre+YwBsVOWVnWToDQXuhVmM/A0QGqk4VX15k2DNxL8/krobuI3k
4JORo08mHKqy1EKy2eZ6NEwTZk9SsyLw7jxberuSiIrDWjAdutZtMTOykPjdbxAujWafYViqRJqu
awwZ+cyJNZM3fnnl1SWgW/k+CznmzerwXrv9sl1Jmml5LBHc0CA5dO/4r+XqDJoZQ4uymbYT2O3N
h8BqFcfsJZoGpEAitkSav8dKJGKpGcoNTYq7h1pI2VgXJpGiPqrwM4lq3b0J16wvjVGiIjAXhK04
TR62UHpuMlsBJNvqYFLs1h50PP+jHLnVJ5h7aSpS/tHF16ydNi/CQ6Vdxrz3jbGmfzAKU2oCqgpo
y99/c6BM+4o+ylIESOJVcf6ak685KB0t2rW2q+OR5a8Vem9iaBkRgVnVKQ8QT3Eo51gnqJdLPfb5
NjeXjl3IKLbHu2ZqOxvtmNX65Cf8H4ZgsziIXaHqoy56Lwd9WOr+rm51Dzixu5TKjr2z8IJThxRm
zbh+lf/Jrlj2r9qgX5CWbW8QJtDFzhwDIklCo1/R0++ajb1vsEO6RSCXm5g2UmjCSIsYo8kxslU9
Pl66Q/UV+SXLh9Rtinh0rTvovViMwIqNUfzMkF61Rx+Ye6MMMEkOGxeRLcbsvhd91Fy6rVWeugze
vL9/KISX0UsTfr6vWvHD+Tq1koXagHlhtG4dCBe7mt5ME/iZ3bpzq1XLd/kqr/I1GlSHjctQtK/7
+yPUmOFnLyT9FrKisY+41aBCgwyx4fRJ2uuijfSdX0R8JHNVgTkc7w2aWKVIpCrQjdpCkO24sJcW
aNM3iEqh6AwlVOKRI6fiF3isu632Jg26AY6nHgpNPEO2zQfZgkxBukPnv1mycMv2VgsHngzdooBX
cGnjcZoDRnSlr6kR5uMTj+B6VryDGpJH9cb33agSgldYJX3U047MOcIGQ7IojCfB17Aham0wsWVC
EZvGAM/KD+5MlkwC3boc69Z4htBqwrxA5k0+tNp+tWO0uPy2aHf3+2tIDx/KUsEV/Fn1OeibS+fy
sZnHmemRicr6/YbgbiaF66CGsSQqdiu2fEjKmp3JOcqRNYo83Pay2THHHP0eniPIVIRPeqXH2tnL
U9zsnyuEvYuXzPif/GuX5iXnSDuqL7j4Qdt68RFon63VlMvOCmUxknZd28T+fChGAhFhL/DKnZix
UPt4J7BjaMPPRQ3xoAG/5lrvNBkYaR12wxtsVRp2cQgGuNEzEl0gpf3MmdWr9tvcuLTb2Yx6nTlT
Jh3MMFwJiHjlfCO1N90nkrIQxol4WCzUc+5Y+Tfg5vXVTD4D9xKAZVijP7tygyPxnxU6rpxLYemG
3oeK1WKcJRcunQuH2KoDlblDbGP7MgRR8x4Rb2oDCrVA1lW2swvOXH28wQgN1ZaK+etu+veAhmlC
2qH7PVUNR3JbceVqG7ojR5PpehqfjA5KVQ/NkAo4MFXc0OY9YSmAj2AfHO8YmgdDRjwbw9XKBxXO
aDEEmJZ+sal1a/5oXG/gGVJ4r+9ObSWxTi6v0VHLDWDP/5RbZjgRIPyZFrHb4m3CkkCcEVYMBp0K
EFd7kSMh4BpNBBWR2GOMVrSe+JOQiil1R6mhUUhb3d+u7lPe7wYSgnX6/YdZX86qdlax9pxufWba
ucgtxV+RjOGAhVj7zDj2SdTuztcL3mbYK13Wilsq/PTeqipT/uNHDNFsSK78y7CRgvAsIz34lULP
DOj3IuM3/ECp/fl4lBNY6RrWb46UZzEVCFRrrW25qIjGAuna8ifp1fGuU7fl1Dtsc1RaRTKosTLt
PSBB0fAvqr1bdyS9oZgORvn61Q9ySuFKIFf0WeY9u/PUE415QSNhWLWWsfuo120KadNHBs+ySyQP
3se4vnmWzzY7FeHMiF5HO/puE1Xc2YcBtPiupgI2IJLob4unvPThoLzYcdqZ4Bt/QUMhz60+0g6+
EPEk2RP/ttKSco2sGZv3d9STqb06UfCIVjoy39HPjtoyqbxgBhi6nFZd2qOqBhPZx0RbBkqSZv9H
0dRcgIWXdEu0PnzYAiioVKRWfpqb51qvFh+C9uaTVfjYgPRY8P27cq5udKPgbOpOC7RcJXdvsy85
xyqSL02fiKa7R8wofwKWT8gV67Fs3DTpA4okIu0m6VvlO1Pthnox+dHoOtNwhasYVvM9nKc9FZQH
XVyCsZNcHcRL2iTRtVvPu2zHNmh3fP87Ap8476JfFl9QIs09qILRbAq0xk9XQpvcHRawn0wRswQu
PUglqTr/PHD8MJDjn4TpDcoMTPkSYFaQnj2sSgD81r6gJ1ziOIvniM4xXu5XbpV1U9Lr103mE7rs
Kh/qLcPuol7w+4jk0ZhTPOg54bXQnMHOYGXNpHhrBUk1Kb47GDpaVJiWA6zcmY0bWnj4hjO61ZmS
8EWvYuUOsWF+vEaVpuXAoPToV6WoWcaaktuwC6NKD0SQW0bg9josmjTPFAXdsA7IUb6hb2XyFsg4
iyOCWprftii0fvfMtlfwgxj2SXYkbNYoD/TidtrcK3//Jbk8Um4LnkWMJju6vb9/PMUriGpAU75N
GbJ8hlVq8lnZK29DZ9a4l5Ll/MhaXZlMS11OTFhsJO9D4NwWZZRMA/fMHE3AsXqmujZaqpD87BYp
0mEPgPfu40K5rMIfsy+SQN4yQCupO+0M40oY+pfdilTbZV3VZU1Dfk+XxV8z+jRHGg2PUqOF4wGV
/6RAXKeGVSrQXbwuUMb06+ww1xDJTrnru9Igrbet+V0phBWz41E2EvokS8f6MM1YBYd9hHNSIju9
3U+mjioAG0d2huo1D5rVFJMNEeQtHGg23l1CKF8ekY+Xhg7QjM8FFy8NxO/Vl6/nCeEB9zhQE5ZR
tfM8ayhrAVcI1IrZYNor85jTZT8/Q3SBG948DiYp1ds4d4V/PFc9Ie8wCIiEn4TrEc6ja1I5G4jn
ITsh5KE+r4grFwN1JingPmu4TMUNKOCTMFoXE8kHSKPoGC55fvFjrdbZPyLNsWKUcLlgU/H7lxDw
Um1BgTep4x8QRkF5x8giA3rn6si0adNHfdi/BVEFaGwABPXphzSkjM3gnJD3fZ/U99QWkVsa+ybP
EdDvR51yK53CXLxd1j1J0FQ00ywyhwrRhsJyvuUyBhzrjHtwyC/iMHkmVfHhRGYi4Tn7Nk7bp0W0
4zAMLU9mLwhcgLGnRBqldbaYfzX2151P+mZeASPpzyDqv8UZiVauc3MD9ZbU5yl9ZX+S9ZtvEnxA
wlFBFECWORG0/K0DPEcpOt4p4SbEKsqw6V2izDi5yPVt/urJRcK+zMTe8gHPwoOC2iEgiwu8GlRM
X29aIfjx5AwX7bFNAH/PknwCAHSkFcfjgcZIqHZTdkqqvOAVvrVd+e/SAmkxCTrqAdOHAN2FMNO8
ppUBtOiJ0cVO2tRChhVSy7NLZTC8IIRdFhKG+XPpxKgxT4B8CLlHMSdlL1qzt/Rby5IJCbs0MwAo
XjwdmXxVjO1DtIlMPKulVr6IAKMo2NAhQ1aD3HO3Qiy8hIOHbqFYj8zon9jef+uegbFHyqtKDMB/
AjYPElzyrfmxmBQAKxGfv+RkYSe7vdGYH10gCTPdR9B5MLzwrtNlebWBWzDsUQR0qqlPDPNJ+z7W
ZFWljTAbnQBQM4cuPrOYtTUtnCywve1CYRxi7qhQd2cMfokQqQ/Y0Tsm++J0p+WTHQ07A+gZOeJP
0oglm8ExeZjly3z1asq5e4UCqTN3SrSL+Rbc/vpWTnmPFtW9CIUBh6QmGDbpv3W43e5bb4rhT8gt
X3nVqSTaMIKzeNr6JHv7bBPJAOn3WZcokuhtqzCz7hffQ+a5w1pfH4Bv23tlppVnEoRgGVyVStER
UaCSnAi+TPburs8qLny/pZ2mUninHNnwYHzH5KBYWAUrKj9E74E/mZrCumXoYbWTXoxfAyJXr8hU
xBUKl+eswgEELlKM7fo3ZsTz21fGz1Pj+uecg2f5QJOM/vNxOD8FktBqt26I6nwkqmeorw7/HL3V
+PFAY58YCh34qh7AzypsuF5+zhOFmSKwGE4kwTOCdEmavJkKqXaq51US7OzbeezP8dfiShNAfxt3
V9H66jZvPlITDONOXWkSU6XXspHtJft/ev8Q4+oWp8rOI4Neg8smtc/dmBYK4+dHhpxh+F6B2lwV
laj81d5ynOrLIKTni/ZrickEBIylA3BWfWjnZ8kA3xf/YEJjvrL0mr71Nx7UrgMQUWhYjbjrBvtZ
axHVt3fExmqHe5OEnfGmMo7BiFXvNsi+/Qig2Ea9AFG172GtaJG9ByNi9RsyqkAeMRJqZDIgcTm8
BJE6O+04oxLL71SLBUcFTPwpuWnhnxtnpRCDzxaf/Fy2Z3zlRJA53lFnOkL+TVtB04Xof043+aQx
hYR/5CBFpDuVDz8apMNBNKq2Sg4EHnux9TJttLnPUthEthN3sTbWnGiAP53lqRj0NFL4EGEFpULr
J104nHsSGjKN5lGtfV7T92bj7F6uhYmtbXh0pbYFPX5dvjSSTNQsOFwHpUIw3kWr/Df+trsGr1yh
UAc7NlOeJ6iynuqGAo0Xpl91VXFW2vstikT1x13AoPcI5JwutcuazqZp6WCeaMDY3ugzm/9CiD4g
A1YzJx9hivwEPiRWwSGq9q35BWPAheCxsRXpAjfzA1w8w+rPUxvMbVa6J9yWGHdNlf4TjD4QC3an
BuTffS9lynlVyzI+Pw96ofwu1LZuUNrmFlITaGoQJgT+ir0+lV0TjiNFeWaNu6pigaYaHX18Vjed
386Vt9NRlIxAGoZZb5I6hs2/rdAy4gmI2B+MMWkRwPrUC8HV7cw9w7e9kv9ATibve9yrbNxfmd1l
vU+kI3c+xDSt39Nf6L44cQsw/F0kk2GRcym2DnUxKrT2p1WTpgr0bthwA7Q82vEv1xp99rTKSH11
kCrl6zoHl87AC6ZptIXFgSMTmsij5Xy4M0sD8b5ifu9Yp+YsFEVwAhHEVNF4NsFy1/HqBtYG8Ahx
2V1nfD813PRuYyeJPKsYnPcDU+uYID8edd2z8ypEP2pSzf2Y974cwOZmsl8ar+bK8tTnT8AR9ifa
T54qHouQORo7ViGmdUoyoPcdIaTEauYK2fMm5mGXGAsndDAZcuVA4blQyFpKTNJx2vPcEPHKMvjo
ECZDTQIaHXoMdv93Uhj4b9FOMT05z6rafj1K6KK1iUrgkSzB0loIpsfLr9Qqo6UOzTUyOleYTHrH
bxDs+XW12NlvXkpwLpNuPatCys5ZYLaEYAahxkq/AJ2cXbbRfW5HtuP91Jin66J21hiMuVZ1S9Y8
EMRZu8x7CAMCfj/W0nWcrTH48C1jKagwkG5NYqyBTMS1izqyRDYF45MzrcRYMsebpCrUQHwaIjBD
CS8iH1iDMmPURvoF9lvbSQ9Es0YP8nAiCbi2cW/zSaLkKWmkUL6Y3mmbK+v5O5nHmPE/vlv+uuS/
JfPgyYXgfD7GxWIX3DVGcNd/a0kWjLgxinoavew8u23yxw7Di/dSNbJFVSnDqgo2AAyqAF61q/4i
ZNjsl7BeWt828yQFK0I7Sesqsiso1VbKYihoyoDbr12wgiUeMMTULWcmw0UW8B7qNwC89MROlty/
yyiIRNB0XLv2fQvseHuh9O9BZYB3hhJZWmwcyseu+vZxscu/Tk+4N+IsyqkSB8mkFG4dUIrVBLY1
/5By4HlCL54XW8JCGEXvWrrwdRvNkkOKT8gbxhbcQylXzqqp3DqGtUwiNGLs3pUeRQBBJPcX5H8n
L1NctOH6aKYjUTNEb/DqDomo8QMwojf/OSCRpHfSbEPHd/eruI6jcVTbftgCgh477LCRiw9UrMnw
lntjoCd+pzGROgeFpGtc2TUbdcn+YYe6MB73gUEUEgwUHLHFRLZntHKsZEBVKXhuZA6HdwfkYPI4
ETJv+CCoxdbjJRD2NSkEswGErGlUb8Mw2CJFwT2fK9Bb0AYGrfxkEj+uwu4LYju3+VBZu6uV/B47
Fz4xVdurAr0KTn9v2xIzugOngIs9kj4nfZv92Hrv4vnCuPNoWrQ17yhBUCKpENhVYkzE2kLzEVbi
OexBV/myxfsFELHcx+7wIdikLehh/Cf5gWWggOoRJJGSUCzH06JKAaIELq/INnvmlb/5yCCvTW7X
QUMX/nMB+LD0BKx/5MLx/7TLGdnfEi5oeu2asFTj9AmKiW4R5eTyH69G1a9kV0yulRYaY/9ALeZX
F6CzHimn9ms4rowuy7AigsNI/o84czU/pGlrT0I+pSKpeSKuKUhFmpczQ3uf3Dg+u+ClujBvWpSQ
Om2hZooWYU7urdVNUKDF3MQfW0vsjd0tG4ib7rfTSQ0GSxAYG6Oh0fn6eYBUX8X0f9oQ0Ws52JMP
KoVyD+8xnDfn1GtW8jy6mvU8O2pf3hRwKmW5nwdqJ/tXY7SXY2AylIIFKewPjfB1fb5sNbyoC+G8
j+BcGwgfgwjw3J6hQnF0NmT7CDJJcunI5u9ohqpZ+fwxdIhDTJNLR0KOTszko2Gw1oVJ2OqcI8QA
FRgL15ycSON7sfssZJT5i2dc2MfxZBkSy8fTGpNLSVsa8RHJ/B2zRQBbEMHqwAioBi6RuejSnKuU
X2i/naGKdiJZgySrSwFAlGop5a7vYLzx0EZhIoe7xMgGNxz5zEP3BlCUpRM7pSA/1zFf43JJ6aGx
4PnDo5sm4RWryQnyyYtmUG4sncyeJMacCz8ZfOkB6eZ0Fb76gHYp4cUP0PxTQal++H7TcxAhbcNG
IdGxR2bmuYZt9yOMmB25ccb9LNKOh8ZEiEa9LbHnEY9Xfh0t0RoeN+pDEE79ET0TL9qdXiFRxLLm
KVXOYATggUxcIha9P/4vIaeaTbLyDQH4GE50L4kSkFQntELjc26BOnDjwTbJVCrcF0z+jrusL5xN
X34emzvTRy9DmuelioLMYSX1CPxJaaVdZ/0HFW82foCUXMlY1YCUTmGw++5RJz/y/NwgZ8aYsvfR
1OiyY1rcj5Uyc2NqWDpgiPYmjdp1G8zCQx6rhC7QmZBG4qAqg/i7pgUGOuHHHQWOl8MQonTsW5LZ
uQgy8VITe34oPT66MByWuVpbUAzuBWj/bRPeyM67DN3rNlsq6jWOeZH45ODf1HvaPsZSl2viiKiw
56LbMT7KB7QayCMAHajpWZ/opKzal3vdHAQdmveAzCs+dugGrhST2YW2a1iGrKHiu4J8tRD6QNz9
OCygKTWmGR7BzvSU2Ud5KhsuJvPLNC0aBrFoveRCVz6F8H8X0JlMI+ggoDsi0wFps33iEekY1CPR
roqL3tjIzvX8wrv5FGrkLcR3YcWcQMEvGCpjU2ODioxLHhehrmnDrmZApKMKcIxHeNr1ZmgsYJmK
aeaHVhiouU6qkU+h8MlBw48bba8cN5oi4nVqrhpfafnFCcahLsHOOgwyL9NA10mpR0B3HqSSKjuy
YXb8bi7kEhG+bgmAqL89KlDzAhj917LXCEliuXmDuZakS+FCJ14MqgPzXbKZVepviLEIuZUl1DFy
lrM5bxJptbeiHV7SejPPJzmI/sWn/UC+SYyOrOilTvgXvWWZCqn4PliP5LM91zdPkY1Tr7WnJzGC
BzEkuGTDRVta9ljrI/9sGxv0T9OLGdADadJmJSI7umh+WQWnRQj8BVAKNzFFutrJDOgFT8ixpHKn
E5EsGB2wUZRIQl6vtCQHkZpAfQeppGAy+xvlMpeNez5rJhMUsBK0nIpOqHlbyKwNa3FzTAwQ2GXo
JxHaIyWzh/g54klO/3g/95yvGkd59USmgpSnNC3wzdjmxov+qVT2Hgj9kg65PXGjoCPfnRJZgr9a
7DNvfSrJ53Z+Vg6kYFXEJM9r6IOpxn0nZobGInqjx9ywRsRnapnutRvMtvPyU/Au/IOEgl/Qljle
MoJO6WQ/jZ3ra0O5Frd5i507y4uKWwoGEZtk2ikhAqT1cXQ+ZBmxtUzxwSPi3SzzQ7LyvA0v+K+5
HfxOpJTjA1Z+zE39YapjISQ1xiQCR65PZ6VsjgXLNujgC3f8WmqAFMsUeDJR5qbUN2hzZ4gn8ZfT
9Pkhqclk0ASPYWjc5BdBSMiwWEl2TmF7ezzjAR+xO6fZqFH5jejBzkooO0eKYJ+qvZ8y9PBd0G7K
sGeG2+N0ThEqskiYRnF9MtAdhC8sh85Bd0iTzoR2aDbrclj46epCIPJI0Bj5WCS3ICScXV1c5i0D
7ptR9nanof1ZKYlqA1T7Zqhf90m3eZMHjO2La0WNg0kQnlRaCMzU5xmEQt/9uxEXdyPfYMFkKSSM
UUrabrAsEKnoAZy6kWxT1b/jDSKhm2CZlAc+DAtO1Pl5p1u8YUJHxEdse/tal0VvkTXztZ8RQZoB
kZe7xeUNHz0uBLpozF00Xybfe6fVpe8+sSuDGfPetZoJ1WO05WUCZaeNQOBdbnq5OTMGjBH16Uys
abve0r89M7g8tolbpDd9ml9pXts98K94ah3ohWBaCRMUo2u93343omLCuLL5lZFY8vXZPgVEPMCT
964k6NsuuDgsDUASOf7FeTEx5H0cqZh90fUjpIcPfqKFV7guwakkDF6d1ZBKCHd8N+oNpdnyYTE7
dGaPhFrHBdyBj9S1BTASulYVAGmolJROnNvljP6MtLLZ9q6JWRfPrzN6Nc4g2Ope7+ciFUq5nnNk
L/6kJaGnDmUZlD9M2F/W4ohTIKPMIyN3prcm4WJR7X0elLVy1Ji7emt2lPDbKXt07NKzUQYylCEw
5/9JRJg0PfmYm4E+2Z5xgkPQ+O9yQTRrH3UYx18SaX+lIn4LmHUNZn4+uEYW55/1J/+YPL6LIPYB
hkOlzqvGKrWZ5fWSy8muwqSFNgUWafhCOyKI7F7/YLO8QKIbfoS6Bf948uEl6EfDhQ95yWKRppOb
HAcO1fTnJ5jwC5C9KaPFueDPJAi0nWr8JJx8o8xeX+Lm5ehyFI4BDV7YiM7oBmD9aQC5BrKV25Qs
/ilFXB+5ZyOhxZ1imsej64d70tOUHHu078VeMSnePiUsnS01nS7fsgHADCBjV83WVosKO0AzpCwJ
i9uS9w6jMVKbiJO6SIXC2h3F8Epz3oSbt1iqNOXezGOiMaGTprS4dW0fYYwNSowgHEYxtVoRdtXf
UEJeFBEMku4b2s5w2zvzrVRIINPAuUdm3iQ3CL8PWZs6Y7iY24IURSddkhewDvIJNScbbqHD4fFn
vwvl7FKh9W7zru1jIa0dtGF++6zDt5EUZnZ/Gyid5STHekLUl1wZid7+zuAK36jBmVgh4O1sZf5Q
NGloOLfnBthsmVeDxiXkD8LnZ8S/mga/36WKmrQYjptoCuTuNHVGLSyHrUjOOwKwBzEQidp5D261
eeWHj3yxyc4kJEotZx8i5ANbSs/hk4Y4qG7m5koK1+sAaZ5kJnTFTQPUfv2AoayNhBtx1Y9lIc9L
S/3qzp4X8sis2/dPMowLfvMQL+9sMehMCq67MfizhLhaNL66bOhxvSDevut6rVo4uo4qntUhaihH
eGEvYz0vSVN9mNojslUzy1Lk7NQ5/LKiEoNNf2P/uFum3s2i4AJG9g8BoGWMm80SaIpMd4Ssg+Yr
SApNNjlrN/Ca9G3xk9YZmGI9JeUFWzcxoINJ2k68YxA9OsxMAl40857rD5+Gxs/pbyjMIyO60Cv+
XVd6ChI7VxzcSMeYOF5ZUVPl6+Bx+AF86r4zWh65u3KyQauZefmzrSzw+LKa+PNdBWuht6D/aQvS
C+JU1g6ZuHx/4fGAmYmUM8FaULIhSc1O+7MQzXkstuYikUI/3rhjOST9A7BJ8auCkMfD5yNcNn2q
oRW+UZx8n94BkPPXx+7geWft8hr77uXgquGyBWwFGguUYkbE5OLaV2bec/2i5rFoiUurQzebIrMt
bTdwPduDElMNa9gO5TSAEz+/9H6HoNtjqQ6FXY0/VNjTNIvMe2BJx7l0hQoADpECi23TIKm1yYSg
falQS5FfipSJJ6ZhysV0v840XEPhxe3rpDL8W88ZX0uRKVjjYcTN/9zVdCYi1r14px1G++jxwhGT
DDxfeZTYo3sJuI6j6kAdrJlEfV5nBz5f+9wn5+471Q7cAaAoJIuRU0AuFE7TlBfy0AhyjsePr2NN
OteFjO6mWGE108Fu6Mg0I+iNgcocGGHdC1kx+qT8Gg7lP4n1pp5rHBCMIRmj9K68lrqgV0po2hrE
p5+v5Uz6LQZIbJur2SiGr8mGyoYZVgAnPPWXZ8fJC+JC+p3s6rUFCw3cpOhgJDQay+mGxcrPbUMz
VvYx1XUxINu3tzDLQrPRhyco/dlsYoF6Ls3bez0XZ93oddq7LumWKVzY2HNVft7qW9G6SUsafew6
Rz6Qy6uz3gTjDFix02rumgomd67SdVESsZgYqNHa0+Qak2vx9l1PGp4F9itH3yiA4d0YALa6FQ0i
gAZs2m8qx3Nthskqxd9733Xuk8yZndsaE7lRRMT8XlpWeFQvrwNCj7jtkBtroeXJnQ1km1l9L5lo
gaWF/pnuyWMGQhqZsjJlPh2KFGkab04Jq7vFZ/yjshHMLT1Vyn0jGVjmeqpwVIf1ohO5O8pPnh5e
8wG0rm+oNXAGMB8JqYs5VHebzS9xu6xvk+PMTO9v3cxLi5judSwgjPUp9hoXTgVCBN9AMmEmPEn4
IiFTtQmcF1w3PvL7go4ZLtkNJ3DITaL5i2TlNJcTtP5SQjmwUFTJZhEjL5gw+DGYUcCOYvZG1hg9
7+gtIW3T84kNZ8a6xIr1vEiC0VZNjUOAdnkYQJvG32vW7KeXDltdRQ4i3nBism2B1yn531cAK4Ui
3DxHtc07S1ea6pvjRc+gmzMlBaZ7HkRkRObmvw2Jalxgqe7BZcSIm3rOChu6gioZ6Vi2pbVuxtR8
3PRjUJ10O1dxPhUko+0GJaYNkoB7lcgDbhBCpWvILSDff5c5YvbwvMbrPMdqDZovVRs59wYbU/Rz
uPkQmXsN4rY2LqZYcLZyfivvjloKtBTWMprEyhhlSIefVcxzNw4HOG1sHiup8ShNiqPuOav+Uvdy
7prphXOtfXoJfzggX9T/Ceh1TNMSlOLv5wCYXKaw4ikRJIWpQbyQFpwu81Y0wXvtdRT8fmN86Wdq
ThRTf5QA853jTptsIJKY7W9lZLv0cfrP5nVv6mhGaP3CTkzh7RAyLiLVkPvHSqO5U/USljmXDicq
8+uhrmQEaM25Z9orHk+bjR6nkH8/lYhbGyFz/eFJIpAG4J4JVMo0gIQHqGLIMp+WIpKhQXkNI2C8
HT4GH5qhRRFwj6yQDbcR4Xtrl0VHhM/vMK7a2DlgZzNR/7dwKHNTeByKMnNhEFiqe/ZHoBILa18d
Cxm/qHOKVSuLfPIkG8XY5nngBsyLIKExNhWR1mWTxlsgmCkz7WqxS8MqPzgV8Sr1KAq5viBQaj8E
Gd5sXCsyaI3wbvF16h8gyNtYdOJYO+/y4Igq1/RF0UTXdYcnLaiPDHwzB5ks5PkrZVIkaKFu3XL7
5lGhSQykjPtAHE6HQazRX5QYjTlF9PSadQtTJk2iUy99aD96y0QCjsFBwDg8o2xYwmFm9zztWKWD
ZWDTX3aJ5j7k/vZZXD95Dw/WAFuYUOSxXFeRgkvRPQKH+EMC5NV3hf/7SoVNtI2zeXSv0DdKV6VY
VKTI7LmVC/IWrk9Y+Fihe4tODsIid8G5L9ZrioV+gxSgOI/RAiPSHC7Lu5I4yuY/BYsuyUlbuWKR
SMOpGk0Hd1VTRl+Q8WUm35+lP0ajIeE4pjrrZsoIb2BqBLHQVMZWNfiVGBgqeDSCsHr9xbZ3L5wJ
uQOBSVuOfh5v/9Ap9r//9Rgjh4HbY4rDJD/ydynrvcU70A3HP0l8/H6oxd5Danl04NbDYNoOIFlo
DDjvKg9rBLDCtAlBFLkZiAbvHO2HbAAxDy34e6MZhcuEQo95i9vYdZv5bgWoTLzPC7bElKCGAAU0
MP4w99DLrSkeCuEXxI44fIBQoNVGI88D7TASpjDIgm57Xm+iD6NMr4oT+tf9B8odnwzrDMZZjc+X
fOsfx3Tz9o2+PjgRQc6y/giTLX0IH7Jbl+gnelqadV6gACsoYZhpNM+RmKEXcin6mFdYezTAW6Zj
VwKP8rzf84nU4rdpfp8i0vYfcyobX8Eofg6K9Yv2Sbbl53GdHlFb8XJmN3miQd+VHxET762cc1Kn
0m750iaIifP+wn0dNXNDDcP4a/p9U359u57SY2Uw+G5Vkvl3Sy+W4oUb8GNjgSKmXhUM3/GM6zCC
uvBSLrUAGPuC6HGD/69J7IBn6w2EVPvqWQzhIxSLtruOKQGkmNHQ2T1qpb9v27pvZJ9Cf8MguRkf
Eo4ct/fSP4vfWbv2nek9sf+dv0eCFVWN0SL8QP/kTHTpqMbRNwHL8t32RC+IRM93hQ/R7MCbDVzU
X0Dwyj6d8pjKZKD0IipWdutcVWgguUf+nh2usH1lNZWtDoOsbF72tqNVQkvT6BgteFB+9KXoqwm1
zXm7sS3nU4PbJLsHm2g73C86+ztSAnz8gKKcWYDEf0JHTD4VbbHWF8MbYkGvtqSgwwoJdlAQALOL
C72pdXoVPvF4Ep57zPib6NE3s53u1bFaI60vZ7SbaoMYFh2hLz0eDI1cgIs2Q8RmoThPc3Fb+W95
1SqWyxv0S6ea22FoZOZY3KWabYcWCG5ll1LgmXsXWqOG6+67Iw45GIr10Olwp3dt1xJTvKuBYhgQ
l0b/p9IeRGBd/F0KsMRFrQTC+gG8nloz3zWIFtSXnPYMjWAJXDqUZGxC33CH+FhdMFBqb36Ewctf
QRH0yTep7X87OtszY/2ih6P+rQScIA9/tmVx6vjuB+mND0mwCNmcy0bhw+V2SceFvPLTNAJa9wun
Ry+dhy01B0Vkd+TmrYKPAkPYwQwWzksOuMv7U/v75f1sa8T9Cb5yQMEZFvWkohnswbid80bwsOsH
fjTFJi30vjB0UnZb1xLkkl6K9RfCeRaayPTKl88LMklTdGHvmgaN3nMjUzhrTZI6dIlLbwISVQ4V
qvOwdCA0JsLWomvEPWctNAJAtRtLISuxryvlWu4/KjwwIM5hg1OOxo7K6T3PuzLvBlrNACK4b/Wo
CdloUooWpM58Pcz4eaYYWZ3KjAI8YVAItS3mPThapw1nZABD5apr2NdyYYR3cNae2Y4cyPY6iWHr
Yggn6XQS0f4AWKQ7q+S9vYtVxc3tqSuferoYDePnyFVXpOZ80dzSuUu9RFzVfm9tc+jAq30xCVib
ZSvozB0CgTLTOt9jxzMBZKv9tGX4CYHkEHKW7y0SCByuO1hJGDHPSIXNTJdfOLbH5tiKS/TtsE+E
wUDr7vMtWhYp+pAOTjT0xPuKboWun5cV7CL29IPQwNx8u2F3IWhKgEmJJqnNjjpnEoeLBKIMOTYT
BBHN3J43kzx4NNIiz7bzye822tFR6YGnhtKKgbYqqczQsicmDWuqASUqxx0eV+vBaeDdq8yNbD6z
9I/YAJZtnulFLj75ddmrEsPHUts5znffZl6uSv4A2znnGX8Qsohdu8D97MkOBG5653NiSgRxVGuD
0OsXjqy2cwertawaNP1z1EQP9hYvxlS4k+X7K1oHoPG+UtN8qgW0rod1FtwavzwinmFDjjXMwCwe
JnfCeqFHB50VpfnzZ54is0edFAqQZMZtCU930rpkpAtm9nlu367VeZtTfle1iZdClrUJ/N7PlFhk
ZcIUocuWCOEjve84Sb9yk6PYlRIZiRKAiDDbCZDjrJCfpC04lpcthE0euqtXcw/JCP1XgS3Z7DZp
rch1b3N8eFCndk8kcmwtZ1p1esUftg3/agCDSdaqlNReJAUNdBlu+YWfDtrqFjplAO9DglqZdYK0
nD+ewONEyRuBf4cveBq8lIU4M2QlYC+psnNtPUZJVw5//ZI6ZNHOQedQ90WMxpWYe2Y7bVrBNRhF
AIMRc4XS9tHjnZpfyEqSiUVTsF59w6AeRfVLdmd/ae5XsYhSispzV8pueYiEzdKswbOpSZMdybMU
Lbn9q7nAUAk2Ksxfnp7acYKNO2vXXTCPEneDUsjD3ik6fNkN/i5UDgoCxWnWYGArfx3Lu2X3rV4I
GZsAhyPA+n57pQ/I0mF97vbhsVnl6VUYdqR7DUttXTUb33ECmKaZNeco2ylSOy4Mv4w7FU/aV7v2
hF+m+nV/ot7iFc+dRMdYo5LbT6dz/VRxQRjOh7DxmA9v0JdVzFG5h4wkkS1iPlvTVqA2LP3HO5Y/
NPojUk9yJ9yMUTCH8pHIv6XDnEn95uIGfooVZg3E3n8z8C7eDK2ZFXdHScf5x0RYAb4uRnMnlzpr
is+s5EaIhCTSWpQH7vY8x83i9BTiN6ky/tmRcs+JyFplJmq036c/9vqwX2RVGCZYF29m6Qb66Qk+
Zzyy3PJjvGbw+UJylSoC4gxMhI+uuGA4kJMF3HAr9fDGDEUUMF/wFaXyjLxfeFPELf6W1kbO0tE/
AfVm4lql22X3WyzZJRjfPzSmQDeEcQgBqDt3Iy+0UGaEqatnWmdIvmMWyzKhW8OjiXGWqrzKsnlk
ilOBqteWf394ZvmOLM0juhqo0Jko/Q663W5odP9utPTFfoYcvoAUsxVO5zbRauqf72uDNO2PuYQH
GrxKUa3v9Lat1ciVe0EuovnU2ltNLRe5lp6aaHF3Rqmetsmbarztel8NJCaL+8Ue40X46SdrGVGp
Wh7VjH7gt/cId3q9WMePNQGLd2PNqaXJA5eC9tjU6oylQc5HjVP6IfrAkFKesSJx6H04Wpknk6/R
HOfTIUUSQmixJ47muGlwMab3lfRak1dzv06/RqgC/oZBcLKprRN+0oIc4irCugE1sVUVW5CsaeRl
132V9Tspb1rCdBXPaQMHJmtkPVdZupgvObZvQDAMoELJBXmgOW9HJrCDCH7CAM4FvnaD84t4czm3
I6zUfSjaK+gpFaWEPCRLIaArWvim+CfBQcLwoD0W9/QsbhSZkwh8JRhr0HyzmyNf6Z5s45Gj3fB9
cNm9iEklFEZbOOLQUFhELVg2DY+6xoIrRqSysmag3k07qrUHDNxq1MYP9d2Web10GDP2caplpLlI
pY+Xn7gKQs6e2sqOjjW1UQuLd1CqzqzCCG+Rfq5bl63Q+QLY04zLN4qbQ4tXbc20DbICFUxx/H+S
ilCJui6QPFy4I5jncvlUD4d96y95/FYnGKZkbVaSsWQJEfeb2s1R7S1gHORyNjI8TTXAGZSr99tx
EpVqglOAg5AROrjKL6X2TST9vTYdxBhjvWGXi1P5JWNIL+KUjtHMp5TpCWZ/i/gcXUDIja5n7trx
qln+kELRSkMSWEc15z+KbG3YAIlSRYGVghvhszB/9DUzn89PDP6lo3v41Vf5SNasAwy6wwUSPc9J
uHfZvWQYOULiLFdldnMMu9qtGD2oZzLyUtjCxIc185jR5RTnhpS2TaPOFy9hhTA4PWT2S5+NCeJZ
rvf2wREuk6Ke4kMXExTfPL8dePWq8DVdj21Mo14N8eAFEKrTh7etIvrHkCuNWMwzzHZzlFWVVbj9
Oj5l5UJgxmE1l8NgP2xXzupSzi36oAX8fWcQPeEO2AEvSbhczur8Igbmplb7w1FCIECJNYBIb8Zn
/7POKblOXvPaBT0LZbzrORXwCciyX9ag9eCq4hnhjA6KecikfpkoR8cQVYQxTXyTWGPR2uWRMOgX
ZvhjsvS89nVyuJuUSMWa8rAgiuSbp3vXtFYb8Sl3hNJeoQ4w8cqSypPT1poA+oeVoqA8coppndbX
+Gclqiv1w7pkbjHH/ytcERpR5ocwjTZukH74LseEsk6Kd1CtLPE+jJOeFoxPVbYdbjFmWi6mnv6i
R/dIYd+FX+e7rSlnJDDewQwBCVPnpicUxU1WfBQd+1JSYqWLLTGJr/FSu6ZC0BThIae5CdylNmUl
f4AvcYxtJhMjJaxIUNyembplgS1V6W65JHcghcxb0onJE76qaA2Px4lcscE+60LtxMHQav4VDJ8o
P/Ztw7R/MAF12E5eFno5uFtLjzpfRKcGVzGxh3h1Y7EhRcDYZfYhR3DOEdo5+AXTrfv+8kdDaqMW
sY4CVm2dSDpEE+1BCWnSFW3CwCajQM/5DqbZNwrOzIsC2ghHuu41Y2aWJGJk6VTbViCgd9flahWs
RXnK5dw5MWkIqO45c91fW6ZogwkzOOOtLMI3bEAJI5VxbKsxbSH+JeWXWzgNh39mUTXYFKH3xmdY
HLDkpV8+Qx6Ex+rK2PqcabULIDZ9wqpvvUIwDS2daREtjmKvsogQrjANT52r075lYVQtbcnDpehA
rqQA3gM8Gt86Vma2NQ5Zj2BFtz11LXhMVYZQ55diCb51B6422bTBqGzkz5RiSNqlBbZ14ktd9rub
CwjHXk9LaArYSWzuakO+3sZiE3cd1ZVg/vZStwSthIfn36Kr5hkNAGhikBL/wm8DUwgZe/R61crU
qTPN1T2kfFCEdm6dlezthWxQeFNuCrIaXb9Ze4qK3jqY3Et121V+CuwoPBWRM4JSw8cxn5ezCccW
jdoABXvyBRbDz3XfmI627BdR5O1gJ/ZEAPfRIc2BhVDp34O049lW2A2M2f5HmjVlgNc8q8NE8+Et
EnsI4zR3xBrX7yuz/Pt6uokcycylKuh+BesLqePUQRJijn26H1o0ZQ14AHsTGfZskMHv0Oo4XNQZ
/7P12SmC+QCcD/qtWJ4y4aZFH+pZ+iGnLrBF97fherFSdxGfU0muL+xrFV8yL3qlptfCZJXdeQTo
RAxMWjdwot/vzpn9Vb0vGOIe28YAsq+clq3yFTgrDHH8DCwGu6EEh45Ajq+nqciNcb9SNQD+oVc2
4Q5PLbmPtn21dGaOXIUSNiM7ZjAKsSiCmixrMZD0ZuDyXtISBVbekKuLWFhNTsUKn9opM9u6OTKM
N/GnKShOdB5FMxFyN5Oa0v8Xs75Vzi1pazbdUw2Gcd6/s5wFAJWzYxRNosstV3qXYlfv1gm3T8g0
61g4lLtYkY1aoM2AK7T6husf8xAB4orx6bn9d6Tals910HVuLUXl9xnIoFrdxce3wVsnRArzKERZ
Z23d12adbeSYurQN7cubZKbTWYPCRBkGUOC0CzEM3fTCOyw/uW/UF8YOM0b3pqcry0CHw98K9MEc
5aHgL5m/geaI2plx6gewiUOqRp5XMgXobRxECFLZbPosHc6Q/CVri0rtLBKFTj1J2ExBMvk73JHS
zPmenh5yrIz+ZCYAWRdzkUsgffO18aq7JRzqJsuGZOtS9khxrtObADE6iXBEo7yEvk8Q09CDpcq7
4XP+KlxZpdKnChgYlrBQ5gIayEm4FmOLsNbAgpASmBEHuz6UqAwZzQOeEPuqhQC2/ctnJiaG5xee
AWUsDGecR4kOsQEYP2RzbNaOZESMXPN/QGwe2uCwTh5U3RVO6ALclLQGnwNPOV1DzdXgVLJTljDq
eO4ysh/2XhIF0zHllbCMafVz1aAFN3r8Az80ihe5cJpvCX0g2d1sgmDlIU28cyjwKiSeP9z8P//6
b28vEkhlccFtiBBLyh6jjEJ6RqqLxucI1ib2A6H21trzwaV40yvoocNXp2UY2hH26b+xQKyusEmZ
JVSYWC/4TswNGRO+mNpFGiD1plLZgwFaDAlp3nMn+rewhSDj4WdjgayQpAsJnuG7WFRFHKpEbYuY
zQpTN7WrAt1oigggk1oqAOAvLwb5Wg6xCG0xbDsm3pCKPM9ng8qGjlT73uE4eEdSesyFiE/7q0l4
OYE5uCoqFkTL/MsL0kdM01EukZjwkoBe6+6KtFKp7bhkBhqmSm4thReGe5BIVB6lVMpRI4v0ctzC
RBI0ALOOZZG79wb6j6gtYrXNVZuFEin6YABzZWF4YCPeCdxtf18c5t4wN5lGhFHh6XyZ1SD/o4E5
Vgwgno+T/AzQrQo94vK7lh4gkc8ZYX8VBBY7eSXloOsMlkG9cDHwZ6Twa37eBQLDOuoUUI2ZiqX4
QdHbZp85/UowSL0TWo96WqAvaPXvEqpQwvTjEuTOdlKUAykkIAdRAAlYTadVcpK3/xe7YMHCt2L5
3LMSgZsLO+v8T2ffv0yu0tAXRP7e/tKEOuoOGU5rk+/CrXK9KbmfttOiiHLmXkRexIoWVDPCFlkz
w5EZV07Ip+vQsYOHYYtLywwHDyflhryFpsjCmUjJzqxXwyCsT/A90OlCUu8KEPkCqwU1uZ268q35
StRmjnU05lR41LJQav7vs9MweymLEdzYRCzmqzjMjxjxSPqcLo6CE/WY/OsX8c+QWKxg8suTycbR
pw6Q9R2qbCbIp3+TrdtEjug5bl8/lMqTq2lZN/ZD4AD1HbHmMldGQ7B5F6Q38h2H0DfAzNwLBHPl
GOd6HL6sKdbqLl7LXxD4cOBq24z2BhVOdYqv3Jc3Q9JCbLmFOxaP8X4EdsVrKEYzKVaA2QOR/a5c
Zfmop9fm1Z5Tu0Yca722w4AHBuyl3bxgpwHlNjRuIJtT8PqGAR7xRrrc9wijxl4Ln5/LQLke5pgl
MgaroutBPxl2hqr0dWdQorNp7A2K7L60e2E+JESPmmzYLyMR9f0EBxPCtalZTK1eQt+dd4xfMR0W
FItlHzKh7foD3Q0P0+WnsZ9H62EYchxF0m2Y6LhTPFX3x+0Hau7yPgqyXaITrUUUQzuTyd0Lv+I2
XmlmsyJOMQEKlukboZeE9mZcJNYpNvZYP1AuifCHmzp4VL8LGJT8jZq3blB3cyagFqEN/z4ytZsm
YGrS2C2sjRhHpHck03At8QUnt0OEG8gLLaBHnmFoKxljNl/0twlzT9aRRrN4Y0My9DpTVrJ19Ejt
lFeZYhP1dMmrDV9qLc+Q1cg3h+vOmzYalXLxcj3fU0+zyFdtt+rwXG+hsfrTlxit/AvU510lWtej
ISplh70Uizs+7Atzdi6aeQjBF3Rj3vjkqIya54cxpa0NqIwotwXUb2RzRlFeJDg8SLlF7vbfnUgy
XtMWBH0yFLJvk5m2hYL4k7Dl8Dniop5ElJodz0Xy3pVY7VMXR+pyJkcnEBoyJP/q9UDM4XYejEiD
EHtoPDBfKBOH61zOlX9tu4CnDMULWWzVZZmtCMrZeQ0RoEEZGnsjF4AsNHDfcZPo/zIkfcmHWfPW
2R1c1d/a0bYzJVsFeqkgW6dn5zPgkowH8Yfo81z4Ul71v8LBnKSaU2fWJVCW9JwbSH6IyeSU73LW
ZTgdCH91z1QxI/nu0zRAvVnhYlXLN3lsPytLBWw1tnLDgb+asyVi1QAT8BFDti9jxYnWNXVX4fHy
DeJpErTCi0ZWOcbURy4aWF95/i32LVmpQrG65B3tkWRKmHzTP+c01koLw1DCe0JUEN5W8RaRCY7W
t2nXOImu1mRUy+xCxVUQpqhcERl8GYAM2k3jz7U8p5/0weQY9x2B7VEsl1r8vHmZ9FiovxTEQuid
ga9asgBc+I0Jp6Na4nEj3AHFI41DyKwHTQCpAkSkSwXL3VdMlWe2PphqGOE9XTnzR0mwcLwdOnCu
x1E0Jb8RQsVHutK35/KDCBnkFsbEn7jeYH5d3sT7A/JaGENLEinD0Q/U/LYaCHqaSc2/WS7eJ966
so1P8COs3oFOcfa0/bQYQUDqflRD0s7+IOoV2e7V5fuelqRg7Uab6nerNK9NwGwMUMhGimcEu9DS
0D1ppDP3P3pQQtWMA2Kb4I9dugIu04fEdhqscPWeO2/pwFZlIw6tKzKVo0yYi4hhTtogLTpT56SA
CmQw4TV6mZOAqLjpq+X43KjQXYDfjP/ae/Mlv11jUzINGihe6NTKxSpErASvlC3qvn30EQ1xNasL
FGBBaHXC8SrXd2F32tFd4vEU3sUGbFAyYAbyCnxuhSg0ZyOdqQpwJZE0y9XABNlKO7JwRDjJ6vk9
N25N6oIbCpRqKKn81+WDwuVL9GOsHqmAAUHaZozyfjb3cxMPtUACifdzk9hfKdTPIf0e+SSDHuFK
PfHAqeev87Ik89vZBkwGxDz7bDNet4sRxSHXRJnNVbfPYL4vRbq8s9Vw6zl+FaoXLgm1sxwjNYGj
wOU9zvm9Po82w4hTkYBQq1kzlSih5zjXfHR299PMAjXb1ZIGsx3TG0e55bynwHL/9KtcQ+b6HRrT
XeJsUtBairL0Z5lvtWXD3nJJ5u4nORCz7lkiXle5vweOjvsoJ7Mo7g6JQ5wTcnxjbXECdyfpRM7u
TKV1AQPuea0HaYAljPCX5F3lWawVZbDb9obXTa4J18xkKyyeHwoB3F2rUoylUu+usK/uQxGH4+js
chont5ILqyHI4RtGSjKblHJ+zMjaYzfmxb5soPi4dj9MGpfSvx6nUwk7QtmMjC52gJ1Q86buyqTv
Sp7HEd23+QJozq05BZURPtG4D0kcuhtCWkEzuVBn9wGiilRI0sRM1G3nP7Sc4/Gm52Qvycpu/gtu
Kz77pe+WG0/OC0frWX2AH9YSch/y5hpj3QNsSwrIghSCxRBTv6HPy+OMF8ucJ8Wkmf3W/qQ2z1OF
J3/paoojcBslSs4YFYLWny0E75yYTxNFJw9CgxMtKCYXPrR6lYbnNjXIdWQXrk7t+FmN7MU/nHvt
A6L8VURSzd0MpnkqbXdVFDgdjRVOOWFHJFH+MQSEQKKulgE6LO2WjeeoAcSWgbIx9P2CYoMHT7QG
juIs+ZS7pd+ok17kwKtDqMbP7M0L1vyzpSGAAeE0mjZDHZz7vgKzBzibf3W0TmtBkqfqD5jfgkDz
sn6nNk3Io40kj7oMlTdbvKHUjxdTAp5rsJ24Y9xEUsHZhm3Amx0VSY2+7Ib4UK8fOHMloNV2Ho6Q
D/IQqERU8+xudnHswel/m0iZhvdERtQxu+3ESjJRdbl7XkGh6OtrcL0xJi7GG0XYzXlbrxRNdlVm
6yuNL9QUwrcUbTOCQawwcIGCeERME8A7hYPiaPxmShSmezpD16a/3CuzuNJQJ+JyH8EV4oBiuap8
wft3TUw3FkdBO/YJr0O1zOd5jx88e7joVkw3T4hwNtZCtqmeOZwrUpirwVbmVepHMdw7tr+qrxav
8e882cP3AptnDXwDDTmXFLmXY4+lZ7KGGw2YnCeB8lA2Z2x7cl8worjidYWMMlB474LkSKGj5ogV
9sAT1JoQjKA0NQh/TngSPhobuuAh7daOighaXwYMQxX87z4ykKQd6dzwE/RT6wrqBXWshiSophHF
/T3qvDg+KQMf850IVYNoOQVUsNUhO7yhURiJke59mkZ4ogvVgLcHDb6t8XizhGw5Qln2ZvqzybRb
53JQVcrv4Vys10wgRLYlaWJy/BC4w08W3hGfZm5TLt+rgIqMi4hTzFgey5bc5tn3Q4OPgF0XYWoU
KTcf69E+tHKpzWPQJEjwCrbQ/tDM/4IsYLuSv1F1kXvusQqaY/slHX3LEvxcgLvLq2CDffrOb111
hWw28Gegx+k3OduvyUGY+VQuTZj0w21d4ES1Kxi1ju5JW5ky/OTN75Y0I5YNsXLe6/e8rVE9xNEO
hu1C7zelG0aRCMyYlP03m7fq3im8xSuYP/ITj4YrlCL/Zjsd7BjntuW4/e/AiGw8BnXKyQelsX37
TFl3E9/hqzF6iJ8zDuOo6hwSNk9NDP7WCocCdcD/ljsty+XyvJVXVytpBkVICxpgOJbt+zAKYfss
CXCZscSEGc826W2aAG2AxychyOt7Rv+ieM4prHkx+oFQkD7zo5aaIB4nlPGEXsZ67Sr/kR2gpFZH
Mw2Sldz58lg/kOJKPmLl27L0/VxUYHkTQt6xEFfs4oWyipWHbcjxlnNI3klISqYGAzi8apxRYv6N
OXPlh39FE+VwFV2QxvCgZcVFtcOtF/57SjK6tjudEpFWtPGhckDTlZIbechK4kS26Hm5cj6vLeeZ
V23VBbx3SuNuTT9YV8FR01uDp3k1bnPbsiqKtSt0/GRQ5NpRZ92kBgyccwbXRyz+bMo2a1ASgwuf
fMAARybJOep9jL/3n+EhUMQAqI9HZJj3l9edhk3kgwA58TavFhxq3cy9Y3Y8kRw2y8WauHK/MeRh
/pKqYXwtX6JQGYWYjvbKTurh6A8taWKFKrIx+CZBWwlRV1qmLsa/xiITF/kFHSm/+4Tb8PKDWQml
+v2oxnTx832TW/h6XWHxyWrjiPEZ6uaIeD7HyF9Lk9beYMymT9WamHPpdawtQVXQmcjk1Jp+xorY
EjCLp5VZ2PEXATpGxQZoJbbl78rDykHAa9qxz3Qz29CgNNs8aamFYm+Q4xIXWT3qTex1Fc01vSya
jzgPQSeYPz/ZG0nAUlY8V8hx6uCnt/xHEDeoyuCrW3OQPgo33k+ABZMQPyrDdoPGRcFy5E/cKGya
MkICdWbVeoTS5848OAhclmUhHUQ2749Wncp/W9lcFh5sEpPWIa0J0eDBQSVDFXTkntO5EPNI7cF0
wAV1JYGIKOid2YGrppvrEG2dn+b3vjA+GPVdssMHVemVB48C+TiqKsaw0QluYkbwhl+CwbAzg2dY
pBOL5K/GBiBuN63VHTqG5NWl4a5Ec02Z+W5Yf3e36NTf9G1woltEZBFH8kFVVQ1rgEDl+c/Kcjim
k39fOD/YNfGRBqFsIEpUeLAEBNVpEJstqc0LUklfl7zbksiNwvhhHsdQyFJBbJP8cW9QSWLJ6IP9
vsrukus1a7/2PWzrIZ/nxoMa3OkPwC0IqMe0hO9o1KcCoO9zTagaLPwmKEcGOwgv38yXKMBVe9Nd
6XILfCmOWH7nkV4V3d89JIho4AWskrygDTKJCwqurOjjvB8GUAF4YOPduu/HIbglEypoVOFs+ZPe
iom3mhpQ9of+aMZfgLap6z2/7mrW9j35rwjwIii1GxgX6yM97IWLrazV4noPYuUXVhNVLlouAFAJ
nTr9BM90TnlfYFZp6i5XBWBvXpo6KWsMPDhY41wIjxg7THoql+unDlXigNnZLKZ2/K/UaNEDU3bI
9iF95oHWsfduXaS4YPuGNpC2cxfctBXIn80bQidHIUzeEGBWa0UtpNzd4CgPJnsQD9Cq4TsVHLaF
Qv8ZKPqVCR/HdSNNU3AOrlTmfvh0RBEPPN3jyDPF2BuYYpfcfZmEfrxn9ELiiXfP0sm9jGTgEIz9
AF5yfQvPiuY7v4kIHJ56ZW3aqc26mkpyvDf/DchE7at14c6NxCoKw8haAkT7LjFBUgvWqj4CBqbr
At7MzPNVHpoYjc+S7ehuwuW0jPc0Rk7AvN59bKOzz6DdtcujQpVV4ZePka57bIDdqJejDUS+kB86
G7mPSKA6jreMEUIfJnXuNdxuvqoNzpSiP5VsKXwxG0AI+MEofr8CZ2Zf0YSTwTgoLVPCMcDmhT4U
JnmJUe3VN06O/TzluA/tyuYM883SsN0MArC5EnwhMhbf1CsM97XlHFyg1FGpyRt1jBKVdTmT/Ihw
wGWGyxfr2+VTW5+BqE/Ws553yd839eaGOi6VlN+dz1pfYf+cucySSeL8wAnT+HyaULwWmiwhc9nr
igygAHO+ZhggB6f1zJkErUNUzxKyplPk6TwmW0uGjifIJdRnCEaHuB8HTCy4X7NQ/9cXe5yQPN4o
IEDJAMeRs6F9ZiXOttWXLnWGvLjUBHyiOV9V7q8ePbw0/45z0/cfOrdjgAgW+RafeQ19L+HIaOlB
Q3+ONBvxF1YkyLj7eg+txhMG/wU3+drHspDqnLNRZOxr0lHjrxSDGUalekRWMUjsyEAeUyqND4DH
mlZkX1IHzpy7CKne0JLab1d3CRPUJW00VRuWUNATLVu4UDjueSoTp6Ztt1oAuxR5A0hHPZiO1MYD
FWW6kdt08fzc9T4niXo7jS8CxhRvTPhSVwG8sz4N/9Tl7vm4TM+pMtz9ZtPgRMWzb9THGSBAcFg+
+iyWxK1vAeY7kmdd1X9wGVTcwaac6OZOgusqkGBcsTVqhm9JYByM2ZD9mHy6NGJS2+aQkGDvsrh5
qhyWawtn5/zbt/N0SYbf9w9+AQZDgasrN00T2Se3nanfRwFWBUOmMG3QNF/Mi/jIAE72vC1LKnsj
Bzf47z3PgVYB6M/Wg7HLethKA4JMUXKmKjnAiYCj4+0XFCO8APYM2SIHkVrXI9pkArMxayklmE+D
qGF7qNhkNZyoOObzAw1o62ydXgLcD1hS5JVDEN2m01Pz170feWpF6xxsnCSjXQNlX9vBuLt66RxC
xunp+jeyUzpr6RIwRtdxnZTHfrhFL0LbzX2Tf7Ub/82zYd+QckfBLcmfV4ytVuHcYOLoKdCmacXk
kuH+zw/nNSsCAvj7FfR+JoiPAiHf+6I2h70Tr7+TN7bxUY1acDSHDQid9bmOo4fRPlWxkYGL9NR6
+EN08zvxLv+WXZ2+qXPxRkjViILqRaUMkwbcRYaUzqeBAIHK44IrDBk77cNdPAtEJLq2CbWcL1ug
2bTlkkNdYcEBIE71a9WDIJTyOVpSIB8y+HaDfE3PIn8PcsL/9J91nVwL+ysrpfZzWaOVApmcNzD7
GgLwf/aM8cMb2VnTle677iPsWfnXZZU8FNzsLObdLAUpqZXWlfmYyi8k7jJSOwE2OMjJWYryXle1
8/6PSBhk1xWK2Im3KufHAHFG2jIUJUVoOPwlEkGvjkNRVizn48BxM/EyjhxYb+mBZcgEK3HWn3K4
aXhJwRGYbpYx9bVmXZsqinFKm8yKbjrPjmrenCiKktvOrRAoWMu3zA/jYppd+nEaflfUYCivbmSB
pXCbLF+mma4uwzBYBOM47hajVCKkPhyJb1ZN1wqp1RRbgv13mdvrmcH6C3jV14NCiWuCzpDP2BHY
eC25Pqw0sT1typsIXKzAZn/ZubIqiY22hOcOAMPPCzZoPgbEgdjDilI1hW5e4ZcjYQm1W83u6T4V
YYORpouNcHSIsmnvAJb7SJ7Xbos1yYrFCp8RgVfF8rIqWopBPdkzJCc1HRBDCBFWMegkFjWWWrfJ
HkSFOHfkYBRJ/XnNBSY4ToEUmTsb9k8BVAdrAXOswGTVpEG76mVsdPQJ4h9zahTEZe2IBbidsayK
vw7zwyaukiGRZhSM8XoKDRXyR72zWnSZvIaIpY7zLRE1wrMmv6w4yS1tceE3m8Yq2JtrEuc+I8Zn
RmKNmadFz0s6srN9oPX2x3sUAMkallG0CAdBF02QMwn/CpoYa0lBLhjo6WNlhqAdUSKpdIxm0wqM
074YGbTt9sGljDbYiCYZRbKWf71CMOLx/JwE37WvUJ6S0hGY07QXkOyvqUS/5TlotQvj7BhXYt87
/NJaS2MGyuDji4TL7jBKwCV5BH5LVqRr9xG5vtoMtissJ4G3u4RU/nXFDJdSf0ghX1gWYA8dX27L
E4WJF1ue81TMQZj9M1nbix7Egkgwnt8nTm63NZ/UpNSLkcvSi+k697vA9C7yD8aU4LyLNxFWwXyL
B54OwzcRZzpsTAN4ONKApF7W9dUym3FzO5K0hKqEeV4KHZra9UlnxSk7JRUZ+biKX02XvuPBJsc3
wgCrqljjBSP8wIPi0cjhDjpzLFf2Qhqo0FVfy/H8jMT544ppH/83D8NCqRBknfG/tokzS9Us9kwB
TEa5lT6vpCojPP+Ww6uyq0wnPr/jQIRg6exkX9xUxMr4GEe1MCXx0qXJdaj2bdMrxGWGU8xHusAD
45chvThczCUkvhr38Lhq89teRXK86qblKv7rFJ9GAVe0NHfodz7O0+oGp3ZWULPMAQ+eqy7R9e/y
DJiFWNy3VOZW2QVs0VQMVreRmzNrJYk9vf7fRGZBntruXs0LArEs4/oC1rfyz/FzdClf0PR/XcDa
VBBHIsUXbl25aqvS++XmKDOOSikWjdkGpe4cd9L0YwY2GkFzB2n8BJ7s+gv9Sr2aV/B8z4EbjM5q
0cdEh09vgWoXS/873/rHD9hB9DqZzn0BCOOf+N8npaAJabVln806RYXBUw46hXWkcrduGvT/E/2S
N4gP05kUwEPyoILWUWVLzIBSaLK9wR/wsCMiE4JChMD2v/3TnNzpcOd/ft979dncTpVm9Fvof25V
2KARJbwdD59xcO4SZuPRx6/WmfCV4GurBpq+kyYcglYenLNro1v89zG3MTJeRjRgv6uWmbrZKntw
dRB5JO6YxYSYXZxancdWNUchF7BgFCmwkPvcWbU8wsyZFfvd0qxJTR8XLQ5ZbFiLaw14vxpAt0Kn
2A3AbmKHaydWVAAZe28PKjk0K0bXe0ySLuspnCMPo6lLdmPKPNmI3nOiNbrUYFcxdzm27g/pAdJG
R7xrEb2hVC1+ODuna0dyc1IbKXKXNdqkIbI/BxUt2xhlUNRKs/0kCyKQKEZm/1K9ARSsu4Tc51v+
Vov4V4wSsRTWHzgMyPILp/MgVRj4wQBD+zG2nZ64HcYJdNqr0cULWvnDXmNoBNNP1Y52NHP9Gezb
yA0cSOXXXiQeSZBPu2SKdR6GEsokP0OWF8KbCayimxd2yhruZL2H5udj3fuv+riRVc57ZFVMAf+W
Vcxljee9QDF8SC4NHGUY9YG5N4oZo47/c6CinNNGfz7V8N52j9m3JzPGpqMEJ/SCaxTpO9x8r9f8
hPV93gOG/Nvm5h9KytlkfBfGO7MyAolkQWESfY8f5UlrZzWTU5W6YMV/JFj24FFGrjb6zXgSrq48
7HcWQV12+wpYJdHCe/wmWSl4w+23hHsC6NqYyBLjpXolbxHV9HzaK3+eiyeCNXH1d4QdRmMtgezZ
seya4LT1tXddbj6lf6wRiBJ2Fk3sa0bQe/1m8Gf8IVVQZYndAJA/GDwYd09i/1pZGJ6s1lrXsuYM
8EgbjPek8O0AqUi2KD5UKVc7bJKK/rcGHTW+3GdAhiFg1FIwNW/elD4DMk5fZLkK8akIWVNzh58u
4joymC8SCiDvyz2HBrJJeVrXSXo9MagRqkpoX1WBl8hW6Xj78t7UQC4TU7mf9qcMPCrxJ4QdWAZR
R4oNZ2sAWCycpuZgClAuaK2wFjk4ovbMPxpE/ho+6M2xu9CYD/ma3CCl97YL6nOZVaqgHKrp7zh5
RTVgl5uOe1uD4id7eD8XEkIong6hnqBR5KWOO8Cj3u7EXQudZFuLD30LBTyKkUH8E/7irUxwdBWy
NgeMWHBa7AVkjESr/H5KWZLFsMsxm2mGZNQpaQJAKNk24Eiko8w6GaCDgtGCe/dT2RxmqqZr1YrS
6nc9wBdkzerVRujMAZWDtSk9b6aGk2JxiQ9HowNEjAOlE845nLQPlcZHYRfgBK4W5N3zfHzhBdom
ob5WIgSpBUo17o7Bggr8aPRNgOYzf1EGc81729upAcizcdt/mvJobW4P55Em0GWRah3UpPJB0pDu
3KNBFIh9YzH0zfttt/a0zqoDbQRsaLw6mF/Q0oNV87NswVXZJnsT9CPtZuY8muU+W56xW0MJhZ+0
Iu3u7vWWzwJlKsoHhje4uQAG15k2LjDuMyuNjda/FzBv3EVLhJOLyeEngnFrvYZqUxfSJs49fq/f
4BfXz4mb1DUBSRTVll9j4jyXFm/dSepYsEsHmeMZv/C2es98vXrnykckiy7MnYi7qNlSSxHWVsKY
E8v1+6348JAqkHopfpNiqEgetKts6IWpNyfnfNKcWRwBidKxmHAM1EhTP6FXfKJR5aImCcW4GTj0
7gaQYsodt43xSSPxy9fqQOqLONJ7PgvftnshDR6VwaTgHw+dn9Im8+is49YfooOaa0wq//co+Wpn
1sFlHtr4dhOjqD6ZRoTlc0Xm2TpFJOOnPmxwUjnR1D15FXKw48zWWCiSGMsZ/pPHnVHNhhuvtLl1
1ItpQmiY/xL0p+rkSeO6cK8ocA/uqFlFr55Ml/XZVEl5yKF1XUyHic18k6PjUEJ+bv30Fiqarimm
K4NR7IGzs5PlZx/HboVqQWLNwksiRbqsTroemjEk4Y3xvV8x4M/YYuSedlpxStCUQF984CxOznSM
F84LPDgXZDcaYhiExNVjYktVVUKvMn0JiuPfNPW6p9OmisfdMhwoDtv7VvcTKmCT36EGwOkD+vbw
nndM+PvU9Z1ntu3kXo9bzuRpNovfwRkDZqy5s+lUHsTp18PU/lIOKh2nYAB2h85qTaUdlQl2Rs0x
sqHJH+w4lPfGjiuojNhtH5koJHaY2hF89nopmbZ3vRiFgovQqHFTAZGUynqdOhJ5OGrpzPkjpwsn
VwYaLY/xzwXoFPb130JbrBAa9eRhVVIoY+ZT0VpYL5UPjfdlt8eAcYwYMgfN1AJGekgs3wboUGKS
TOAujxUig7Chtc//wxali0MAWlr4RN7jnKlnob0GqZnll8pKebyzGyQgiXG5Kqy+jrAMd5n0W106
sGjegIBURRu6O5DyfJKIViElTtavp+b/sho/8X62R4rtBAzsQrxqsF8QRGoY0Rl+iwrICuCMgf3n
Zw9EQhesCm63c5uHsciyiJW3gNH6PSSf9t8MwxpIRbtIR8Du+SERU696bpwAKj9Ss5kbZQHGuUfF
fSiRwRZ/Wf3k/Lz1L5bg1/FAdu8W9jgm4mv/Qta/CtPnwTp775tMrv5rVCLG+n13KKB6kqiDxMFH
6nhIMEWCmeIhxQP2r+UN8GinVaBdiRuM0yFXtNBR+ZP0+hWdvc1Gh9Zgp11zjrz/CzaYjmkj+7ke
0Mvkd9/mjqu0DCEcC/t79wbSJyLIYoGACnhxPfsENwT89QCCnAtW8/PHf/fzrywDtRrhDFNbmBka
Fc4Doeja0xg01CHnGWD1vXGpDTPDicWV37yhr3fi3qmoiH3RFAc8dpSYQHh+PS2kZsef705/3N4/
MVC8Tep0tb+9QdxSkpp1jg1hNjWXbMtSWIVY/VbEOGBd4CI9uutdDjrapzPHogOekr3ltqB1EX4u
NuJps6TkQgVmB6DspKd7rgAzt5AxAfxfEMHE38cnDWP9w7XL1BlM65uDXg8Nr3vjbvghInQl/32q
+xuQza7YTDGsXcsxgrABJKJtrctnvNoNWEXdjF7AXeO585NLfJpTnxk37GCXVyB2Ppmx7sDF8l6m
lLYOGlJRQu+Xu4T7LlW6ruMUTDoLNDU8k75z+xHi/PM1dm0rfmvToY3UgNpmSBzRH27rdL3YXAjE
lyxv9DikFf9X/dlKVrWovqIN5LPF+jQH0mbX3jCAwNjpu0e6rrjh9/Uyz53HOvp0bcHHiO2dmMRs
jxAAkSDJvaBEwa9Yqi7mE6Dtweyu6M9i3dwONPrLFz6QTOK5FqizHVM/LnwBAcwl+QCHtNcPSPsz
NViMG9H9T5X1e4b+it8uMeHO34fPdbW1bEgUpIqYqLyAGxSHng5iCxHjxGz6pjynE4q4f6ip9RST
YGShtF6o4kyo5pnyukV2rkMq1/Q97jOGrMjDKb1CgWTz10xXxpV2iMprOGinPPIDqNWNAu/np8dG
9wTcwkXX9t+uOEjMmx5PZbc3Q7pJB2CY65/dJs44Aug2FPjwS3kcfQaO0/7Pjv7fz9K8B1KFqZO7
2Ers2owUHTLKwimXFoVyjK1oy3Ue4XkMqAZ54vWDdozc6pita4/EhaHogNNnCGCLCU86RxaEsWWg
VdwMm+5mDxREnlyniBFCqJCr/469rKWNEkPCsmTgXjYW+SrfrIyqK0gGKYhX5QMxmWhEOJeVA4rq
GrhIJvaEyugjDA0xTgxOeEp0xte9jLccfI6nsqhTspLCLmGJu7YP9LU0npfVKz24iztC32S6fFrs
XZ+jQKt0SaBW3UP/WPY7A/5IIdJIw552PdV8czBsDy0tXZ86yA7Kpw7VgtUPUNQ5fA1ee4i9+yjL
EZQsFk6dRM4CPSf/NwCBv7byTqTMMLo+I61i4E1xN4gRjtb0gSmueEjB8XoWtE2NoviC5w1RWJeF
93NueQMB//gbJOTLb/7bQmv0jrHSjaha3/zrdg9j2UOJKAIfHDFwY81hi3lcKtgT7GLwXxEv1BF3
yWX2sskRjR+JBoTRcXWR2asmSado9hCIyzCtgaSPJ2BYtZYVSl6y02WldDUPoBZ1aP/rSG2vik9V
cFSl+3/NGZnAKlm30PeatnImHd82uP7KjSjabIcPJxZxHd/cmvBnoJQ71ddH5XaY/PY24H4XRF6F
m+ZvAcc4RHfNViSgFZPDJHzJUaX3ETRf0hCUR5obetk1Oa699+oOgADed/RIcMF1BjLJATc4GHBm
Wonw/XBaZoG3P8xo6MfbU3aLnxSIm6lLVZ0zWU2tr9WhVpQd+kzmO6pQa0pfg6PafUoGR3QbSX9Q
5mHxyG6Ts3qHoZof5NzWPVsPXSjF5xaPUqZLGCFpVeEYracpxzLLh5nfNr228cKBGGWjlUDqO1jp
+6ECtYbhBoaQ9ilXNNP6hIrqcEpyiRIfVWunkTV1vEm1Z4U8MGFYr/rf+GwLz+xAgKrla430ngvZ
OogkaB0x7Qf8yfQr42yMue/SybRZfiKowVl8TyxhQ+HBt5Jm1xkMEs+ruUVHDQHoyCBVS8h9NaRG
+xWwU6gQh+mAyD4rpPkl/PgEHm6Negi+6lLtfNDngSG6bo/oG1qfCxFq8otnjYbfpt/W1zlmCwOq
tns3OGyE7TD9DDvfXVKMUvhNW2HsgVctRkRWfJRfhiiHIgVEGBNXFLcL2QxfkfEA8eDnQqwi1WUN
6J9hEqUfv6lYv1DTex+WOkpdkfxMqSq7JGrFWc6cg4xi0BoVUKYXnIDqFPeOglYrjQF0V5jlIPBZ
QvxbgdlGRJJTDDHkNl/2OrtEvQpcBqjiviC/z5rXH9+Ug71S6xGmktsOmWm85Pw0vSfvCTZSsfkX
svjsIqp4Wzj77OL/V03YInnul39qnehgCz2Po78e+F2glCzo/Mz4+TQGdtxNE+Zwq/4qwCl8orq0
/Xb3naSQKWxIj5kXhDiXVubT6dfiJBhDk7m9QNn1QUnhLoVv5S7nn2k6j2tM1gDn77Ee+Cx6YRzQ
Z2RPFwKSaMbmyqK/jq2f7pEA5f83dlWvuleJKBKaM6uoZgpVf7sv8Y9vhwKK3tFJQ5x1T8SPkB7H
Cnj7IKDNrMVz4KFuv6eKXnAla57zshSG0SbxXnUrNaLeWYIWHV6UnGKgfB6+Yfr7N1L/40a8dD9i
Ql7EGkXi2lHC1wYVR1MpDhxfQ+eQ63ze8Ixrc3Y5J4HJUvj/RSe5ARKCBvh4+QqLnFp/WJa0gp6k
5xhO7iggFyvY9y99ugPSoTf761hPgoIZfSZorsmaKT04ers2qG2kFLEyDyy/pGBaUOtN6cwvZQ4K
PqbFy8noSSt3IADB78oUTFrEpHjJ6cGZcpcEPgqdayzNhQRjFSqDSHGmyFTpqpjSS/OoWf5FhACP
M5uDew876Nez5J91TR4+5yhirFp5ToRgCDdeCK24QUKGWZO46KVcmClusy5U9/R56ZVnpssLT3uj
D/gjG9PDJnFjWmCVL3yFKMrDMWKWYkycD+/z+n77KsalJ/Cz2pAX4HROvYO/fcuJ/HYhNZlYYTx+
KwGZuOmATaoFdir9TJF0NR6tUb47WruzjO1tAi9W6OVtKkbpcV5cxm5qPdDSKrZ99KDbAKAdGjne
/JvkDMrC28MuxUPl8sz09hMNadXInEya3K5wn8rDF6WvP+r4MjR4Y7Rb7Y5Boxx+63r5gVe2RWxW
BmdHMFIn2KSEzY3i8xcR7and8SmiS4lSLItQBK6yk8V0tXP5A30hq4/7uSAPJttRdyFHGYlo6XZd
j5/17malHoDOm9fTvjc1pSmJ1nQWwKiJpmsJ+0WU7YIbPmsh4gL579UhTJmfGl0ACJ9affMdpEAT
tpucydB2i3+LlUUy0tQDl457sBryyWw6VHmFduwtZAKGHCeL6ymPxNLtHKrWpXiMW7NqJFzxIZZn
P5jTcUpM9VFSBF0tSwRleJdvXW6e9weP+Sp1sjCbF6vs7+nzfzUKCsimtM3Y7djei1JfABhQLgZp
N8/0r1btkcbcIAW2sxDZpdFiqRMZoco9bdixagncC6IbJ5r3qdGb1uN1Ykrhmt1BiQEy4dhyRL+G
PpivAJAPCtmQ9M9FDC5l1Jx04VhmXQtGFSQQWArc7D4OsqtzAgdFGYbxVdhysY6PFv91kR399fpv
m3QvQr2kD37uoRCwyTXHm7FLF9r6TOnYQ3KGsPjUW573A8540/Qi8fJOtlPcoQv21gtwYU0PDQYd
EXTxAR8F5ci4Aq3C9qKgmPh/vYgQOvPgNUeClH3ybUhG9eYvPZYL0Zg92qRNCQ/2l2O6dX9pgaM7
V9fLoHfQLqlHanJDUlSgFj1BtdUtz7irxTQ03RQpQDNmPN+qbSnI98cd7DP3FRsN/mv22timHLRQ
JbfLv9toW1EMaX3yB3oiBduHNTFSzEUxUdoq53NlFkGhIpubkEAlSZADdiG+9dnsNhxdRROarR43
ASajiqw8TIUkG1lOwJLanErnI6WUIp2WNadSG9aR8JDm6TcS+L0umo4z4pAVqfXmAHEiO9e5JuMx
Jg+Dh294mq3FVBY29VjgSonVAG/EOcEJ2nMz+H6J8BLrqMurZJ/+dG0RH3l1xseVy04kYxTzQqL8
RWJ9ALAsvUGkXJD/7lFdR6jC6YuNLUmcyk22P5ptHeW0tbvoLqXO+W+hNDRIQCI+0S152nt0GAo6
xc7twMWVXTTeg9zZB3zQhNhQBhRtrqH1xELYcfXIedOwn6RwyHnCcawygeWlXGC255oB7jW67sjq
Z+jHiTXY+1twMYP3rAoAa8lIIc03aoI3gs2GKvm5Ij62CE615t20XNUGjog+Q04ikdQoHQ8nJdfV
I1G6yI8NNxjv7Kx6Ww5wUWcFsBb2tCkOKLUmJb1CWAh2JMmh1xFcok1Lz6BAIY7WubbEEmIC4WIu
dQEzu/JixKFWEQDnXn8Av22H2eSWzOFIKUla28kWr61Pd7cVc5dJ+tf3oi+ag+hPpqzQm4dFgmU1
J1Yf0L9P/EXRRNL9TCa0Nc3aAgvUKyV0iUYuvehKEt7Pg5uYR53ztbRY1IBCGSH0Qu44pFiKAzpc
r6Bjt8InVxYkMFsNseQMh9K8pJcbyCmkG9LEylGxz7zxHTbAHB7Ahh68bhM9gmPamqtep0ikz7EN
sQndjUM265E7TJsjDGj3j/LrQF3BRnRu6KeacFWjkJwwwqsgew+toIelXiGqECCha+3KjtjyViMd
qeaAEOeJa9E2jqKGf1URHVq3lTUuAPv9EReSY6F37Guol3LzYLmHzpLLvHMaXJTJWura5f89UXq/
aegnISoPuf09LR1vH7QjsGIbQCHAz/fH1wnWQ94GooDsu0ru18NPEOdbZ6m5lEkQyRXKX1RCyfzn
8aYW+IkTz88nIM//pznBuqbr0/utHccKEllJEf7WdANxccEYdhmi+4oFa//1UxPwqb1oK0QK4E/3
5caw3CIolYJqr3XmpXP5+lE9g2P/wtigYQ6N3ek0OPgxILobmtDOsAHIWupbehsFeUU5hZcjmY4m
hJDfAAH3N4pSgApEvsTnTQxlJCf9PbArMCz4YXUQlqOvyotPUA1yuVAQMTowbFIsEWY0jhPkjJPB
pJuOBtEmVu2FRuHdEnwyRjsVWrDWKlOAxlQjC6Dq6fGLI2bRI0vpZkXL24ZM6t3pHrCVB+ifjB2p
CSZ0O9Nagf3vtCFbrJZThJ/y92BA12iyU6tFXhQZKmaaJ8iVv3CHU9OeLHSvEcwmFSY31todhbRX
ifOtzkaG+mQCsLxbjmfck49pKjz994qAdIFkGylIW3exwzGCqHepB9I56Xg3BFxc/xtdIXIn6y2q
+VKibYrQ1CYaCzXw2XzTRtvCykvfH58zIicYhlFqrdHefcQkq21rXuotgzP5j1ehWLNxl5H02cbJ
CQlZVbSUUGCYl1EUAjFFbkaK0DAkAvetuvd3cVTOEKeZ7658pcbXGvjbYiqwFjDRWm47aMmpggc4
H2NIrPaMYVFKsCweaPuVY2lbwgShJZt0CdJPsc5C0HKua65SJ6rMu9oVhDwkiZ12KTT8rfi2XPi1
b49+Xy8O499iHjDHVcEbA/Yo9nFrfmqQ4eDO6wtkN/T3QuuY2YoxF9j+eBc8A6DrD4jGfeAKVpED
RrYwADHGMe2tpv2PsU80TnGBt0IHkcid/wa5t/hswsi3wAlW/0Id3ZE+3WCzFcgZrHLCMrI0DBku
HeRB1tiSG4c1iAsSn+OMkDRKTlMUZOzkvd45oCYDH8SEsdSgT5GgSkQjKDrANWV8/zNueHpKTY1u
AbETDB6plUgyKI/L5NIhutE8SuBBn7/zpyondmAY0ExxQX8iD76/Uv9oOyXADZhhgI/vmvEW/HDP
aC6mPL5hN/VaBtJ4UJEU5AUqioWFAnNWABfUNBrSGNAxkx8Ek4M7fKq4YzLQyj6wtPcuiGEqpxU/
Lw1FIteFlfGxa8ktoaIpwqjTzOM06gmo5fkHDAFwcv2A6bQ0FTi4AbSKZQ5ZzG/tWxlNtHD6S9Ti
3j1xx1/9joU/sJlTOS0LSeLy3KwSf1r2IrMqojXCpZ4b6o8JonRZD7OT19iG+c3akKmB5WL5kqfy
WpKI519gwFWJcwp3282wrOR/McqFZiPVzV7jLTy6by/eoYV2EU6xxBHpiuz1YuA3X59JytcAQtVA
Rta8qVePswL5YgFqvKAw79CGXVpI4DtRwmLdyAn4d5C5yX+96O8RCj+SxAvlJeDycCxrf/TEZ7J+
8j1EB7fa6FC85Tt7JPH63AAcNKBwD71fz+CvNynLVY3d9F4ibxd1pR08JuKIhh2744o1uHgkM8A2
SdYjd27YJKLW0qFt6uXcNwIhwAOv7vEhgNkNGEukVY18Vk3Ifo/yZf/MlFIZHzJ3QESFp2Wdy78Q
eYuWxaXy+xyY3AJGCzr5najx6Ss0DSVGHDBENLFA5wiZoKPgfJ/0TZ74KtESAug9OwhscbVsbIDF
BDRQEYdvIUsRUb9cMdN4K8RGC6kq80dF3j9kK2qyM+dy3KJqBTlBk4Q7YmaR6Tqncl2/nNWn6JLZ
EQUeqryWbzbif8hxzvmGP5pA88nxAU0iUX6t/ukripQCourLSFNdTgWd3BtN25K9MhvdOPYFDCE3
9pccQ7+11x7WdlUdqJrb/2cO5MqYFjvtLAYNgtzKI3T/b2AFPkvw1LS43OA08hhZSsnIC/TpcNSq
6uEovY0TTTCzcoNjz0018/5DaBrcZgfyllTpwFeSh/KfJuiY8lU0fHP1mgXlIjnGGd/cchGkfwH0
aHZdk2CxJny2DiSUJi7N3EimnDuqI+GYMWJq70/vFyUVKXhfm21A1tMkkuk8S3nMRR0LMAJnDJ+x
JsgPH/6xVKC4amooZt+3SEdy+zJ/4WfNibnyfhreb1oMB6QCXqjLMMNJqI/k/HTSuZBDSmlHhT3a
BXkH1cEN88b11K0tmj1Q7ny61tus9sfZcKIL+7wXbivbwI7geWTBsBF1QGclW13eEG96tUmhEtWq
SVA0AqlPpmpOYuvwAk6QM6pxZdpJtDTdsAQFyeWdTRHqR2yEPQ2FCzFGDCX/n5T//7CWZxVV0nZk
u7YBGDV0Q7AvTnE79tFigsKtXYBc+6OBLp2s1tOlSiJc0BMQ/L/lRwAQDMfWSV0x7KSX+H3S+gME
CkMn980jHTEF7a/WOMZ6MzMwRvzrvyUBvMq2XnhQdOfSrxCma5TcRb7Bx1HfmFmSrRe4GCrhP75a
6Y+/Ag83O8PGGDa2n7fhIWEWcJqJPHGbLFK/+1G4i+kuI1SRPd+WGRcOvVgNJWACp5zv6DTLKozd
lriBI0qHP4jE7Pdw5IHjeVatIz9nRWQkFFYQALDje8U0+aAhMi0cn70nqh10NEoXL1g4x9ovzmOU
wgjw0cvhvxLXY58g1c1QpBjAw6QFCOTz8G9nkiz3Jycm6RaF87sGQUk+rhNhruzPKpBvpsMtmaAO
Hm4YuxW2vaWvN/uQFRxyKhurAFhyDVKGfd3q0lxV3v19eMEFvPVeGfOIpWIEYwvpm+2mrdVfamSv
Qv5WgLy6L8AS1FHF2ocAP12kjJUj6BA7RvipY6oohL0/qUVkoENdTuKi+kuN+XFnBxRo+2hdlXD9
Zl1erzHFhXQlUi6k1d65SddUFWVq8lYT6CUx540+JM0QsjCCiVvELtzgp+02Qevz6NwPlZl7XL8H
tB0MmhXQzrSNGapPDhXpunBVh/KrGAp58MzvrU9xyU68O7Bxq4TLf5KIG9IoWIOBhZ20Zdt6JXXB
EZLE0Qg+zdk/MtVrnrLFchuiLd2VmVBRlPH+RDGks8nzOXS6fZgBU2I+V9Hf6upKWWFSSGAT2AVy
fwuSK7uF9qI9JLTzPqc5TF1bDCU5SFMXg5P7QnfAeJEtLrzmDahEXnlUES1CvC8/nB/Pc6B1Zl3v
AUGZ1E5KAc+1ZMHZ3KHBRVQ+f/F4Z2XH4HpNF31h9kBT2G3NPV7F1s4yizUNhVGBr69Dhvr92Eub
SaC7OliTTRI2wzTpiUuGyBjgghbxS1vaIeDMYgrDg4FLL5CKXdF0R749WuGP2S61ofo5R+KItKkW
BKzBVtX0raTFOvoqWNco+g6f62Zncr7dG40e4gNRIdEwwzShlQjKGZnxj06l6snV7rrW2IRdZjhP
IgSp+pFLbzhseV7r0zMVEg6YsZfE8zsnUq4Dgfvqlr7ffv/3UuI4kdlXtjZx9bqTMXK/LUq0hG9S
KsepD499ftOnM/k0X0jrx+M9wbAGWQZUFMZEFtiYy6PLMRVdCg+BiVYDFnEPSCoxWsxX9m9Vx/Ul
V8vq7c38J+jvJskzKw9gMVwCOcum4Cj0+4G8GXJfnYFfdP3BYUjDMKbupsqaBzG7Jh8dBoJHIZ8S
xkjGBLfAwQc3Ejq1PchkDK9c8hZkYVM9ft0Rm/z0oeXZ1b8O5zi43pt7JxZmnIdFRrmAKhD7ZVle
fkAi7yqld6Kal7+vSzBkxmYkrk1u+3mUqpAXCvs4dHY3o8xQ+Ab2dbNIjG8TynuuE5d5zY2djvBq
2sskWitKkmfTlsq6whWsWR55T2UuM5kPvN+WkQxdqQOtESUerCeF314zzOjdNfVzUg98KL0V3mcj
BegUxZPmSEF1Vp0PYw3SPyrPB1+ng370Kp99HkXvGJsF+r9tdPwsNwxXUPJHAaix58aCTEmipgmb
++vrW9ksr7xxCJUJkIE2Ka+SxHBXTkL6wysK4AyqYyNVac6/7iBDKLAihBFD5Q+Ew1BvvQ44Vxig
eWv/pvyDQhuJ6sa6DjCwh5848RkBZCdGr+97592FMByBOwV8YruE8rKQ305xuqgIJZbWDbu13ZLp
YfpfrNKjQZUFiQ3Atw3su8XAzOo89xLonmtRGqhs9nDJ0zAT84oZ63O9+qHVBzg0QDIgzmDwxq4e
ibzJZKERjihwO1anpAOXAFZWxrOexWKGq0QSD7IiTjuCb1Im4knoSyKoNvlVYHlMtX9TfFIMej+H
tFn72mgOjJv3IDptmiEUTQkNxWuM1ygg3RKezkixhRHexK3qNEsqLMajPZBjFcjuG89OxDOWBLKa
zkNdSgv8Ulf3TFcKw3mXzG9f9bB1rFZy21UBLk2E0ACmRgRxpNkC1422YDMq//O0LW8F+VPZgjG7
P6l5Qfiv29HVNPnkjYjhRjR0phjwGz10OSpkRFWzGqw0pqUKTisQMHjxgs+rUdZnS5e7z74+jDsV
D4Q2YK3M7eHjkM7x8ShpiJfWZc15UkXKnndYC/5JRDaj0xnNSxXfEALb0GoM09GcFsU8GCQug4RT
hHSu1bbyrMK8EIDipYIlo/nilpGV5HMeZsr12iA6xFyMg1F9KzL7WoThvIqdkEUiJ7M58u1mKqc8
HKaH+NNxvpUD+bWb/WJIZ9aUFHmYy+46ok6qo8aWHISF3Qatpz0o8B7sBAU1SBUai4DG1lWLz7Jz
opGwWv1d2fQJ1bbGAKPK/MDQeQmtBNkTWd48MGkbPeHyK34irJ4JM+zAU+oHAHnfxA319kAWq/DM
PSntFsiTmzdb8whK35d8sXnHYes9H+iG+hgGDQjkm0BlLZPz0zmVxNkPDQC/XkEb/6I2Uds9/DJ+
dysj6M7Afd3c43pFLpgXnyALF+A10c+KS9US4s1Cg77MeBnGQ/U/mZX71bo4JtiIMpC1cQ701E7S
/rHIF0BdnlYwq+9j7J5sDD+BhE8TGLkOUApf3S0V8wsXlsUx3kGyQ9hY71K8WjdLoRYFZyaFT48H
UkFRCMzuxe527y+R71kobx1h3Weosrv86tqfqTj+QNw3cTxE1Ual4yPrZHehZiTF6KE6bqwTL4mD
qI3PTa7F2yMmTNFBhu2LlUYPTxLIwMDdSK5yyUttn3wHCP1Zk1HgMvFS1seRsURParbaeXVXTBUG
xoq66PwIUHe1fKxYKNFd/j2AW6S/GEyx3GeopA+biuUc1+eynEHHzUQzoCWCOgCyLVbao7YMvM97
G0zCf/lDerwClIgZh0wYcmhwVExynhA+gtdFS5WwiLYpWpOZCf3CKH/7af53pU/MQCRXMYexllav
D1CMgLaQDDCGJnWZLIa+y9bK/N6l1QKuSb6DYX7o/JUUvNw2FfnOFP2oLRTKPoVAYabvZJs1xJ6M
vC7QjehYtEOVIsEnuMUJLT9FjUNvHnjwI6EAJr/MQhU27uBevp9855eIna8fUtzBHwHjtrYrIyLS
gqp/0/woQVxvLpqz4Ca7F0lHLWvzPcVAUfoSFqSKQ/Y9uR6Ykg8t1BJpxk1I9JMZAraEgpzkUgBH
rw6Ie7cpMmIa3/h6z5P2/3LLHIc81BkoXjyi79Wc24Zy3fODCn/6DLZESyRB8dWn9C1pPnEcJhot
Diz2PCXsQL/DOXPe+oCpvGQ628FjthEOXz9TmEGtQflg2SQG1C9+eApIL9OSD30+aZhzt5yRjdA0
ijqJjUQEoYJ2WPhnpnfT07LfShyA19hAAeBHKvrAQf2Fe2uslX7aXLpnLyMUbidKYs2fsk4zjaD7
X8tyy6Y+D1Dos/J7NX3RsA91FnYpZtrA8FrDoPZashdkcesyEfKC+26k5mzW3oSDQKLYPwIDuUBf
w0fEPIsUcJQQf2ZlUz8x+ai5Gild2Sm4U9htDJ7cDYWJ8mCZs4uDPD8yeyQSBQagdZ2HFg1fs4L4
zkpnfgJ+UJbcoFQ1nbUt6wMZy/VDLi+YeCiCtufU0VYV/LvOAYbpZMeYCQuqfY+hQtoqB7Eq14nu
LeQPlc1A/zrc/K7TYD+MbpDFDzxtkGkqqmzIZPV+DIOTx+zWqYsdvULWY/DUU7DWV6OEIcIGGxES
6OXriLpE9+kwhdCcum/6YxPY0Ig2kCTpIY+UAXQZJVHHecSiDZ4+V+HgfEYiOvvpFCxJ0UUaKcrQ
zDccSEDmrhg/bvb4l8MqhfguELizjMsLZycRM/cEbiOjnVOWkdchD6UgROMrQHMG3WQEdgqsagb1
cqh5qw9ofxyrPFzanNZsJX+dT70v/0h20jZf5tXi/078q5RSbL/jcTGPQwSEv0PLGTWCOCV4wya9
vZKai483mOe/s96rtP4Bs3YxBW4IM/OZ9EkK8enSWqY8AzZVAy+lnRbLgV73F5ZLg2zi+rq62Rdc
+aAUXGCrcp5aHyz+YG1u5A/cpidVlw+a31kCkBMIZjZDzn2tDdiKE8zi+GjXul9aY1nfVMIlf/bs
NdGIg8TKjn7iDuY4+/qtvtoGlgGY8vEa9zX0tunNbkoKhmcoVouzgRhpJJZvPRE7JtcA9Qbb9cP0
hVI1buf066DQvBdcpbQk+3Sm9/Vgjf3DKUsVY1JeKsUdkhQDHGdjn3ekXAOiqtBYcvjqOBWAQnRQ
VIRwemupT+05sl1v7kv0lDo5gkvB1jjEKs+EirJeHmIZ0ZhqlAGTSqtHhekqzZgeVpbxp/zBLnBP
ZzfTET0E4q6o68L3PmQdiQfqfgto98gzXqTO8/i6xlIOwSNB1UfMKqg1CJgR6vBDytqQGtgW0yIM
Cals1he0kSKNzbn75l7TeOCUkBxVaPmQaDUGGPRF+GaEad91MGg2KaMg0LZvRfm/NubWMedgVs2/
8kRv3wrskZOd6VOID67jzOBHqA8Pf56Sk80qHWchewI4Bo8Q814Hh8HonJDn48eLGNBOsFlt+6Y8
p9FtImgq254uFF2MbqebypK0cz/MFhJHQfBMRmEYGn02htrrtQ+WQUzmm9oO6WFRSc5eYsaps484
+J0a/vpeHC0Adp68HIA7K2EdjrZRvzw0kA9NRBVIx8pVyirioLe3szg4BUkuMv89uWuuXU1lv1hR
9RBK3l6ChCn1HFs6b4FOkFrqXIJFU7v7y327kAkBP3yW2QNjrXLqI/H8UzLa+tOQGel05rb4k2k5
9zWoqvgAV/H+LM2IilIJUmFqJZkC5JbhrFy1D/PRVDRNEGHuQUTthZiHGfsODM/s1hwBtsespnnH
k0qnH9/xKSHV2JUpVuh+BW0WemUZyTvAHKfNRanNMoD4I8UJKNt++7GPUIVR/CEI7KSfc7Ynx7iT
ITZVEUEjuGvqFOo5W33AHz6gI5NyG0zjRAnuvNAHr1VhbtTUkHcV7oDmnYrhAfFwHND6jQ59XFEx
cdoJ7pa+VuQjA672IFFpViX+mAD/oHcP5q7UKajdfDfENwMOn8F1/Hhs8M+29CKIGG6uDjFr4TDD
dboTgPgVUbGyrT/QCd39fYtVUCMGRKfr7LQcHw1BDIHL9OzrQNaW3wvlQkWAuNufSLzmNftpyS4O
oHxhDRzHbfljfbh88ePsGIxuOpijQ3ARJ/hdYewgeBJYBnRHcOLojHfL1V77xPmDFnlRi6eHzwmO
TQlFSB5aKsRks5ogmYsgQaYHKNOHX5LP6bVhRkQiJYZ7eEJ3lyW6LTSLTQ7mo21bJx840TsXA1RA
00Wqamkq02oUcw7lgH3D5oIPefRJ0CEOh25ya+HjJpJQI8EJX9OeyhxjFwhJL2katIW6eqBpn3XI
391nJ1Jkl83YBfSM3XuVyK4/DNarTsH6aP7TsyAkQgq+bTFo9ZFvZW2IjhpzBIbVvp2bbQD6pj4Z
t8NwXLkPG76tXzveTLLn4AzpJr5aq5o8JA9Fgxw3RVSOegqQE/uJWzzOF6GR+ZFccFSxp4gVAq+k
xReoJCyFNrLREqKDAIS9BpnhaS6jav4saU2X8mc8ifcsMzcIv5Qmo5HSzxPE1W8TxO6w757RbgNC
S5tcqLlBdLetnoaR2CpT20V2TiRpKAum3LJ0QiPbOZ4wKfBuJo9oulHNl3QB8NF7kd6q7hkgG3Rc
MKh3T/uHFQEVOmQj6Tp/U6REORNrjHMgaIKK+QQWa422ZwUO3VxLpUG5zqMfS7QAiGu2BOprp3iP
p6s8kQuBottCJQpTZrm4O2UnBB0GbWTNIIq/R8VWx45MwGmhzt0oASpun3LToIrnDGXIolHstAfN
6Bk4xHzyJGhFLgP2/jVbAkwLEixf6XGn4uroSGYqBRJVN4gcRhoL2RGUcrGfIw0DNBJY/LaE70Id
SNZCx55nrWwKCE7TjWTi5GZFCZNqKy0iX/AGI79931xFrckkWfwz+sVp6WNoS2wNgV3Wjr1S7F1T
SlNo6SAsskMKckG4VdwiWjKy/yYqqZX/oEiXD+zMkEro3fuMThUjm8RGHrzl4RJaoAvRrs5WL2FY
bOkgiyRSvXIiBDYFo93ZzOcs6BiIQrC7LMYRQ9tAYeas9bR3spzKq+WeDkfYJwNcLkPq1PBfWNQp
Nd3NgHUjWzpQr0NWF4nBx6IjBJutaaLSSSZV/sSRWk4HK/1z+4+8hJmqvwM/JShsO4raNh4ciEUH
AOgKdi2taEjeCQbyCdzkgUTkZT3Kz16RlbZWU4DOe7NXt2qTi0wm6MNTZWzo+f2aQXeIGb4x5p/C
APpMncpKo9/rihVVHnnShHmiomYtkdr0i6aGrdcY9BZjVg4i+MtYPDtp2nBScYG1RomMBv8jMxEt
I3/5UoRc7tCsCc0i3l93BmcgDTsMc+xNRuY5M+0TSwcLi6IZtcL8VzZijCqE7qp4qw1Jo01OthVK
MQIvpJYgPAeW8NZ7R7KfbSwPzOPFmY/o/2x/DNmWanzrXO+Zk5Wrm9LuCvF7aZ6mg+YMgLMow91E
lHXMFUazE89KbNK3VLLo43hCiK8TLV5EmAkjP9YR2jTNsypAPnGwy31PGQJaY9eO0EpxcFYTCEdn
rKwOjeLca2xqtMZd6AXjciIeGM6ZbbBrF1DI3/0e4u3D4qB+JMsyW8uVOEjjIAbYCYxhCudzWiah
yXqnnOLxqD79rfY3zfkotGerNEPywTOTkHPfkDIAYq7StjVm9Y2t3Eu6lWaxv502TTVOGRFShr/A
1uVtBtYOU2/x2Nrk5Gmml9szVw/5GyC/jw9G9qVrly6lCcFtxK49KOavx1Iwtilx4lm5vbJnHs9O
tujSuEBcw46cJUkS5KfXh0EE385sZ13hftkBrAOJAEEQAKP39Sh3Cb5EVc35w8ygajEs6BfC6YUI
7XFfVGQWxH+eFeQwNvKoamlmQRJQ/vYdiKfCoDBHyC8RhCD0DJ6AbbPreRPTTtr94F9DiKqRjPNC
I/Z+InanoH5LQGyhYteVDs2OTNfaE1fJkGw53b2b7IQ92Mg4oFqyLiSK8LyZvMqzV3nK+8BS4Ypp
PJIJlLHbhPxAc036YXz/uqhwqUiyZOzfzbBoGNCekB9si5dmx34A2OU4tODUt8mfUQDCKtvM8t4X
9KTMHGBtpji4ZHO6JxRezHH0+1wryUmuQDFmPkTu337JU2ngN3NdyShWxa6DB02T5eg9sDhi92zw
OJqbM/+KUEg6MxFTpvkhdUqSK6FsoReI3j7jDIlVlt8DSCtQnVJkSoDfbPfKV8H1wzw9NWNjh6yy
cSHdBGF9co/YuECcYJvThZB2X5vF/x+7K/YcMpi4afhzsaXVW494PqH19xM+Bx7sx6uDvlKKAlQO
T7cLQcNYbjAmrOGgs4Tq0CRozsm+wKfuvH/UXqV38P93wXlGYwCOsd9UdKTagpSJCWjZrH2M6zeO
dU753Eyp5xETnGbvAoud/1YyQvI85vXDqZLnUQ5EfuD+EIyZhvsll3TCYLx176kNW9fnvV+AF9S7
v0bbComhQTZKTi0lkSk8VqmKxc3xRX86IURYkyrNBTnyh8rCo+fCvo9UclqAa05EBS+fhjdMwnRo
lXJnqJKakz6z3TPuUbvztl/0puWuZYWZmAb6gKQPDBfDpdG2n43/3BwwoFO6ajHTmvflv+LVxyku
9QXezWxdYgaL+95RLnVTv9q0tBAd36RNOGDJopIvYDtDcqGJWmUxtpM5+vzr2ztUlJLTRfUohP/I
DIyenvqPi9UqRwQV3uyRCoSvGE8OaD/QKX+CK1nBAbVL8kUB8BdPm+Tvg1TmM3xvJ6xbcDXpALGj
Yd9L0wWRZrvx8cUkI5TZp/hLOlRmqjCnDGUrzklt31gLholowd5h1ZSeQnBd6J5CyQjNSA3SFjb1
yccbd8xhQhVQJiCzXv5tR61QxqmyKlAmiGE6rcTUEekFnIT9SihkGOxeyK+O/s9knfn2xK4yRDO9
M9BUntrU6sV8d74s/DfyjEATGor6bibaHIQ0c5xcVS31hkGRi7pQteIW048bTS9jtjVVMQX57Onb
UeOWHVJ3umkq02zuJnQ/xCRqleDaHiWd3kUA5XYcOg0AY+WKjHJzysG71emhrFiGTeuwVvLJfX9r
uDiV1xd0KdFvHa6N9BSIgMu1sMLZ9l8r//p0SB17h0C5Xl7boSw4TBzgyY+UZ5U86n/0ROyywyhk
Il1TQEK6ItlNaK4wzIcB8z5UaannuWKrXxGGc4IqekzE5fAh4WsRRjWTHlQoTU5UrxagD1Ykh53B
/OobDL8SycH9u0l2Dlw4+cu3CwMndPhHGNopXZa+UXf/15A3v8i1PJjak7NAEOXjCgqCH+ZAiLkn
GVXVT/0n7P5eu0fkIRG1vRGAOgZvjZAnYbxRAutj0n7CQ9Oggj0IIOZnwpFOpCQuUVutv42TdPbC
gjUeuprvMjw1PlToBasubMb3rFURxVIVQocFgINjqMdj6lFGChb9MvduTbm3eEcJhjmjzCa9gCpm
1FZeqCjTbCuGPx3XyrRhQoyqWOHxclGj/HLCJjmhq20jYBiBdNyY1cmv/MrQIP+9WPg/GEUgohBh
cTIMGqYnNj5QzTbfPtoF0p+HFnhZQJEryu/Qcz3Bpc6mqnEEfakELQg0bMfEeLbSLSoqzxEKWJhs
l/FWaoZLvakcWmKv53SR3cDySgAqZZ8nP6yOSOLux6sa8y6/XPQezgU1fEGB7RnrYGYG/aSaDQ6v
WkEXhY/ls4yji0qIJrSa3XbIoU6KdUU0JrXoILOlafo2EyVOWjCYa1m83+i9GFvhfZHvA2nRqOhG
+ujH9Zq5XkXIKP23OZft0N9VyqDpeH59JZ9sbv9HiOzMyaqLA8ohZrwPIPIB9PIca4bXuThu6wuA
aAImyk/km+TQZKoM9c3G3B0V1dTE/1HOZVC03d7cQIyW4ujdlmRBOnURvI8LqXbuoBZdXd1Fl7Ff
xOrE0xLLgrcy8oUmUwdYrjntxz6FXgRwvj419aug3smURmVHXfNBj/msIk9ZsTXlfUYTK0cIEauH
t9uzy3q+0wGG/GkWrVr4c7awRxkui75YvnMlUlmmMfmB9Iz3TjLFO3RSsYsA8+s+lItzK9DBiLo8
hVD7jk9va2qf3X+v2VoqN1/atjj2FjG0rW/TN1LVmvEoouTcv1xHbZ2smWiEV+YokeHQzwxfLf+7
CiPQq5qy0Fn8r2iqU6tS2ln0OESVRPEEttFY2EGhqldHypD7EHoQHZ5MqlPT1FmS55LHglvEuW0o
Nyd+TsXuntuXNZJkmvsL6Ks76FJ+Y39E0aro1Rw755Cy3CMu1wDrX0P6pUpZ5Y5bx52rfNNo6XZb
vdxFPE/m2rfkyD3bBnf2DRFMQL0An+gY/Z/iZSvYbBTFsyxUXvEEM6vYQtKiQQ24Uiiv7toLiKup
5TnRORbBKPdBaW6ARMNY172Ltysygg9TmdZvg7EYd85Ba/VUH63s4sZx6zjgM3aMFnlbi+vyce/R
WfNsO3Xeeug1UdIN+cSvybZto/5KHoPlSyHosNaiC7qUvY/LwmTMa66w8en2ugoOkjJRdaEgfS/+
WEc0dfS4BWTapwHTwKieDT/JeujoGp+EkanWtEkYfcQVEx6TGTMMQ8VSos0yDGzFP5B/Yr2RW1kO
1+OwZEngBu491FjRuoEQTp8z27vsuZAugz85VqXpJKF0RLmxttcGJhRFWLY3X1Iux0gw/flS8Tdl
9xKYqpxDFXJzemntLxS976NWVbwhpbGeVDPfxfqJ92HSSv34X9hgY0cAPTbFVoLbEdfAhYgOU1Vi
g6A+1E7Bs+q/67wCYbkhc2OsnsdMBwND42CZNF4PW2a3qZqaMVSqRxnm8rChpYRBzo8HmErhNAo+
dTAiPVyuaPWvJB0KA9cllF26M43mZI4xgE+yAiMyxm6jIK3eE+Wcic3w1v0H/NSo8/0HxAHoreWN
Y3RAa3HOFvXfrekQiC7DeO0MG2Ovi0HF18vwq0k8RJ28oz7Z23pyPREqeGOpbKA8ryyvC+IZPi9d
akR2EkGdytH3JosMZ8Wb0r3fq6z5DHRmpwkhiB8lUcI7x+Spa3gZ+Qqos1dQ/IiPhcEBRrL0vyFh
ZtX/B2eH3D7MrQYmXCDxAQdsV7bgtPM11ufuh/CbiT3jKHEpzynH6kU02PYjeDgNrZehDkqG+pVm
hMI739izsP5KQeV5wrif849wx+W1dmFm8/+oub4KbLd7yQtkw5HnaU32y8pwsTPl+hrgynTytyu3
Bk1+BuGcg+RQLRhiJvQfm7sDyc8TpUvw6K7x5fBV+EgAdNODOGQjoCKV/hSOCdnh5NGiovVDNoyj
5Lpdka1XvzOZ7sHZFiOFVSg4DSRiAnVfM/YqKEEt3oqc3QDtj0lsQHd8OI7mupncfIhdEfxTDVDl
XaAa98CRVDYtfpKWVtuR/SZz/AbNBsMkF4oWE4h/QxjyF5Z0X0STpGJEjPnLpVyjFMMxDiifhZSS
KR0JwgdKzPAHvbHJzDiBxjE2XCBIb1gI46YgGAvoPS7wCiU5SgT3+UQHPdtwObrDF50mZds7Vlty
EGdgfYaawoTYeK7hYjeskcSuuq2liFijAThL2AGp0Y4G8girgaqzF/MGDDB7/kCtxDiUxyRgHvKL
CPPJvx2Yt0VfeZOwEn+NJZvV12I/ElhmrrG0qFW2wLXzyaxmzqHNQ48keMFDYLTlWWpC9KE3RtYR
6712uL4a0pMUGoJEyX8uPRp/Iuci6QjcNoH6oEG03EQ+o3U7xTq98Fm9PFtBnoCQF7ccpLj8RL/e
qlJyI4sPa5L9hg7F/iApOeIfq6mn3ZN83smNYGDD69lfGtLkp+hQ/G0lB2R6NrkZ8V4nxlwjypQX
KX5y3raozjGBzh8yqwPVCDdckKXCMo5cejgAUASDwEqiiePjR6zO1nKY2SPYcw9r23sENaZnMYZV
ZrNzurRRBNmdYHL6kA93iauW0OuQ1qCkinLdLFrhYauQs/Bmulljq9AM8lTItSFqSgKLhp98uroW
LOhtIX1ggNbh3lm5S7cSaEiTV9BF7tWbVtK715Kk5N9Oefgw4p2GYqI+Uz5sfbbwxVh+B9/eLQuC
N5EUdMr2JOiJCvLD6KgtbN5WMWsCLCz/ST1FoT35qVLtruzeRQfCC5mu0hJpB2ZPPBcZ4Xq0kFb2
pqlv6tSNmp7m+EEVLn0UUHCgsTp7WD2U7k990SVclpMU/FGpcNweIz3fYfl/Pkv0FSjZ2J4uJxIl
r36evNRDjkXD+4VcEOQ8TACfULl4RYktY9GvmNxl6KhXBvSxYvQx9V0epVPzICl5G/GmGq29GDAv
4ZcmiAx9F+b30wBFUrgF1ilK3Qf3GNuFOyO2m5Zz8r2NW/VftpAD334+s3exkwuohMZNhuQ+0Fn8
JL0sNJfKR586h8pZu78L4vd3nbslJgt58XbQ7M5Cu6XfPm894bYRWwqsYzLr49z8ivEoLwRDiCYu
WX5SHAgzBTIFm7P/OkeKua5/DofHvvQvRZY1+zsfDzzC3ivYPcN4jLpw9JmnaIkY6LnrOOM3+Rk9
ZUJRrEHPhwgQkU/8YRffQcSobVvBjDs1i1WTyNegdQxOxDMIzp33mSe9CeOIxvh31AOeLuAH7eqd
+8MFuWYUwOAgkgSostHctT9Pg0i1rZtq7rSBZhR35YtWh3DNwKplk1MVjsC20Rs1OFQKkUALLINb
DToZJq4q6r13SCAu+iJUa8l74IQ0XaMwNgtiO2zOwW7amcIGwc7rsnsIjVVC0YPlfghA6uGqFPOL
jP60F1OwTDcRtK1XkpMwxsvzbikMH5XqfQpcIsIMg7FXRQtFgURvwUw/wbD04ZPX2R+OZ2Zc0NP4
5XpOkhJi086in92M3HdiSZNKfEiBW+vwHQZwxwWx65xkpr1NFsI/QQY2WEFwT6ASV5XcEkEQyzDM
b+mYm1Z9MKCu0wsjCAX1Z27ZfjIz4imnHsbsPWXthOi0shWu0R0obBy7pL7JKctAg5dkKHFXHDKU
oy4ybcmlAyy/QkiocLH3iDM4HJwv6kJFo9qP4FFKReRJlZcGxZv71RV0heb9FqhcnHICW3Jh+ERS
IYIZnZ4GLaxFKrN+jfN2IJCLoM323zfXFYNmA7CG3MOz/9sgoJD2AtHS4ZEA4pfY8J47LtNEaBXl
6BYAj+AaFrzDjSP8ihyEhQ1qo/b4xd4ZIPdhJo6NKJWKwocJzKwHFuL3r6c7C0sNNwQuIVTAhguI
bfvxSwIY1+iF3AQMHtrbzwFxa9kTxX/5nzO9y0/l+Dj1xIXi6lCd1zmmX9hMQNvRUgoMJ2MJDtME
jYHsfRFyOUCOaKC24sC8l4jgdLgHyGZyANsQUkPbFB7klVRe68uM6GjzxQ2quLhFlhboI2cxRAMf
giJcjmo+MIjNTrsqTTULUcSS0a8VMKpBiWLak7ds1VKU7TmiuutMN+q20ibO0mEuW2cALx+4V8/7
m/S0DU2KQ2DAYnwjBmPdwNisoWC1aktcPcYeYpd5KtFv7eW7/FDPI/nSEGv3pK2YDV0s31DR0aJm
ff4SEOBRkeKqyJz7Nn+7zdg4kOq7dOV1c85DW/g9n23+9Ow7S6v7j9hTfaXet+p2YLbYOFbNBZ0B
QIXqSDr25GNTzVljqYpIf27DepVWZBkdZKqwdo0CkM0RX8GJEs88w6kZYuKtpUAZ8OS7BHiwpjaw
ifFWOhrYZeyFjXMoanbi8NB3qVz0wwogkWF+fBRWAh3jNLKNDtBXrS+659OemYEoZTgZm79n01BP
W74i7kIhOCn3eX0KOCb8CprhQlvDAkeHvJKk/sZStAafFvpeFdk9udZY707z/ZHeZIvs9B2abnbM
71pC92S3sRi41C+GXXvB6riijShN5uSKzq5jKAQlfFbLvZ0RZpnlqEkm8+MDlP2jqD6myyOCFNaX
DDRrZ7xB0Ns+7LrdFU/ZIYiFFsFVdqc+sVo6llNWK8KWJi+EOP8C6oAOUKwnd5RCgGsqvKhE9VRF
4Befm7eSwIT4phNyUAfqOmdvbTbXGv+HAOSBGmjH+RAJEu/SmTl4cxRODIlKX7Xu86a4Fdxn7YOF
F8sfYOKrwgxZbK7VCuPiBjiM4lSNaTfHEvk+4/RXM5dZ0Xn3iJKtLkr7NfnAG9UyVDxDUK/difJo
F/cAkxPXcx8YR4iVeHXlV57Dm0WODbKKpfgRzsLoM1myM+GBnQ3UGhZtScsTFQkQoRtDMoVx9Nxc
m29UVz11IGIosERq7FymYJQCa1Ho5o7cbZ9Wwmm9EvOdZKUR5OIIBmVLr11NVGSon2JoojUWU9l0
SdVAdBASdVZJTFyU5xSjOKw3Dtl3khCteZ+UkbwJ50AJR/hgvOFsspOBdPfQy9VOx8RWjMw9+e/1
68MGppyui5o/Jz/M5YRx66dstQz7yOO1eIsN5hEUgp1f1DWcq22ozMRo6QESBEMTgs0SKyrfsalp
ZssQDms95R9bDyUln2wCREG6MFh0qgaa783JQBxSOHRtkRL9K16Wq+6Gb6XhVz2rJPF44c4AhOoy
4srLSD1pCTpqwByN3D+FzIbq41wgazBSK/x94GSR64nXRVEIW6OLGsDpDwgZ9FAJnECRvLoVY2SA
rJ3tl1OwdusHDi/E6mmFKvf2d/puPHD3VKVq+XqGzYIWknsGsZ6dvJtRKQ1uqT2mGnBJOfFKl3r4
byMOhiX/pn7peG7zp/euVTxzVXX4xxzgVCscsArTKUlA8qT6iMun8LwC/DTxaIUe95Hac7Lh0LCn
X5RY68QK+jRFYfZm7OGakLRjdrND7jIyF9W649jWjQARw8NIesHD37gQpeMu1ZfRQHYRc59Gztno
5QAuEzm5NbI5XS4izoU/v978YGfh9Fn60fteDuRWKrQo/xDCv/sSMiw5ltwL0wZJWDxGeM+kfC2e
wb/EdyL28sYkybqp/YxXuoeWpS5osnVmD3KrJeM0nP9TEPl1gzfum60ZfgKZNm24H6fEcca8/b3q
crI5PV6bGmCJ8zfZERgJQCKgchZi50mPOisSAPVTfCeiJErbB6WDJ0GV1VBmV8ECsfQheov/DUAo
z+5G61tZHT6Ro0LKtbk/azXpqegljkAqQUC2XXuSCt7oD/p9180HLyK5EXVMMKtDuKiDEgLoHPD/
L0ppAzCRoTFI+JCyiijie9FhH+fJv8DHUFJG/y2lKTVFA174SAocIHr0icavFrRLUB7mwIYkrVFr
6E9KJfVazK9nu4G0JDXeib2eOIOFKks2ejeUccucfHAxroUYb8/33FICDBOVijsRKaUoOHRrN0oi
in5Z0nBsWu7gRu3hyh4lKrH6Bz/4Gjawkcxg+HLR1vHGfEb7se6TCD7GAPYUcfAMiOARqRJa1Sbd
v6Up/Yb/wpiEDCCWK52h/fAyA73bDlkv0tomhauQ6XuIYxdyGbVWAtd5MWcSvgKr3sOXwEbyeRq/
K7lRktR8BHJu3wfiP0PDjNZP2OzHzCUTonWSE1NQy7yDIMQD3tgLOP6oWWObmtcC5EirjEDcH926
CUtVEuoz+T6vHezoeGY40GBuzQW5V+Muu/tqOfljTTONHpQlnfvK2Ehd/mCfJsv1aBO7iOSulek0
PbuVU7mIFmGLJwGjMUEEKGgnWPQfZ2LeDJQDD8/ksb/QfTiQEYKP8lZWdE+jvQGDDcaYi3pknRMF
ymZTkg/zbtcZgojzgRN0iOnHNnUL19sy2q9O0GgXNbblXAey5q6qRsJEJMdI+xWSZ/ngs4BuPaWx
CHOTKXKhCjeiqikzG0ZmH8usIYSojOiNes/RB4u8VJxrsSVlyLFhprIEVyfLATv2kt+hH5hCtOqX
1BorEN6Ww2rhBdtMiH83wzRMz5I3QqBz4p/6MF335m1J0iQ7f3iLCn+SyqwDpzmDTcWrE6C8W99N
Nep9fbhggq9is772ZeY1ccVVDqCYn2ynNQ23hZT+I+nmO/OH2xpvN/WnSCvs7nPidRWQ5fEvF/so
6+gR62dVOlzJwxg3grCB3eulrjsZbMjIhomb4KRIVJNWUN4hJrd8Kd5JZK6NoWOVZ+iQ3B11Ckfg
gHpVfV2KRmi2b3ZLgpS8t2M4f3TmK8LTSymV8XxTcOYM5nlBjbxnsUg/pvmOAmN8FdTdQVLriSFw
c7+e34kaeKA8aWE9DL1P4gm3SpL/0Cvo3EaK8YcnvvzLvKLYQjjqzzjhW/8ue42ecIGAB95xU2kv
gdbHA+G6gs2cV2+9ymomt1kRUTL9a9D88KV33rvZKVX5CclhPyfAqeXs5AkIkm8n6RCV0RFm0gtP
7ncruV0ATNM7PjwOMBAtCqFPcW8xgnYDbM3N+/0WEL1EK1dkXGtyrp5dhQ0PN9A1c4ghDw00FxJF
HadGBB9uteUPfScwQTChzkGH4fzWsIQE73MMWrQ4KRsGJua3rdZOCU5Mh2/gxO58KGDMCDGVCs5C
EBa7sqzzVHA5FUnKh/e5IlhEr2XOuRQTCfQPevMSbXuK2t7dxcxS4/c3avxAq5iKJloliOwTXdbO
9u2VS/dG1DYphZMQqecS4oVxFYrGdeDuhLIF1Q8T/0j1tLIsF4J8IOUsW6SlKTOU6JnmlFW28OhU
ZJKEfKQVB1l+1yei0xFY2ANwsWzvDyxgjA/DEsK9aTG+rbFlMhrHuZaSiih/QQaUtGwy6jPGK+Nx
k3qcHPgRjjVlV7G8+fWlQxGqJq+0oTp+GG/nokbVhlyF1VHgSK5inXAUy0/F98gCGcr+BcFkI33C
wqEAvi9lBdt/oRA2USljKhcFfVdc8Hp0+eN/e3eoxe55E4HrWvOFhUB4pfoZhn3L1Mxxaqh3sJac
YGjfpb3vE8bSJEDAke3SfFXZ15Zd+BNNv78FTxAiEFQxABOtLbYHGfHJbZ73lY/Wcc8D4C50pgDr
mkXz1vwd1Z0wOytEkm+IvJpFGb70BMQCvaYz7TBpATfbLw6MfwKQ4AjmjF7Txom6yofuMaO5ceK9
pT0BXz94Lu0FisQUntlP6WOTfaB7lkBODf3STz4BSThWTvsaRfJ5nZausz20uKyu35ESc4vJoL6w
gr/UWVfiMBNoauE+CwNvAX25uVc+2vf0q6KnQM0zGvSjZwiO23r1+5ywabhmLuVYfu448otaICO3
rPSGsUhy1cdqDGMEYkjgsOKj3YUXDhDMI88bgicK9KKByYCM8d8JQJ9zkTC31cJLsDLiLifKKn0o
tSP6jad+0v2wcNSP3BY27QcH6OK2qSqZ0dI7Gxq+JBscExRHzX8SmKgIPXayo3APXg1QnzIPNwqB
890KYBc/P/Xh63jeEzRui3ux1jtA+vVK4g2aBXDU8k6Neas3J6tRaJux7jdUmEEBe6UiEWB9wdHb
Ik+1fhEdcyG5reXci1TgXXDqT1sLrIc82vwLxmIIMA9QSqbX3qzrbvGEuM9/f6uKk8JDOL1Ghl11
Qe0ZC9xlrLB9nm7NrdB7tPPFmyuUCzvhB8A5JwNHIqeU3zUUJfl6xj2C2ZOzNXl6ujpzrUEt9NbO
qsFKFzlpJIewIgNmwEBruqKHp+1i/USXmAuN1Zv20fY0Isya0XjCi52lDGHWkrhxuEO4MsOalaYJ
n2l+P6JyMndEYU8QH/x/ef4KepNuajQ5INh/UtnV0mbXNgfzeY92qtX9nJNNaowgfDaFnuP+WBx9
ePcIZM90wQBP6yys5SrWP/pKQU+CawxDPPZWJrJ2KkMcf4GpGRubuFmPw0l8DjaNhxrUkAyLnfHs
a4AmynmJ4iYajbvyHbeQ9KgJjWqpM5awXn1XjQLSQGzkEp0FJZZmblKtTWf/E0TG+sTPJu4mA3pt
lNOeUtDJT6/pwX4zfOYQmlhk94ay5hObhIilcMZs1Q10HXHUHde+CuHOwQUlPYjXQ4Du33l3o8kq
Z5e93TiWTm7N+pf8yuraLFFponSmLY26fJ3ryoizptId0NZ7R234MeGBqHTIcnoRdoGnZrpSdbCL
3QcdYvE2bVpcYtpp6CwUUYxAaRn/QdW2CGgj3Uz8HSXdpb/uWaNRueytd6k0Lphh8QXrD1eA+3EU
2QDMoqn5V3OD3AOEZVH7+zqKK01P8MOZGvPaYGN9gAkZ3Qr5jjc1+QmsyZ8Lm9Y8mLRnWOMTqcyH
/c7ft0Oa9HTxYXpBOj0IcCsLcxnEiavHfKh6uddNhi2dUrInSd9pCNrfbSZzoe3Qn3Kdmt3muLPo
lyt4gGHUim8lArFu8VrtOXPgm1AJP4sg1M0GukmsNUVtJP0g0iSGWqG5uChd5uFnWmqOYANQ5oE4
LO7jKDjvEYplYo3aSDXDp2C+Rtctt6BsJ9p/C+/P2haueUHKUBshmBfqqAmnAFwhOxMFF4XDMfDb
r0Yu20wmpPFDXgy9+brO4DAkoGyHi+k2ZZvlYNnM/754SiCDXtV2cxCc5VtxSPhXeoARrQfzKxyS
gOAg+OnUz/TTIG8lETcZje4PfTpoNXV95vpUWOG65qrj+W7T22Wv7Hn4mlRgDqE3udpxAwarzJeF
CPX0LAlxGVKgWgt/2nT0FNNglRd9aQ/asceVkrW8DBtjXVw0qSfrNNvgGIgbhLd6pOGOGusc/7IK
KsNwFzNlP3TF+JoQMyh5rYi6IPJMfmAtvciEtytEhkEq7I4fYHQOZ4EqYci3T6DK8aQgKgHspmN9
2UNgukb/9PRS40R9HY9ihVXSowWjjXiyEzknUeXmj41OQNc1Se+8+p/UG/oLnlQ7lNFo2Dc70tja
HOjQtbJYNsGlDlF7Qo3zUY+FMQeBGi2Gve7mLAuhq22AyeQ3x7KIZqOkeS+1AdICyL0u2RFV/QTN
gWWgZFlIAeLoO+yV6hzqM6aOXzYj6QKNPxODuFOQU5aE93oAjMnWzvbXvmzrQ9fC2AX8gxiSEdSQ
CeLkBVo1flSRuLC+nDE7+/ip9byynC+6NW2/K4/8D+m6Kcb3bQliH0pynwcYiIb95qV7b20TpixY
Nhz2Lox7Wc0Ziagb8KXSNWDLhMdmGJgeIRCsk3mcoxhIovpw3y1dcEG/hFXCCQyAKcIFLjnn8MwZ
3pQmVKvEbhHyve1J5f4uHFr/CMDGHlV4peR+2t1QPJMa2kG8X/2kVRZk7NllfPS7PAr5t4yBtyg4
ZrC3y8CPM9U2RZ+SuCmmY3CSCAIURT30+zCamS2EpV9UNIYHjLXA/dXxUhxL+hA05X9uwU1gF0XK
ndoOBPGHPMTr8/6VT+Ikj3XC/Uvc32L3Awv1qmxhKGPZ/vYvrX3FC31mNT8G/FxxPzEPr/rDMEMJ
IYmX9kRFnA3hyh91xPn2Q6o/BzCHj0eNrl33hDpypTEk1C8d1zC1Nx+iIWi4i9xW5lF6MOnKGDuR
X4KVmKGIDNl86Ux36ixe8bmQVjb7yiu5iW4FIZzaVE/ZsXiNvUn+Y7G2Orpc2VDDKQx8rig2YZMj
D9LUZ8w/0eL1t8DPnY7QThWjSXyjtkxa211855HiRlaxQ+DUwpt45kChgeWzVexZzgp+3IR98GFC
HmTxJ6ANSLv7FExO5W+BLPyELORlBt9l4RluHNGZS9ZxZFbiwulNDT3e6a2YlG7gXxrCkPZLGL8V
kgLYs6mpo9SDCcqBEywRW7nstRZaihZP59sBenKty4Debg1fQxq1b1JEGA7eGY9GPQbcgu53AEHy
AP24WUQDMPXwOdRCz3SJYE8d6tPtkF4AyNrmR/Mww4na00hy6DsCrHgs7B6A8rD1kTY4Ag20sO8s
UvUeCG9zed+XjVE88ysBb0nJh+1oi/3hghU/kdpFmc7kLPBDpZIW5j+OCMHqYb2i/ftWtA9LgCDJ
kIDbTrC4jn2Qh2+gia6itOYA+4dZPI609l81iwwoCxIW6+wezSve5u0m3AIenW2+Tu9D7riiElas
G5+7aG1DiKt5TMFc2Lc2f5qacAafZCHrwH1sYzSGWJra+wn9bboafDAJNaVSsPTLej+kHhgQTueN
Yz3/+APIIU+PgHRNGCPYtHuFmYOA02UKM2LfS/ZGL422H/zs/KC9SN6t+ZcJCvwwwAREY9f4YF4M
ldiQWDm7gwtUQeC3pOcoDoXRcNCaw3FNV3sDkzz/s/jhp2R/sgK0xw39MNs5npEHF8WDEDTXQGp4
XpSY7sdzoRe9SCJQInAatLPnByy91Y/WLoXZbyGx7FJNYu3MQ0S9X2WUl6ljzooWrKK0yJzEwGiK
eNs94TRBcyyaT2Y6Ej+zYc/hlZ//Efn7sq4Z6bc9sZOy4eWrxiBwdhJ6QRjFN7roMAGwRRO3R3QW
UAOx8LPCKwqkY269PO7Ct9OdVCdMY1qn9GEHjWgvWJ5BTqQyhvQ+oak9HmhQ7lX2Ut7nNPisGI8Y
s/j5GenXxkzOwc1dATSkySEKfeGTt4EZE+/jvcgJ+BEADLsTZ22xS6VDC89gSoo1TEGh5viHMNJe
EmsBiNhe7gZrwxwToStXGAy5zu6ohRT4J2xLwkc6lFacGxo7M7mmKQAZl9ggPo7NGHLeOf7z4R/Q
93YzrDvRDSxhY9B0ihWxukRDmty5pWnSSbKdM92hLQXK+S1pxmJdZrQftcfFcPYWIg7dO6phFw7w
xjEMXaObfHBWmZZh/5TqhmLhRCm1DyhSlrMvKkAYXj6bzDpnwxMTMbhGPpEDMByDD9BDlIp2vzfY
LOYSwA340MOmLx7b6uRJZc01PhPR0UCGyrYxBcWgwiQPqR0GkzP3XpdjF03qqrq0BOB4WuUd+QkD
wIFiraXjR8NxsSRr7nv+Xr7Ydo02VFVZnMW9cnr0j12C36fILpo3dgbd1Dn6UCbtRQ+sOieh2QNp
n6RzziilEQ0c5XvStkEL3A7AJmgfrsJZjlnYOaGlOviTnDK6MpfuyRrqirdA2R+sNl0Wq2+nXS24
UN4Yf9Qh9FyU+quPNMJ51XZQMppZWbzIyKY2E7HlWlkzQuLZTzpjh4b7NTFLDFuZXLzO2YjlVCf4
s5ktw/I5U39p46V3Cy5316u2ltrzKZV9PIdWiGx9R/vfpFV3Ab8pUffTHDOrN9mtu1FhxcS0Pd27
hvLOGnehEnOsgYO0Vh6T5SAItP9z0BuTzPhDWR+ha5EAl3XHUkxAX3ce0KMQVGJbr4NbCZ4TjBeG
hpPrxa0fKS8iPD/R2oxkpRxKYLoTNWB6Dru46fQ0ShoIJtl5Zprff8jMNb3V6xJZ/iBRfhdXCC7T
Z/ZKnYew0RitcRvrEwQhFA9dDr1ooh3ncYDyIRM8Rpk8wPod/uvFe0U4ZBq3QUOmf/ag6w37vYa6
GHDlHx0sgAUq7o84h+1Gzvt95HOPpQzfJonrcseAdFfjVIV+i2luCH345Rj5Os6Dc4qOem6nlMhL
Qz0iM3NJmFX+7eygSOziGwDT7iBzBadMKWbgLFBiJ3VkT0l4UGILjcr06Nc0vKDN0t3y+eUd3sdB
nkm+uWS7vKqZmhZwIs4L/QdwL2kv16Kx9fPFFoSMk8Qg5DYMJi045tW8eJmzI0MC04QxhUO0ZvD7
jSZWrYJTiC+M0VSB6eo8QkuLroH15ROVn6PC2Tz+lZBKTlsH4jfl77VKfeFqheSbmDk34Np/Asd1
wY+agS3HiL2Lm2a3+PfmzRRBsVlUB9UjRectLP2FEmkRExyn2gM078xEglaN/wp7pjIjL/OoS2aG
MnwxuZlDIL6munAbJJfMDnUr00BN9G259CdcbBGODBA7XNy7G/kxWSkHFKVdCbjR6Y4N4tHmECAt
yrWfbq/jsyqiXHR5Y43WnTcS5Tbr3qfUfrZd7a6ZcIglMJVs6DEbDKj4EEi1JMx8z9qt1Ae7OyNP
y3+SPEHtk5aOLXk3Iebqi3MzQqcTd9y/cR+SYX0Vs/K4sMbqJ94L96MaVlwbs/Nv1qcVrsZB/UFF
3cwZRWWKOn5jeneU84MuglaL9Aqqt5Ow0s0Vq1XjeE6vXdi+Sie8fKxyfbt/juAdbwIeK1KQa3Mb
7uNgMN1cS69XRyWFC66X/fWp3Cj1VuwqSCmY8ryZCn8Og3BYtIRO+UQz3iEoR3mertu7VeSoDFft
tqCkO6un6lCwoU1o78xrUUC8xE9C343Z7lJjLfqosl3EcMws1kcCt57ugm05Q/8BqXJNvgsTgkDt
efmN8cqRlV/Z5g0ZjVsm+4Pqk64ZRZ2VMLhrOdU8Pc27PIqozGQezBUdtLodC6xGQcs6eBp/pzkw
vzcPs6Pht/xezgakrHapzU0Kp2CBkAKDYOV6DhKsoD2AMB4TGM9N8RgyQzK5XdUshcM3LlwkCBWS
ncMgZJQtggTM7BOkSwYUpvririmTy+R7fkqkVKTvx4ntBpS8y+XgYzB0v7KvaHosq269n1nJyQZd
2oLp8T2CzugGKIIJ5LtJQsLiloULhiW/ejLCttNWGFIF4j8LIbcoth0YVvLQFqWYd5RFRdJ6sMlH
swt77erNWv+7FE4+W8RvS2zaEjHxSAKborGKf0XD+jSYOuBuuHuaXtCJYLAdYKCAUOYgQPVDXdLc
8LjwU0KiF+jwJjL54+j4fSCPFnKaJSDnYFXORab0ny7dDNdQup9+oGupUMsm8AhGXqSpRVBYZUSx
GNCZqwk9gZl7Spwz2nksXHKX0afU6mi4qsFaQw7llPS3ey242zhgDZ3tM7Ior1beX/JjxxpNKTDh
BJfyeHuASxBfO0rF3NxodBT8QcBC6rbrNd1V1KZvpljPrRedK4MXzJqYnAbC5+2zzdz5doy/7XEy
NIRmGLYTfH7eiBA0InVizg+vkqOtJYjQ+PbbeppMrvv2KjTexoz2/4khNv7MnmHUUANOxsAu+M/K
pUNT2vJ3Oqwh9i+V3Oedxy/wdeVnNSfsuhf06Rl8fF5iXZvclUAM277j6puPGDPD1f3WNkQ7i5bC
5N0ReoVyj7LeLBCh+RYYvt8DLsclhlkfGXd1twZwNRwZ6UqJ5W+ONesZCCfM6DbWEObrKrFcMZca
ncNNd/lV9+RdysBAr2Ri8s9Wz+v2+ZIREuPqAaigRIiwqVBiwblTtEidgagLnmnEJwCLN0n4BA2E
ORb5OZ5toju9r/wMSA+yzm9HcaaTTQtjGjAKHqXb/xAqTvR5zoBUdkjIq9LE2X785p7J+WuH31rh
UVd6nqduL+OAKABDZTzCHI14X+kHf7sv02ALZJqMsWIgcSIzgoVLw4mrTNmJGkZh3Sty43nUi0EU
dyNJi1QEukAeMhBVgXBpfkykOACzuJ+IELIBSq6wQlOWCUZ5EI4nMKBUlaWRb4AvgRJLYZzS+zu3
byr7F94FjvOivZn+xF2g/uq8pey6gxOPQRvqJntL0Qk3/5NWWzXLTwktFFhL2A55VISlYb4mOA6x
53YeiL17BsBIBLzRxG8C61uf/0oF3nroijJbE4QR+d7N2w9k4KL7+yzAVxXL0Q90Dwx8webvGV32
xvUbF48Uio4Z0Zkg9APTgT61e3JCOl9dmNwQ1lMo2pDaGfd0xIkpQYN9Cuglqnht69QEzIhNXXDe
o0dInlH+8z+Wxs9529vLJ+I352WX+lKBSzyhOyneRe8rc/eF6/48qep7FimLhKy6Q1vwdbttSLqd
kwke40GrOsKYaVIbx6dEMuLv5SDk7Y5lcrxZJwqxol8aMNua2GgYc/qE/vbmOa7h4Aj9i0pvPujX
GXVVZxyEvXu3FrbLTjF3DX32BVIMZMSSa1aMxYCi4s3USlSiXN09y1bYBIW+s6FAemmkm6SViU7A
gGSJUojbJDien72g9kgqIeB5lNgGVRYf1+bUPkJQqx3nAqgWTLHau0SOEqu8csJ8YffMbhEs5oMe
YlCiXobtVSE3AY6FU7Xtr/lmGqjko5LLDI8bawQzdwX2Qbpuq+73xO2LzMxmsv7jf4rdkyaE1HbL
rvN5mIEjSwJmClJheuOmnZ/cRhElQexKnC0q7JnUbyHoOk+EQcJJrJnZVWSYSwlhr8qy5sC3LvmG
JNBQMpQ2YXpcUNorSxEXPamhznAcwMg8hq5wQ6KVYzbDPRBYOYipQ5ZaHtjltMqcXDofySFZdaeT
7oVX55saCQyIMe0JQsNVsqZeTm3Hk95aXASidKSeiuEpF49KNy0uTGVxjQFeaJJPfkuC2bWfXGHt
r97I5sE2+EGCL+TFdqQr4H0OA/+JB+HBLcFz4afW39AyqsfuKhfWe34J6bZYsC4kv0D04RJYwWQh
YlJ1JuUBFjSon6Feh7ipjzxEvrrYUROA5ytq6cDDraC528OHWdleWfw3VX2dCOh7c3FW8TL1jpKB
pEwCEEUOtGq0CJMfsLMbiQN0Fe5niWMg+pcvXwTkeyQb4QUCN02OFJDHdj7gtJq6pV2zd1oCiBcq
gpIhCx+q2+vqiy+5J4ZrKGxvHOUtOcn05/siQZmBk6EkEM92lonxhaHkYfbemf9FFYLX7mtoFmC6
vfMEItW4Y5jnQ7Bdasnu7SejqBbRRMhlYR40qGAJGRPr9UHnbKZv2sPih7QMS17NNLGOZ5OUDPOd
kWVCLx4VN8T+oocRF5yF+eVc/ZZtBBr+5DXnwWZ6NQ7rlURZw3tJvzayBnH/Ns11ex0XAXv06z85
H643u79qR+apPXFaBrPoIMcxT8C+eGx/LVBqGzlZQtQbKCxrVJgaMyHvmUHGeTEkbB0nXkvROWPD
2eKYU7nX2jvvGyExrxi+CgY+zwZBoJsOec40t56RMZB/tixJ6CVjuzLuMa0nfgYPTM6aey25ZxHi
ZI2H9TK9mTKGLUapWvDdsr+jEu0QxmF7G5/oG0X7YZOyUqRhLbBv87GqsWED+pYtIqdLoc63YBE/
Aj3noFTLUVK343ziEwS6ZbobdvdkjCUpixfpcdraF2Lo5jOuVZJBZ1lz5um9FSRzSOhgaEdF2IAb
QoBLRtr9JV2YFab9Oi28p9vjuptTlEEEYWs4TzLZHg4JF3+FKzbTZN4hO5GFPXTjxYVk1+pXxuC+
Jx/ubU4Dy1C04yMJx9bH2Z/CMULGP53MI6NrnPP6FQAh16nUttV+UDFBom+nJzGRtgBIeW/SBhe7
kU4MuKnFD3BmX6gkezWTAb18ZjEgHCUVFzY4ONhYMnPe8t+kVEv60k7xt3WmtukPEuWJ5AA3WiC7
5zTU3rWfVfrNTIWus1XtbGGPU7y6v6Th8e5wxrlD4NlWbch0cPSO4/V+a94OpOgCCQ6IywGvNDOB
faBnK3rrbSAT12pbjxeEo0SNmAK1TwvYsN5Mwbdd144GMzIvGXEr24h8/ZFRgL2EwQAvbtAEoBLK
p+hRmmC25hIN+wRzyiPYhfOIFV1ZY7ofMb5X2/8aVHlN9eugY8hApUM/Cf8ovFxHddNZqes3x68v
WXiLYtx2NVstlsR21vkQ46zRM5K3GGnXvwT9fhEVfB7kc0cz6n5xVGk4xCLPVqfgEx/YzsDG6nIA
LCywhqXpZrNf4huc0AuESNNZkU5omMOb3e1Gbej9GYKxIMXG9qtZ1XfJTotL3JgPOFkN6c9f8Cq2
EvipcxxzoKqiikXcvSoZ831Ui/1/0+QHMr84MzJtxrRq//Ocf/REJgKugysFdbfqzNMo4l0sc8mX
cvMcZpdpC2fNuS53ZmEYRZlmMCymui3gTq34CQRuMEZk7oh10mWyBJbGECqodsiL6piJZ39V436S
BGvkBtO7eaVnYdyY0gsjjXE8Oy3G9XaMUfNEiKYgO8JRD9Qh2bZbB2QINQ3GRKIucxuZjcqCRv8+
u9CvvrwgAqIQ3dQTAdRFqUcNC2ohTgfaE7BihDaMC7ssYfedWc2+JLjQKW4gW5bNGcrXX4t2EVr5
UYt+GQo0hOSw7/dfcivG3QrhhbEdXYgOsyIQxE4DnCom1rOloYkOr/dmNf+xYf7fPhh/FVn5T2Wu
xbP7Wm4T38gOOVvjMd8zNURbrWicMQXWHlc+uzBoXUTtcUlMOmcXJzE0octwz3hvynkRui8dxWfB
eLWLUsROmRZ+hOOZuQSCEHzVmsCdHb4vuJ0aPRKkb2Q7672stZoPqb64YFla8ieLFLnrNyt6UI9K
Cd3SUKWgkEpZkWJzdLrDu3ATWVzjFYfXt1m5bNgEZ1qcIO94c9EMF+ut+EgOtMc1ueKftFatsE32
iXppsf6XpdxTABT3RWbKJ/thUGoTLzlctwlbzypi6XdGurBo8ex/dbS0bFuXav3s1mMLN+8a/gUQ
DarryUBWE0yqc3pZ0tSXsi73fM606Yb54p7dSEMzHzk3QKcd71YsH8z3ADXHd31RGJl9zYgfHAy/
YqpcyZq0QEZMdH7wDvgk2PvSOHEBUslKORJFFxWtdBw1a4StTMSVNx2QGYsoonLDJkB2252StBIg
+oufggDLRa9kL/y653yShLSpyD6GpMB46I1vpdogeffcQHm4wWWFCateqk1w+2cSyWRII1iDq0wp
3kjomH0K3n85hAPCcVLxh535IuRQqeJmrzgZCFxeqAGn2h/QMdioTNEaHllox/VzUAP7N5gBszfN
PwVvEsA8S6KeHkE8wwFYrrcIW5+dwr2UeKWEvkO0xxtQvH5qFCi9zZR6jse8I85rFvI1+hYZxsb2
c6CU75AxWEHSWo7VJXudvqagyfp65TGTaFWpiSFQh/JVL7JDZUQUBLwMaAv3pCKjiWBoU+VKh576
bsA+1wHNHULtSrLJF0PgY5NcL0ddx/M+xpkLLCZ/5hI7jqfWLS6IrGF7YGUfQ3RLj8CuUh/lVFz4
SttkeDtcwNhptbi+RJw19gRDvXx5D2NufGFTvZHvUV+hclCTkA+mL/LUtaCkswPaHthdIeG5HRLI
IEq0xgYurrLU0MBHCOCmfLaCbzLxU6Cl1hfCSZo4bJNGujo2bQBydAv+Q7zouHUgHjfen3x21AO1
l/vbTF6SeW/9ocfBaTW25uk6W4qsEsiqhN8H7dtYicKj1LgNZaWjj70zhaCTNENVIG4xHnIreU9D
lpgPHcN54yXlRZSkGTRoZkJ0SDDQaxEtMW/Xqkhl3Tj2ZsY0qlJ2fUn4s2oKdQ7jvkXbANObF9rc
qfn0Tp5V0Iv2thPVO4T2fobqEgPEDzyA1xiffoC9KQt65oiNxEk6uvoWTR00+/fai0kopSBta383
JF/jWYMRuy3ENO4SkFWUK0WVP/V0cKbsaYGvd+IPNrt0kicT3nH/wpBunei3ez/VOSRFettA7LXy
/iYVYbTuJeLp9K/gi3H+wolfLo0J+4sJtMuTh/s55oRPkuBjswVLE93asJNMM8FRgbgnDpeNdA7Q
CI3qdW9QRWwsY99ajv+Rzc6kv5yd+96NFxuKoHxxzOV5TVQ8FWYuLs0olcUx/kO26fd7zujDCpGu
frzOxVBdr3T+xKGqi3zIMAEqh05qMoHpjwDuczHOQZ+04ny3lYkA66eKUieSGOJZDVzhhiQ6XWaR
nQatYWA0pu87qR5fytUohpRR3aG6Lvw2rDSnFcdBW4RSgKwPfzWSEa+2qj8Jc+QD35/XuBWOUI38
VehDtww6HntA1ooHVUCQXibv2dmW3Shn+TSKP6TvSzcifNr+8KYkYgRQIhWByltrv0DNJEbPIL1k
98zsIFQTAel+7nVHQOPNPXgXnopUHy/t7TJiIpSa+O38bcxNDbS0NCUPRsGHgaM2bk0mq/uPsDvN
CrPEHQXIMJd/fTkhQNk7YyxPCNQ1GFEaQbS26outxZN14U5nP6+042yIhb5Z+/D6m582/z+WQfmr
GQjWBBJq6FryH+fKDCWqBT9AYsqoUjlYFKF9vKSRyCLw0dLCr518+ze5S4Kg+dcKxiV281c9LG81
JFeUtBzl5wXh2o8VPrWb1jfDaGOGLEU9r57TVGiwYQGTpZSzXrU8/7/pOUD7ux9FwOkpjQsKqQj/
xSZh+zHg1DqhTf6WUSUzD0mfqDa7fZultkWFbqBYdoykD9iSfEPIWc8nI1f/I/F9SixMaXF0D0ur
2NJ7yazp+aCcUqoFTCqbi/mWjVPET903++VtVCVeTjKbmP9yZBr48fxbr7ZkOc60u+2TPJFrnwwq
ypIG//hXvSaPbTQ5Jb65DD/WLTLAkAuL2jc+TJjK9hD3AJAd+crHJlVGZt8Qt3HNSdw9bmpYNSJQ
XbpnONmDP+ZdgHQ4ZJW2aoddgDxIormf1CXj76LJlYdaqOPtRDmkocJPdHytVCkX+GAAcQkSncP8
CDypOJObpNlHO7X4K4yXm02BWU09aSx9ATPEZ21c3jDcetOw51ckol/p6cgoqrV9GMFJCHtdf0Hh
3T5YtK5y0gVGY0aV4sqg1ITXe8C7M2t+BNlAp9EXqlvWos7aPhHDZa0BysKYp0AE5pXDyBSwda4T
9hEPskYWQ4IQ2L4xnHsly1bENakzzQg7OI4qqvdPTK7ypbrh7b5UxlIedFfZqfeZWFwRwXdg5ad1
4LOdgU3v/3B49ShkxzPsYQImyLtdhzXp/2wBE3pnoxZiBo9VitlYS0pzmxqtsF180HljDa144W7t
UbVs8DKny4xum4jkL+4Wders4NK61EFQh4XaVb6cYBsZJE06hM4OlMKROtpp1unTWKNSTVp0HXw4
a0bWQ/wnOHiSGt6UKpLnDrJiSv1/MBSvxS0evDJRBrQZRAUgxCGSuSbb++Ytqh1IETP87B+I4CcS
gAJch9E7Vcw1yNTh44EkYoRA/SYbiSEPg5VSLRZSORnrtcAZC3wUNAdiZ80bq3NXUcyFa8Zjc3g4
f8ZR2Rev/SqRHJkCDcfkxpk6hufNe6ypwe7Lf2SyDWGyysBOYNH67trI3gjWhncjiO1HtJdO1uiR
3D5GvURt1PkDtf/ekOvydwPjUq9icULA7MmT8CzRxjLts1kK9vY/SVdYlHf20fCyOycQR1xAe+S+
PjobK0/e+oIKmbF0HWfUtjKx1TE35kKLZb4UcVxrQvwh9lCEJOfM8OLiNg2x8NSNhg87IkneuS7l
s26G32tk/1tRqnRck/bWD8GMhjRrJjwCPaZEWiCCCiKpqJkRISaUh/kvRVdWn7aAFmYofLZ6TkjV
zxuHC2wNVRSfW804Almejh9JghIHqhxaYOnN6WFa1nbzDi6CHK3GcAXWc0fB68XCkN/QeZpwT8Db
ltiLrKrZ2DSrlal/EopYmH97gApLPaK7A7ksrNt2l15s9lGNF1Vmt4eaKPj4jItIzox8CnYhi1U7
oCza2Sboeam0NuhP6UZ6ymMGKxFbpHw1sWmFAFiuHEnv3/CmauNbb9RZm9ksnBoijC0xS9szEA9P
4Zo6lL7dpcukfBJndmyHrc4SGlx3HIPRtzwFXmfjvDQYJR9GYO8dtWE+7suAUgn6W5DQ4WWYxS4F
0d3MTPEUqtxm3PAOzUqBc//Uftkox8ZAOw004N7e0BaVWIdZJEvwqwY34C/JBdfkfszofvUJ8hVC
YSVIsuDY0LOYfKlPUrCs8pvV39pK4ug11YYB1gDCdgie6LBOeh9Lzz0P19iD/b/de/mxFYTNNbdz
agjh2PjAQfqCzCrFtjBQOMsr3kEmfgPJq4HOJo3eWneuh/NaEDeZrgIkG/fYrILHKnZjsdIdNbzs
Y6sbiFYdxN/r8w/hE744a+NT4yq0i9/6CSrIyUG4U++c7xi5Vbh/2GtZattN7wEag2UsVTEDHRBq
yvb/AB5pcl6QHJIdXlLcgIj6H3SwIwopTthtg8NwHQmtAI3xUFt3iWkqUavwQohWGlIO+DnaYxIw
rAdHXM6QIlzOFxnWkqgXX/DBIYt/rjt2yPSzQh1+KmKhjuZVGBR5K8XJmnBctpPobYo6P45SR5S2
6VrH9NyDNEvbWUlGnSXxA4/QeqnwostkJxC8jOMfjDH3P8ahl5koTfHTrkiuM4x4YoGyvggwmLtS
UtyO9lHfaTIlS1Va2iuEhdZ5YOCfWmUb9BeR8dzaadntaFZaOc9836NEcKWQUdLZUiOS0ZXqpI2T
Nkwk1Vi8YdcLnTZde5vQQUsC0Q8D7NKVrLEUAvdR635gzMerCbGNr+dtvvADZtUvOwzgYl+PMyuc
8O0vPGrqrSz9gRzHzMbOKuELdlhwsuFRW5dlXcJcc9cFxKgAoMJ/ScqtvSi1A/TrDBUv0D2lplOi
OMdtFBd7YVYcxERM6oGuh7qpiQqoAbCBF5TO0oZllAvlysy5q5hMPx7+bRTDSiuI6zrnnjBs2tCj
kBjBVcZ4ucGIAh+rxdShtHfKWnzQgbAOw9pzFG1FUdM6PJia2dtddYYokQ9cjC87I5bdPTnqGbyF
XYXC4waLIu0hRnzIVm6lsfudjUXRe0dDXkIRapoNqjsgiDj9T40ezxbOVp8vth1eaZZwUh/nnfPq
YQuMnZOH6Ip1bFi4EQK32qlj2aao2s3gu2GKopKiNLVaNEA0FghxNn1ZuO7yCDPWp9CwOwHwHCMK
uIuF4pcNxMdbBGkyneBr+dIcN+efG3lN1Emw1mln65AaGx2rGeKLZuRqwLGNPABChqH3COTSKs38
z1bxlO4zc0K3OrKW/TqtslG+9LDZiHy3P5Hls9JF9NbzbESaDNZjqrwrhMKRewMwvuh5N9NVcKOp
KPgwKN3WChbjLZtwsNHHZQRVva3LkzY4SsAlCq0YEvRQoitHLpbrmrCFlu9iSxRHR4hXHTdUUadX
hP7helcKMA8qVDF4Gdgf6eYWq38Rwl4VdcuO7uByVrahYVX7KiBqvUVx74WVBbmGacUTOTnq2Adi
1x1o94VV6OmE6c8I3h1T1aNASl6HZU7KLAbNtBIQbEcwLrFG6ZFYmA9A/rvDBiYGBQf+zUqiIqqX
CVihljBjKxO3dE6G/fbVzKLFvI3E21RMyfTl1QZDPVm8YsqPJ59ISSp3WuU8YAPcckCEbHQtxTN7
SoWq7UFgJt0L4z+Ey0UmU0a0Ed/+fMtfusiDbJf0ShjEv1Wsj2BxD+d3PVuePowZg2rjfRu+prDd
lJ0lspQMtzKut9FN9DDrCGtBm/kaoPoKpwfPoGQ6862N9jlXkx7GaSXw7UKZ9DHArVbfbta9XJQr
lqoWb8MWtUKYOTjSibbzUhDFCigOvpdns8/uP0PEcqEVoCh+fQaeIpvYmDP/o+o/WATMETjNZQ6l
9BxnZBZNkbvmF+DGN/Wo983Xhv5LP/rQaU5nqJo5PvPXXAIeQzFWQm8thpwQHtk59Xl8XyrCkLyB
mfU8vX3TvLMMgDcJeVkYMD1m7XUGQDdINnGxgFomfA1kIF2++hIqZkdQXYiu7IXifCMF8XUAjGOz
fp1IhIvh9PzYTReyblDkLO0bfhks7Q/58jktuMwuQTlQeY/CtS1mid57pom3auNLN1MOBnBK6k8K
tFPmjoAs1k/aSw2j5Txx+t2DMdzv24eHCw66VPvdgcUjKz2/TrQKbIB9K8ucwZKP7WTJbHlezRkW
Cw8B47EpAX3e1zOT6T8KsQjbxVOuMjVE+OxsG2oWSOhnQS62fz3d6CJ58PHxpJs/s5LYz6mcVJgD
8ka+iKArx2rvYYAxnrLtYRM0UEvvvxDvQXN9X3wSdwOo2Al93sSYNzqR4zDlwzSYBDcKoLags0R0
zVnxdINzLgK1efFFu/pPs0t8u+gvD27jfPU3Tp3M7wWTvtwhZHq/vVZA3lbBtBLoWa2qo04HNdtI
uVCwUC4MiUb7Vru3SkPcTmU9RSDle4h7YZccZnW6zryiBuqUoGHAjk4yDCuZq0d+9fgCR4/2xaxx
E6Q1DzgrJggWVCr008HkbN4r9wD8iPqrTf98TWJPfJ9uDzXG3c2+OTK9nENVOg1KWExnpb8M9HcF
3kL2Ek/SV3rNA08CGKdv8Y86P8kuoBgu6s/0vU9X2JOVTSUpnCJZrGxk1jVKu2Ky7wKBLLK6n1sd
o/iAw5URlLK29Vsuu0mmOVF7EgUxNOR9PRwC/gxon4lLFTvSceoendO/dydkQlQ/Puo/H6MC78DY
pBU74lsBBOCEPJYMn6UUjPolNQ2FA6zOxKYe55nDc+mE7drtjDJ7gygo5oCF3dVwqgVeLqRU2Khr
h15VT6kvUVf72K34j7N9s1h/0Z95UPj/zPmNrdR2W02BYNHxtjaPVne1sObAcDwNUfN3XXDvL7jO
ghlGaHG4SgaTtQ1kyZ+hj8/bP1ONDMa/dQ/mq+vUpEIPz/JSIYdDUpTbenGtSV14amAOTPuLbI+f
2N2eGs5fc0Ux7ixWoNT6RiLf0PQHVcVl7SruRZ5egZCf9NyDAXEGN/XaS6zGWVG82Xw+HXYNERzf
86gzMFArWiuvLTdEgG3FzNZivW41XP01ktkK9z8E92RS3q+gWsW04GD28iryW8kqEAd6TcDFV3Y+
goL0GKn3xq4z+Ucg8a9nb40SObN7Aikjvj5mHRxgmpfUvt8MpdWCGtK8GiRTZXngZ1NCxdIhttcf
Qen7pMHTR4oJRYuHdNIKSaClbmb+sLhCvVVb1XGijditf9hJrykHdrww88w2pn4E8HNs+OAoQGg1
2gQYrWE9HU/Q90US8kMxEuk55SH8TrZIgv532Khr4j5Av1EuNhapuq//SKhBfuNcIxEwo9Jipb2d
v4qVyf/QY0+fsDnj1ZALd46zTF+uZl2rDXHIDWLPM+bESeeg3j8crYFEvyxVRSz4hqiE2bpU/uLm
inrKmGMBNgYhCdITGyVlz3gchkgrMN++Tl0e5xU4ukQ/7z+HQbKLlYV4rNo50zA46cEg8O/CIkvT
DEABkWxyvP3iGmy9qXhxp/GPO+E/eaelfJw/yGma5v8SJQqxKIms0YQd36yQC67y4GIc1m1tA6BB
MjThFZGLYIfCXR0ZuOxxPXQnm9QE64Z6k+tbUhQn8OVMbJwiOpkBoJSijTVnHbM5v3SllwrrEY87
LaOAbR3NIlWhW77xm2egLFKZfoSuhqzeQzA5ZkpmoT0S9E0s3xvLUMfBBHp6sCiGdIrOgx738SVA
5LM4qNitZ9eBdfz5eLMp+7Qa5qhQcbMgZstwD/spPcySL/pHwYXOyWWVh9ae5TspJkhI94yDHiKb
2wXqj64AE0LgiU5lzBOD6tX7S4sNyyYWSVljN5k+2cFNDHTy/Witx8DFXi7aaUtD9gl11yroD68V
MbT/xutMDR8tvBoHsGk/0nDdQYC5K+T4v8VoaBvl9ImIT3NIGjWlAVTwAsUD0HSNef6NCiOv2wLS
wLgquoTZNZgblcGdcpdVd1Wx8RRBJ97FR/ZF0a/29UZQ8uIY69ZwcqYtFJ3U9YvVsb+Ns7oZFa2B
6vQN8+U3gU6uxVXZmTZyKapC/yJT7YwCkL1OxRstYJsIAfdstg9tnrs89pzNM9Y2UdoplMNnEsuA
Byet0Qodf7sEcZu6M97c9tk965Ic/df0V7hF4nuHiQOIQrjESNGWp143jAkDUtg/gScB4L1jSYIx
iRpVPzt3HbDDHTh8widZPcBSJkxKb/EUkpY0rVPTc58weGxp0hpdWMZytmlpL5V3Z59ZQBfzAnN6
qJc7UFHBUInDNYh1Jts0/DCRCPxqZfRXGtfGrl44MsgXJSMtSlpNccUXn+Icg7SnJD7ixBlfEn7g
sv3siaxoxMTiG9VGQljC25BV/TwfsdOJG6zRaWiKo7KPstwnRIEhPjnjl7lwMBeM59OcXa5SyQQt
0nP2ZWjxfzQAOXnhhmNmjfRV+YS2iErYxLSYvZ6C8EzdM8adTcDfUEBJLIjFmh2N6QMlQQIlLvpO
HFu+shAyYmE86r5kVCbPSUyUuAkWMNSpsaPIZYLOaXcMy/J1aasPL1NDmUvWHNTJZZL76mxKlG5Q
/KVdYxFIpo709XzTagoD4uVUy7CXEGv85NZ5xt+yEmQTDvgM2axrHZMgWY2WNZXMogJYOSFWcFJR
J67/ZgDiCNrHVxIVbxzAuvImcNKrEDLB3tR2FJ6OCGk3JAP7g30vHeRVrsll50zREeLPw9Pg4cCL
65oRsry0HnXGoPLiQedEzMPC4sG36lTvWfzC1oPJxkNLHC/+w/DE7NjIu+m9qLDQGjR2NBu2n4Yl
h7piNy+pYasH+4I48vn+ci94Oe6wLt+3+FXP7+GIG7krEUP8IfQUal4wGS+/pUTpRi8QpVgnrdt8
3sH1iFwk6ulJLx0IhNnjJHbuU7ZE5O7AGCj0/sdA3frSKQKQbebx3GTWHxQW8bjstxhC4ix+JGSt
/ZfMRPEj0MViuT3G/S75ETUBz1Uf0dQ0qDUUzORQTmfVBaB7DvecNPds0PCrEGJfgCKHE8MCJnbL
jD42e5QO8YsET3M1hafp8PtHSeuFxmT5XoN/pTm50YP9e1V3q7jxple/OUOaLiQd6kej7C5ZdxHD
ExNNEkWS8kixxETy9LVN6v/if27EvLEcAwmv4yp5w7lm48kdzUWe1WXy9cDv+DpMZqL40QNP3Ufv
Jd5/N0ZyuMjK2wTWJLWvskk0W6IQ9JB3yGvPm9iWHNf75W2KC2D4KK7wJj1uOEe+XcFUb3o0NFZQ
Qdjd6an6hDJvQWDOdhf0TXcalSxl7B80qJ1Nv3lMxzPQfpN8ExNAmUrhtBzNK/QBjqjlA33ZY501
LC+Jwz/tIfdt2cmgaaXfkClsCWbHhsOUZB8E3NYmLvwBs5BL3t3QDGvmW+fHLK4FxZ3iT81y/eLW
53JWxFL0uazkkc2s3aau/flZsFDkAllQ573mFnkQes+q6KokQsJ60lESAYP5bcrkIWR5F9o1Jxht
cA6CMkKhcet6sM/Vhsz0ol9cD/qcg0Zk1drfVjMzLnstBaz4NgctlVVC6ru2deEl246Qdf/KO1wE
JdoxPIMKsijFp5FH1JCvTQnMBaU5URVRZpKQS7DP1pif23qnSpTpng4bvDF6uNsqlbPJZ/jCFDa5
hA06Tj5eO1AvPEYMk1q5d0oeTPs1wN+VBUFHnV1mzzLqT2dkFLDcg3Vy7V+Fe8cuWuZLSld0yLlx
0O+Z+7TzIVn1CiQHCO7PgtDxt4blzqJJrz1WV/++iPK9IzCMlhkrEHQSYjY2XdrJm7+65uBJDsGJ
bLNt1gwvgUNu439+sIw48jvZhYlrbmzi6+VSdCb98RgSybNrzDJFphqj13z653i456IF0B+kvVTC
yALrLiHGH9Ls94gYKlb6Rv6X/zZPN/YSpWHIEu8b2X+D5OZGAPR4KpwNMjnTrJAct7DI/uNjF72m
mbcXOPVxxpbQAVgwuRAbAK9VeVNmv6fNsHMP/zuAmnMvQoRp5x3T1fdUurSLyhoR9f9LIbcodn6V
BbOxdTHrcn0m9Tf3sV/uZMNL+Mk5/Hl075whE8zOzlxaU/ReDSTuGZqBS6Epf0MlQaM7a6qtx4fo
qiEhXq33Sxif/4jvnG1lAmWLXuLFEWacWNJbzQ9DhsDsTx3t1Rj1QcHiBQrXglMxdhoFj1z85SFC
eLmnoZyjVIG1LGuV+teqc1h3dimBx0sy/RZexDA0xFb3V8zr91ABynCppqZsCYAL++DzlfmgEWkG
E2rIE+XTzH+0ki6bmHgw//cepypfS+Uoo7Tcxr6wlnUBQabpjYJv1B2ATMdDt2h/nPztqsLztFP/
4K/i3pueY22kJJoQNqvsodqu83TVPZD0F0UXEFn2JfS8M/ZWOszYzOVXB/S7k9eMpfSMwDtgQbPo
7PUOeGfwFy/+7x282RC5KAsXjWdRbwSWy8R03w3/Ruvn45OFKru8+/AKQ7KhWAFeNIqd74lXsveW
CPFTjlVe1qr3+W0xJRoKgKockB6gYIil31cPKXEEFTZ+XAIqVP53g6xdvNm3sHvKhEbQ4JB2aAJ5
ZQKZ43f4uUSHBFr4LUrUeABTDZHi7nuJqC0/P3XLFM0R+HkcI13uKYP0QoLUFo2iC4hyTn8PrNpJ
Px833hFqFoNRm3+GQ9kcnPjUCod6IYnOhYL25aBbvFTjWj1rnWACsf2SxSvbm3ItFhu5wkTDn9a3
Sg4XzoOv7cbnn47Hs/5O51zo16D/Na8p/1J54J7jZJv1aI4HnmwWS4S2XuqghZgvrthT9XFf05XJ
P7p35M5ggk5czHKwW3L/O3tPW4unRynoHFI8nJkNiqtbdHZzZV1cMUWjKOQq1G91swA1o5XMlCRE
KqPK4zkbRJQy8e0BJIC2VLVxAohvH+yMKSNcqSQu7Qwq5ZODr3aWvMbQfZq9fKI1Ia9QUtesBhuH
kqjOUwSZapQ0nzTLMUgDoWtrRKFX4OEU0uvKErksCyNRNZVRJF6JtraI52FwpTX+gRE0Yj5U/Jzq
dm2FRQ6i4qPOPifgvysXyMzuSo+wmxivVLA5v6Qo7zoMXyNNvMmudRN5sGpnpKsXsEcueqUeG0vB
LHcpy/R4SCxnkVt/OKvM+X2WN17MkE74NDL2BgPz8fMlyAngs1hBj12uwrRuIZoFRESFesNZGsb6
uw/fkxTl6twZI13TrzLLw7pJ8malb3zfXinhI79tmekRgTkS+L3ahu5G/9okMXkO1yUkbdB/09Zf
jWIH3WTqm8ae+oyq3AZzniS9H2ZKexNkNmCK/6OcYcIcPnl4UfPqP6RcAPiFooXVy3crlIgvPP/N
J6mPQnq2XW8SRaJoEm1qKVLj2WCzXywkcH7H3MKmLCwaDLFh34e9RpoYNARS83ILH4Ldzdy0UyPe
ueo/SwSkZbB0bjbife11h9XvufqxuzYYhAv2IKSPvwSlePtGkbG8GfpvANXL4gkZWTSZrC/MQyWG
7C8AnP59VYqZxShOiWlUAXh+tWq9u5PhM7cO0yP8hjjrLbpEDzQUsUXeQJWfb60wnZO5U7VXHByD
bThPp1oip9utQtfVoThCH1ZFBNqoj+AVC4fDKKLfsLIOlfmm8KD29rB/ZqXEw0wob43pncKnDj/y
lbQNsntorPbY4VyPLHARM88UNmREivWZPNPO2BSW0kDhe9429W6LdNMevPDT1XCxhNUCM+0bXoaC
UKBAM9ZbGsB3TyZMFe/DeGQrlTnF4TXPebA1tCHM+qIeVrayk43tcMfFluSl1vPL7OQH0+75KUu6
xjQYTtktCufCYTabVMomUk7XxpMSwg31sgYaKjUCdDk+LoTRfFaMf5eLXHSMh87wNrB2Dd6CO9Ix
jenvGrqhxe9R1wBDE0JzSR+iyr1WZmVz9Rn8cgYiNAdKu+gVeIES2JZwWfIalr4qjyC1i9FCfcRK
9j2QxrQFNYq4Qe8F60BAjYfGRfBEI8UhU2T4Y3SIudBTgqLFDrZN+d/UnNZ0ZLilhCkstMFAcdlH
KQrNUbF0KUFTLsc7eBOfxJgIJs7eZHaLGJ73Neq/FRtn2zU3YBqb3xcQomBSJ0dl1VnZSEbHFX4A
5Dwne2wkHm+E1Zod4ouVTaMEUfDU8oTpS7V9NA6SDpeUaXipbUXkjGKsaPX91VTsXOeyC4KAeTYU
dcRwO8VgoXW0M9wvVO3nbIGlyd7M888wZXKvjDZX0uWcr4obwdlvpB61UPeRELkSi/A5Kqq+Z1GV
grlrKECWh0Ok4gXK164nmYBtgoDh0rJ1W746scwPterqSyn0vZRcMHu+rmm+Nkqj2OBejfErNDeG
suh475v0j7PDxBRw32uE32RT2zu3aa3wSDHcRVNs2bk4WPlbxv5wVNF4nNDlUYyz7aFytH3UH7Jp
/XPui3q9PsXpNuQekh+tnqIjvZWUApVBczlLRLUktEXw7QGBQ9xTPAswUO6wBNU4smG3jJXtzRP8
98AoohDV9ATQGlPXSrpxEcvI8Xc5tNsFVsz4c4Hd4i8RCupNhUvvSzYwmKVBg7nGnES4NiF1YULg
DkGDCa5yJulBJca/KeEfDqqsobitaGmKhiHm6muum3EurJYLFZyJVWgBo6cRcYGhxqcehzc5FHaO
t4sdB651IX1DNb65E1F/wQlaD44iceDE0xvN9B7ZgHQwtqZls0B5cdFHLRoCsY1mhggV6znNglWR
RLJ0PWQED7OfTmt8wo0WKgaQmr0N7zrG8Tcf0YJDWJxiuth8rnRZ7PxQPtMj6/krCYhPPXcD6OYL
u6Tx/i9nACOXyjZQ0qLsn/EOtzP8yqyEin0D5h5/z0Qx2sEy4RVHFpr+pnaKo/VcnJ4f7Cr+1mfn
iYH5/GASAyiRLxc/f6P8V9h5Ty7+FwJPtlhJFaNI5gijc30wDKcpOeCIZ1/1hk/sAOdz8/2ncNS+
SI3jzrhza2RpA0IKhEpeQceEdzm71ygD2tlcXzLH8TDHY9b1lcnziNPCejFhqclygWl2619ftHX2
kbisxEZc2c2tT1voU1vGab4rxuoswUnjZM2lsSamVeHCNGESgQa6H4JuWzQP9nPYr5GlddWJmiUH
URYdB2iYpT/kEghlLJ3yOfqtlvvBOXiO5bXiTDDrSolXFDGOwnkOXBQcbRXzsn7oDLtOpcKKb3O4
aY20IWaoE5PdkasrhgkMtHcf7/EYhnoJe5Nfo2kpQyggy2FwWpyAkfMN9mGev+pRAiEON+juAWmM
LNQed7BZNSPzUYCPAtpnG/DtMi6KtH7/1bAxLiGh+mrQnAlEZvf4qHQmVdqDxF8SEXo5tCyfI2aa
1XktwpRFyJci2KpaLrnYJXSg7bsSU3ETiSETi9PGeyinMkzChic+ygPQbrMKQ2A9T5bWP8zglgC5
OucF7nzBGH3SfSEuHbdE9EVSKflOJwMzC5B3fFESapgBmoi7oLvGwKEtQLHGYWlSadnKH+YEwv1T
6jcjJhcdcVGYVo4x6NpYKSMhqCdR2Ee84eWOWJPpHGrU10d35mIupRzl2RGGEqNxS+I6HO3/LFTA
kQLTileh9MqwXiLqEYsEyUggH1er4nogfGH+O5ohOIBLB4aCVIvVpsnEdxWpxhpt8eERUDIU5Ozr
EV3xMkRPeBdA5wkRGbPe01R5sobwOR+4O2xBF+W3liz7T38wdBNDNyVqu6QshhwkCqBczw77DiVo
Oc1gpQimfFqqSaD+sFmFLTbt38NhA8gytM0VS4XpvQ4heuZFEmNGGnotyRWQ3yLwBfY5K7rrq7DL
ESbXN0Pil5qwanWZsNmOrveWRJxn+aO1AtvH8cPV157i/r35wFqzxMoVpqZcNVkfgOGqaE6elKqy
6YJRpHrONV79+uN0i7OvZQ32vUXrdKSXuObk3tLyUBSC8FDj6cT2MY08nx45tGTyB0Xa2G+0xqid
ZpTstTa55uqi060ihau+Z7s3RCcCL2R/VcHhRK1hHN0DNb6kFOB/zsIIO9NHBlc/I7I6lajPEXIR
PKShe6Ch+pvQfoD+CVVQUdhwJd+FGRYn4Ri8cBGiusrT+8hXt2hhvyAiOp3QUHRDUWRR+gj8YK2e
rW8TnNlnvv8KBkSxgZZDRyu6/2B1BDST7p9nIMO2ZqjyrNeFbLLf/9PW2w2kgLK2lFpfJElqCZnr
b5vWOdt3EZfJHlI6xbE/4qTuaRLgHYNOGN7IxJZBLKfUMTqHgrOypACHx56EkMJmE43YhiTXM6DM
gPnHRHumj0FKOcp3FU2kOHBF7I+PEqM9vSduDNfTwikroLgOEDTxrVrv3R8qx2bgV6G16cNmFs8U
2RWCMtAMOe4oojTDca8Sbx5R68M3CFikCeMQgkfwqqUDIk9GtYphNRcinYsAWQoJD9ExNnanDWJl
3Q9AXbZ38lQv0Sord+TR/Gn45w7+VYM7Vk0vRfwz/i/Qu2IrKkwUzoj7dICFCycQFeCG/vS5yrPm
q8il56BnaJzTZ4SZ+F9gMp0XwX5ktuMzhnoEr5b5niiSiL38D9ezaaTZgnk0zs1a4jncPkvtrXG6
EiMFLT5gL2OtVNFMvuvREweD6MN/Rk9l5fKFODox8JRi84AvGUdshXhv1N32XVOrvkfn45ZWfUOh
B9+DNQI7HRT7Y4U6Jwo5Rbt9sxZKIZrMxZHccnDvPE3ykp0KAjDyjOVwvK6QOfvrVOAJzjReOXtm
iuwynBjsxVa816njR949h0Ytay43+7gKaS3bWyseGd+gz8c57CqK/ACwC9bxC39+CvQwfKE4jqd6
lrv5XfoFvryMEBjmpVgG/ANbxkUm7KUIyH2VrmINvjtjsM50w05XuTuyKwlda/8DG7k3DFMjjN6o
khuuAqN8ZZyShtnSsXJzXiJoAb3fo3hGlWzXIrJ3aDShvXIyfewvi0Iuqmxcrl11dr2gthSZfftJ
KtPKfcYiZE6K3LNJIsnN7qe531Z+UrGeTQo2bAC56pXZzmp04uJb0E75i+cvz9tikH0hsQUjCxyN
+n3uhqpwtpeTs9oi7iPuTS8VU1obqgGdknzHSJrF9onWc502shyZ8dECFMooaluwua9lQIs1YRdL
xayAFKEvOQsUY+1Jh+HhSXEyXHOnEl0oABon17quxRDL20xJS79Cz9Nm6YT9Nw9TKGSLLsgSU7BB
4z6osAXLJNNV0ZG9x0gTX8e5sNY/+LkGBif1A8u40jaB/j58g0Xo0wsUgjjQXEdD38SahcHMljog
83jwHdEGWh7O8xNOdVvPez35QxussScONvzzjF6+akPsUapwcTpKYca0r6TSK9W/jDUzUh5Mmdub
0N+HMEc4+j3RPfBMKqOybjloeDYznahingv6WBFVTMal/Prssnf6DzZBlTmgLDCxaJN4RDoc3QHy
q9n5tDlmJWZohtSdULWObDpq9COkBAdvDCrNPnFeMXYvD7B8QFuhDi/4l6KXoMUzmmBNPjULF957
xDUbKgqb1gIiTBesJ6cKME0rbS0aUSw+usj8uq6FVYBqpA2vbHPCV5kq+JiJh4OlheAaJFHJdIPF
VFOk531/1xIcTbY1HuLvqHEDWESnmbBkBf1x/yjGzYio1jQmYlCm8ANomFz+K6crexDYuFtPj53P
tf1Ool8Uccg4YMb5KM0sDrfG258en01pY8UU8xJY3L9hFoLJIpgyKXz+Xv1A/W1PK21t+zMZNu0s
IEpBIODgfvHZhaAkQltaD5gKiFaQMq5q/d58TKRQZSvUjKo5+b7IatRyIBbGND3MK4EHvl4K6Bbx
whqC4Wk7aF8xc1s+u6J/l0fhwQ39kqtth3IUoIvR32fWiIT822GDw34RRCXm+p3tLjEHDCU+yE8D
85xj7Vs80B6ley8+K/UTajScOKjGOmxdllwHOKJIUO0iKN8EH6/snpPiZk21SjOcW7gQwrQR3i8o
pqlv7bna72+GoJSuA/NpDz/Yl8FyOcIDAgT4OaF4k0TTuqWs+AD4Z6annxlqSRiC6nCc/u5pkbuL
4/sVYm/b9guX6b1JiND4v6NofZjWCmTcKJhaeq6mzsIapY/mM44+QTaJGHmjc2VP1V4JsMQbQvaA
wM/IgaCI3UkRhCEFMwKeYZN7PVf59bGdpA8xZOQV+ZgrV1BK+yXX70we/1iNncULcN8ZH3iBfRrk
xuBIAR3V+XC5/vnTcnBn5/oe/RwtjLur9lfI+RKSEVzvKepVeSV8YHB2IjUNlWaUEDxZppmSMuDy
/gNcXhYcGjp5rC2wjpML6o5vVUwmw+MpL4qpVSdU6uXMj6AYT8id+6bp12CrzgKcErDZsvmp9g4p
rWajrcAsUZUoW/seNhIBPVtHddFIOSBNEQbvFbFC2PT80/0/Tvy7G3ll379+tq7XIq9yirkSufkt
lxUmm168lq8k3CkZNw2tW2t7SVnfOh7A9HiyzhE9mzS0HfkSnyJESKd5WDdn91XMt4rB1ewt0IlC
FZgLH64AlI84edCUnmnbWdOPfqL8rU1sVnsg9OB8PtyWiVWDGwZPmLQV+YcN2ROhSMJj7GhdJlDt
scYUKf4fUDZnKaEeygTQMxpq00WXtQjqqfkz+ro0ejG3IAT8tOA+qFq/AzvcGz5YH1HLMCQ0Tz8Q
A18kRMA79HO58Cosklu5qYhGdLGqqVH0P2fHBlohkmMd6LJhXB5cZis8o5TU9TBWDDxh2kZomC2L
vRDlZ8x0Uyfq603VWVyc2q5CctdCBdTG4ebPfJaCWmEeyfB1Vmxk90QF9uXo/tLeNTi2GBLd2crG
+1MubgYIfAi2WV/6BtECWKZFj05Z4BmDGlIQo9e2ZHwXLAgcEq3dFziSyRRXTIwqKykk+2gurMRV
X5UA46Nknc/X7PZSeyacXh2ONCPfPHGDHqngnVuBFn6RD9vPtzf+1VePHq5Jhbx1dBSG2xodRgs3
3f1IyqjfYr3mSUwPKSbLdoaco7YlTjWtyaevC7Mm5/EQg8pS6y15ALwTRmoVFgkAqRSDkTcl3YRd
vKxheOvnZftWCGE5hcKzl9hlJzTJ2RgpBkDtVdnT6CNnAqCKICJSPy7Y4Xlsr/PXZfa1k+0qHAq9
R2QiaH8lonD+S0EwoiDlT9lQmNsBCjaHJjSz1T/JO6rQ8OA//xaAeNQhfR5WZPQJDaTXUw/g1qrP
s9tNdM9NU6WTqdmSBdhzhyCG9ifsamcXo4iOW0sJP5xHMCbl4fXVnotwYUAbN/hghSz73G39b1ZI
xX1HncgwfyydsAAv40Yb9RSzPcUOvVClqxY+kB5WY5iQk+a+GOl6Q236Bb968MpdXcP+4L5NEo//
H7mRAjg7z/tYwX0t7y3PattdoVZU/jm45XCR/GcRwHncCtj+PihlmVyD5uG+xEjTaTCQy/rFgF9V
g1d458FZNNTQsOYtEE+KNVC2CqNwl0E/X+qoCM9F95oNUssHS+bZJeGZqypDKB0fA0Xs0X3dYQG+
sFyW4+t3Tf4eotagIBfX95LctvKHH02Phz4Nx3rfMFshSxeWwCBM8t8IeePIrIPVAHwhcZlaPDsJ
Ac8qOmnHD9LB4g07x2VkJCqisG57hnLPvdS8s55EGNu8C+iq1XcCis/sFovbq3I1nXiOU8IZkb1G
86XALA5Tv9jUwOzw8XMQUvt5OBzumfJiMcnXGFW4lohOLw2CJsAGNqregEr1l/n7NrnX8p+35uUO
tiCqXjIjVKypz/XfXLV39ndqrFdW/B9nQJPnu16zdDLy2JaT1O7t9qBNL87mht2Lux5E+bw2tXN0
QEeU2977hjdzrV533fkU0E6GlDhyaFHAfwv+9mDqTrTLftw7oOJvZrx13HNTCrSxiO9mHDfga176
7zsXS97Bd63IkwN/9tvBvbdFwUXLgF43loAS3F26LocVB1T6hV/sd3iQnsZXyH6ruVBsBnWJiVXr
vgRxSac3NgIuJkPuWQIGv8AYtuE4kvafv+dX3oAGjmTKumSHlkkggOLyTrQB1cTo4XyOKthJOped
XuabI0yPJmtphoQ+HCKNdSQ4fpQlEvhoPt1O7+GVatL3YCeAT1ZDxObv61XvgUf2dlKkyJkerrs7
jnIDgEXazOTCR7EJ5Zp/l2C+kB42Tjp/q6wEusBptRiEAJigw+upd5T483gNbjWpxO7HQxq7kgtt
JGl64j7EPQJzy5FClmp8RslqU54G13qxpvZYCXLpO5HTvmSrjG8lgF3IThfbpO/of/68Gdp31ANl
7Q74s53F1Bfb3A34g0UpTCUvFMKvXG8No5D8c+Sjzdcczt3a/YN7oAWN65WXq3BEraDCt4LbKn+5
xp3YHPyg3P5gCnHCsBbC1sAstoGDbnCNQY/nNZS2kiBXnd1jrh4O1PZ2XQvR5ItweYvkUqxR9daJ
TJOlJrdr+5Pu4W5zflxafcBDmcICqMMB8hqqoRtJHcLVotonkkM7tVM1NzBtcSIfbDwb5sEGb7JW
zUKX0v/qm49W1j7TNAt5ritGGN+HT22Xjw35/wdYDeSvsYMvhER+mGnB4cCEEnFzHFjMDjvCcqmT
CgvkVRdZKW+OmvDQivLanSXvBuCO98t7gKXJbkaUDTeRgiYwnb2zdjruupbSFBtZliO7HO0POY/d
K0EqJMKprI06JprpCcubKRcBA3iwmuGUew7/KQNqJNSbm9RNcORCezOkdgDw8MpBL3FHfhMJiZI7
UJZkHjnGn71QBsAbsJtCXU6iDRgct8enCIK8xwxGnVwI/azUh2oSU4P/f6n80S2O9F0OcJBXMOEn
dA4yrk3Rhw8AqPrRP4n+vLdJvHmOkQBAKuKgRwBHp43FgBSreYjWnrZsO8zERlQjMlQtJwB5Lr6o
iCnVoQ7oxCX7s+HoArDtk/McU8YOqBAOI0N9WqtQJ/kdJpu8/JxgQvtaG3GKsZPviCM5XdW+YDA/
utpfr2rF8aslcUlwNT38qm5ik7zUp4Iuhf3q40Nk9cDXF57e5cdWOK1MEaMcrlQn9WpMLBXAWAbP
IaFQ+GBBwd9D7+Jph3hwOi/8sWOnu47dB1yLrnJptT1KKDsT/ZwZQC7V3VVDBdLtoqa/kEwVAALA
El1r64q0g7DtDSA5IRNkPC9Ux+MO3h5rY5fZhm1+ON0pQ67TduWe9lqfv88R8Cr5fDDhSvUBdokQ
/4pJa0VrIk4SU9kJ3REYYtz60XeKDAH0Zg+ip6b5ArvBOLnrJTGfs//VVZr7W/LS7QjQSuB8v48d
wpgebt6PuQI29Pi0w86WJaeUkAFKGOAH9RG60Z8OQq8fERGfeFzrYsEJZ3tUP1MmtEcyaoZ2jS92
Fw7oVR4J94otKfGZGf43zN9A/L8PfUMFXdvBVycdTsb7v6e6Zp+jKznTt4fUMlx1Vau0g7Qyj0wd
mgPDHmviJXxPf/A8OFjkdANiQzwYiFYzOyXNmIC/IfcTQ475c3Q7/2HQlGsVqNIcmFWn3MyoFakq
8mLm8QqZAG/WYHVkMlDsRyOJpbjk4cZHPoaTyzjsBuzLfaomj5hdMFF5zrl1g0+Q4u4QYYMfZg5/
K6GMl/D6PwqEkPFxnUPICZWWb1uThc2hPzQ5hW7C2k7VT++83mc/IYLGtIULp+BDSAx/h0Hpr+PQ
V4l/Wb8BJREL237GXILfFvwQzTYZjtCuKZzpttL9rXeP95JpiT99Ov3PanrZmqJq2um2DKNkF+mg
pEv41EO5P5J2h9A2e5jkJrZjy7hMtsRD3hazW8pEhpgwLpHAx9riKQa0k/0T56WmRT/hbvw+suxA
b3Js9J9NY4wCda/TWblixlpUcGBiTj74KPrYDUiOaO+/8+KHrO0e/xek5RZlK+G//HTMkdzOP3x1
NefDz88pUj32z34mJrfJNsd6LFI171wgaSo2t+KSZYrxmtzh+J0i7Ea9tVH+09M0btaTEGYeuykm
RcFwoeIA9lIOWHlfvk6l70IGxe+132BUI0M3atHe0iEwmXhAnBIRmV9rIEnbHKBIFPxoUVTJGvBV
mOGZtm/S5chMkzP7IiY4opew9a3mrfBbW4k1x7vsIuXGGSTllK3IWAiM8Qt0weu2vQAaKVn5/mO1
Oz2Y1SsOP7RTie6YYA5iMqGuklfmAT14fJAw++GQ7q3sC0jAAOKE2PLOuucYFWOsi3D//TZHBLsP
xDugoXam1PC/Xoi4sIcynARVZi4cvVGJevIzjbblrXFwGChahz2GRlxy7UujNr+HUlt9tCmWdwUc
XEq1mlGIuQ7G9o9/jUkfD9i8yYaXLF0/SqSeNo+uSt8W4q1MeE88EX2aj8SOMghaf5JJxrooVFFk
4FmVI1MsIBuSesuBzyy0B+HOhE9NAW1LqYfU/IOLwVJP7Dlj0duAMvAjrMU9mpF6rJ6bUxX+xpBR
NWoZw7F1uR4Tgq9lE23GuEBN9zAvChs8e+Acv7/uKLeLVPRSAs+0CBplV0bJde2Jspunw6xG+hVz
kYVkbDjw1JJZeOnNDLIe2R/rN3JHPNRtVAQzcE2y+cv3xRm6BeZQvVYVQTlBLi/J4xpQyRbs+JyX
n8yW1lNB+lg8Zw/n9soGk8RdjPlDiIC/SzAYURGpJ6iHx75421/5+8MwUucJ6gKEOUCVI5CpDBM8
6ndk3aXRKWxjNrNMmIxmRsA0WcwB4tF88gjXYyAGLK+VwVTsaGMXqDFe0fR4f8WJFzRRNXRK51Hp
CuA3283eYqJ+zeESeGVoArzCrpyMRi/S2kbMiA/ygLIwjNMp0bdJxbSX6TR3yKQqU2KKZUO/R6sX
dmFyWeHQEHyS0atb9F38tQhpAA6BZextbGMbkNoRWGZZ4J0ZJqSh0I7sJ4MciDLkaZ2OyyaskG/t
f1JnYqJqM+96OEqSA2CjoA/+S57OzXB1PKsPhaVUCjJtR7GRWdBDTu0zGV+pXCvD0MiFgeqbz6SO
tuALxlnYYZmWH10+LuLgE8Za017AWAOCCHB1PTyMTnFnmSHONbRooWb6PsC66j8KSigZvWQXMgyt
XLf+nclvUROJZG2whHf0Vju4JXMLBbFKHcM1RnFHIAGct+Yk0qsiO8LVRPJFZH/jO6qCyWqXwVcS
P1pDxmTrgT7kxC+UD78oSNIDa9HDR4bKdgQi/VehBHaLinvu3mwMmf4CJ9sAxS2HG2POHTrhmcZo
UyFMUZQ/VQKMG9FpLKoOlq7htYCp4rJnwh7SHemhbcj+3/4gcEz78wGBM06TRA43tzVhcE/PnKx2
0XfkVpPddPEDBeN9GMRu0Agnwo8OVHPCxyWNv2Fzhl39n92cPy0uYbP5nB6DFnBnTSvo0aiEA25R
X42ueSakFHIBvrFLUcKUnpiZ2NwIUAhgX98/txGEtMivnHN6RMPKmmDuavSOissSWJ5fkA9X3bL5
iZyEvmCFrpz94ly9Em3slwijVBWT30+xzy5iLZ+oLEwrOmdEP/dJ2++cz3Kb6KDY44xSAYa5eHzO
1MRQeIIhbMkBBz8fP2fhA/OUgy5RMl3PU//aDAHjzmYZTp+7VpuzC6QmqEXK5MWMlEiTo9UeUWWx
gA8GeB025shb3CFuF1TEDr2M3qxPTYI7hwUGJv0xmg0olYyXHEa41jnSTi6EPHGPKdTquPS7hewD
XP9VfUZyoqh+7IUCr+CUar7bG6pYDTXi/api42I1igAfhGl6krc3vP93nSRObqvZbDgxsXxbiZJS
YqTQVjs+W3AAL4K/JQbzInZJmoe2ptAUGTsuN5xhCQ4CU8hyd0fN4PJxHP3QZLE5bZZH9HS0O0vQ
VmGPxOIjYXjgZLfusGcUFw2vVK6KNsSfq+JFtfbGAXg6s403HD5bP0D5Dnh+DT7o1PZ43eK7oPs3
IPzuNJ+nba5WUdWNFXBpPgZMU+DUxYU4uDM8QkTEGqvyYVJhkKtGCeCyDaSgMWIWwvjxlZNGirLu
6w1RNTJCWQip40rroNig1+p5skAF4guVee6haZBwwsUB8vbpVKU5OzGmc87WsJ2eBMHxwhQ/J3kA
xrT7FADi5WYM35JqUhqnq1qOezGsipzlfKiL4ReNhP+s24QS8VNSgt85rXzb0I017UYUBc/R2EQ6
lFVYCfOUAB/B4xoR7kUyoeT3R1xYbWqx6t65nHhDGXBVSVdhjVT0C94VcrS+3+pEqH6ru/WLcqw+
XKVJOUw/O0Zadfh3KWFF1UcA8r/eLTrfEKJJED/EUwPqce8jb57dnrKt6EGxhZ1Gg6Jxrhk0PYzO
D90CD0kKM+bihMoqmBLiQoIzwFRn9XS2IIO/R33nMx7PHZRUb+Kq7Un5JrWErttMl882RG+ujAWi
7aaZV9RZIxLeisJ4yEoybZuuuna13JpMdZVUXCuioxJhPBwBRs1v/Ht4BFfQ86mtMJ17e7agFtiB
c1WwMl59MSvBnVKo8IhyjgJZZ7TrnYg+MQNn0Y9l/wQvyEGPLdsOrf+JmwqyOFu6hJWJgUvY9coP
akzuyIGbyp6FoXKmMT6/yj3gBb/hX5hHX4E34wLii7yg2Ig20P91LpE1PuqIaYiB5uGC/w34etaM
D9lKry+bfNSuwA9tUuOuuWuLdFOCaFKS3qGqQnQkox2QBgDjlPDucSBmcBxY8blfNrsxoDtIrAey
sm3sTPfZURQGt9nyo73kMbjRuN7pmnoNact4kFRjin/0Jk1FKgQp3zBtkCKgieAQwOUM836aqC7q
MD8TMigSpdqDCBf0nObjXx5jB2LmOHh1pSEKEzsZ9rtBLaHkg4AzpuXk9Bp36hbHLoKJaunF8Dh2
MMYZ6YxSRHaDlpDKX1WfHwkbDymiOa/4B/H0y+AoJ26zVhA37zs+UCgUmob8wIDvUlwJKHVQVbcA
VGc2aVn6eANfvkKzgrz6CAunkPOcA/2sHALvWDRFH4popNNR9QNhu1TDidYnRWYW++RzBvt1Z+WD
7gOBhrNb8SXYaZ5x44lceFUz0ZY2j5QKeYkOOoWcZGPPA0gwLOLi2AvMJmfh0DmP91zFpUq6iHyq
PRKralA5roJvE5tiAsVzxgJsN2uf6QAn59uNx2hZzrC00HKsiGDsrh8S+WtWuyv0VKcMk4uW2s9Y
vD2dJQ+P+qQWJIaVfogi8XSxKhteJ5Ec7OHgTX03dalE+pBjS//tLEyBkFQoaVXc/9k40LhUe12s
Mg6yMnI9CgM4qITKm6OHYKgzcxiPjV8vzg3eLz45n/JoK4PUP5OfGsxiLu8Ub3sA4yg0t49/lNot
Mxipb1xz+J71eo5npcRa2qQsVFo9J7kQTRemSg8vZXE//4i5J7xpuzmdWSRjDJug09Dw4wRX1qdk
oD15ZBwS1pIBXy+SruxD2TUe3AzcISpnZ7TzCh94a41ZBgwwfj7JCkzkvyQYOEDQwFAS5YUd8sBQ
ns9RwOdfjE6ACMeOZAfkWVbemPlNmpJBJBMIvmAeUgHtjhuZaQQUQ1nF3rfjh725Bj4+lWechQSS
xjaOS0iVJFX28SSA8HOKgQFYXxbbtKUTIQjkNvIzrygEJUNzSEHZ1T66JrjVyqkAC0zdTz1U0IvQ
oSsNhupfWkN6hc7dbAf4sNKm1KhhmB4WDJf+VIhzJReWsiHZlQIvMVjahDOlDDn9ihM9DB56qbP8
HS3LnJI0K4aGNM1MBHsVbPb6X/OrL1VHInTu1dbnYlpJMdyhvGjwk+O2XrO4STbQ+gZ06kRMcfsK
j2ceWcJdfEzHDizoSIMO2do6TM97qFsimWQvspzo2FWKYgd6OaSqODe5Njzs26jucdBOmLPNZELI
1cZx68OsgyWgAKxuMGSgmeLW53rQU1Z1Dee9Ab+cTpoJ3dri+iHlafZP2dMVh10rGWImdWeSt0YN
HeNVpcyW5XrH1gQgl5V8nHMH2czweGJ252Kf0ExRQs0VirBEc4JauGtl+Wgw0wY4kNNNM6gFJVJy
7XDzscJ9gmFpk3JpNdoUsK7sP8DLeRZ5zjrLPOrK9rpncgeFle8VnRn2jP0zdbjoOK+tH7QSlWZo
4DE0LKx8XxUCRC8BN+fG47zxDlEdFiV15LanB8f5TNkSYdhQ3TWzZANjFV+c8Q2iTaQr1uX0L9GK
Hf3XOdwNRk/l6IhlMa07AfeUTtEmvzhKPcZrzwldPIiK1tnY71m3CD/B6YgxRbj8DBGsxFfcMFAP
+T6uLGL0uWxhxor/9UWZio0XHVks0FdqTaoMGrPOqF9s3T4jGXFej8MwePNVtohAheNyWQik2Dyw
k6M+Abb9ygCaUEKXM5EBw8G3yBMJDFCdJZoXHK9MtEP92e6qNkFokPxDS809DuNvYUzKt2A84Goo
pvyVUVq0d4c7OMukFBd6eNTOH06BqF72I7zPFoYJiGdGUsrejUFYyZV9ZIYGxjnWkFUQTLeWL86+
SeTiQOyt7CeDDeWHDgP4Pk8Vc+htNPlJVTimnDlU7zIGaMD7e6hzvStFnPWwZ+0RCsqhGQ8eOO3c
B8N75FDxctUjAtOcjH3Vqc5I4NrTU/a/IONFmWNOYZz7EuA0xMQ6914dcCIn93l0IR6BU6V8PXwQ
bOt6B17t0sIYSipYGRsV3xpwf1Gjq0KYdArcb5si1JzBh4tMREqP4T8GlkKeEyLK2LIA8i+W5mg7
0WseILhOmTQ3e/mn/nhd6HHfI6Y7lS3cko6iw2hevmV9RebvGgVprGfWIQi4na2GEXFiZbf5fw80
ZRHN3zD7ziAr748t4pL82joqumVyK3Bs9gl67T4tm9wshmvl26XJRbnFEpN6phJdViRex7eIxRYu
p75AZpcjoChoNzC1rLF+7TPDvvn/BWyirO626H0llzKztAdYe48Sct+sW52Te0sK+XjlL4ZmMdkB
1nqm0zJVf5V9vhLF0GS6rwBYX9ALDjzRZOSfz30+1bntjGU0tKx7GgZPzDp6Bbx9gn+UW6ZXFBVJ
94iA0dwb6EVt4CgYTiPtvso4+5HN13eWz9hACiIZ3Qo26pL1sZmd3DfvdwJF2hEb1wj0uSRukrl2
UdzmwwpL1Lz96aYwNueSO6D9kkOUwIjCMlI24a0MwCW8hE15i4VQOQDiyqQlz6+rOC4fSMTSGQty
ZyTesMaWE4WpRtBm644bKVoJ02zhY4ryd1E8bxLCYq05+mtl2W0uT0JqGUcrkH3+TUbA+P9lGbBa
7Zu5v/Ta+jlH19vqltGfkHTkdWGydQ++auUAJhpm0ZyofOymwxQQNQRp7zS8PmpGSWqRXiLbkqXW
Y2T9HvMm2UXa19ZGj7v09pFQeneXs3TDvxnSyD7jpxQMjnAbOrVIOC9XFYRLgV353BYMKsPQeuHT
hjypx1BXaxRnQtMD5SkjbVpfz44t4t9O5nlP8PeUBcp4DsST0ijA+jZ3PamPPJZotXntesJjS+jA
F4bu1endlKWAl8vmml/N6butVjlxk0cbM3TRgStJh92Mm0EdYfbNXPf7xQDmn1NXwtD2adKzEpl+
cnlIyWT90jTAqmukcOSxtIlVJ3l+osG9V7e6+y8GM2v9uE1TsAHnmifwprsFEeRNpKGBCXSXB0sN
1phK9D8UkT1W1M0+Zm6gNz9QhL7M2Smg7qoghBUq1QXzlc2WcThK/LHoGmOBvfJ9XSEW6YuFjy8u
YtVanyiyiic2ZQxLv+0E2RxK/QIS6wwx1op1/ciqPI2gVJBam6Kz6p8zWN0HzgAy6sjMjIE+dnQ9
RwagpHB4dTQtSUHwzRjf8e5NHNxnDaRVfNkauxmsh4ycsT1NGtuIB0brBKQxqtk1RzuRzvn7+dMP
fbP107aPjYkNQLVZKgKsbzGxMAt9cpJ1NPafZH4xK6Z7q6n24RnnCX3gQsm5fYU5QMnh99PwRvpF
gFWExWxDwuizMYpyl/EdzTABIpXRsFGCZnT9ZSp8koaq/wuD6g6KaweEj3efzLwtxk3IPgfU31IE
3v/2zvFRFkhbZmDFgZZoGe9Mkl1wzhIsdZwGB4mK82iH2YT/SblKRY3BVFRpI3v8O1kDEz+esf/o
W1/ZbEaTq0FgQZPPCkfTbqJPjEsp+9U0jPlySCYgsZz7QbcTB+ys7LEe3SY24dIYoDMDpn2QxeaK
1+J4i3osXl/A3iUQydOkPl5ULUi8cZdv7AP5c81xzZePtdk6mxxciMU0V3e1yEgHm35Oedy5u/ix
uDUcN1WRjWQUvhA9mnI7TopFCu3SUe3Gdw3nYW9wpElugCy4XI3+RWOG2Vd8ZMgT8X6ciU8sSYeA
CcegU91Tzoco4wJ0PfDwPfTKWhhGUZ3uilN+SvWMEpsVF/IAPj8dQKnWpGX1DC73EJ/twv8BtCRy
FjgYrNG7MAVq3qjT/m8PwRlBAxJbddw7ULvO1SnqHnTSrzALiZqvT19Qbp1TJG08qpSZ2pSRFEa9
Xch2Sf3jr7LRfv0qHV00WLx9zZJIzLikmVK+mWITQ0/JpnKBH3uXHpqQyTBQW/Weq2JRwvY9ZKl8
zjOdj7pW+Vv6RpVF2dJ+M86w4ASnTBWMefnLAyG/74GDp7d79Mdx9ZK72ky1qyRKgE3BTYnpUYb/
umW1vY9Az7FtW5A4kis6mjFjitKax/5amT7dNnSv0lm170/HtONLhMA2jYl6fSfmTUjfREVxQliR
wrZPqaILm4/XoSFk7/3ns+ThEAKZU6AQusMsZUFYWqKZq+MXfb+DjEjV2TkM5xZnHt3g+IhkcpCl
GNpmyXU5p1C2d78Yb23odqFNVoJIqfvIx2qdZaYV5txjfG01aOi9imZC9FWmpwU2OqaCC8oy6/Db
EfJus1qojdU9TiFkJC2NfWVo36DMhNGIoYj4w7ppLPMCWhjzIoApjcyluAGgZuvZoFvCZYuwUSH1
ZAyeJSXWXrndf8RWypQCZQA8i+hBP8x45NpH6bRaNADKymu6SZvHNfcGkmXijNHUQFtqSECFyhg/
3aSCGIftlzWdYX/ujIDzS2Xbvn+rinVfYlAL7dW6UUHiJxdZKkXIOxARwNxR60etTc1F7i0osODa
WtMKVT4b3vpthNwKUHDfQVigv4NSGb1nLd6zlVgILiHMAI0dT5ZYFtSI1M4GcUBI4C7WUAGK0YRb
o85940DbQZT+ErSNA42/I7mjN6XncNO4bh4bC+gLIvK2J+GcutauOWETpWdCyz+ha9cQzWQYnwFb
11OcaJur+IGgTsaPzCyQ82rtQl3Bna9c6jhWmdyEWoYW9rik/5S+gZYya4yavqM0H8cBsbf918mC
yuyCdrnNlBXu0USDyXHEqz9yNvVdjTnMd2IauARWZbRcPrLSFBU+OtlrqQDyR4WCHnwx4KATO2/X
f36VrW+DQBRk8rL1v/N87ZDqI7fwHiLktv7SuEBy3JqYeVIKe4Oon2Ayd8A6lZiMQMQfmyNLP61C
oTWqEtwJ11r6Z2C+BwXIY7K+NryC2+9pGLxbcXsOFdHxkMTiO7XXUm/QcRosKjIrsRVaoecdBrrA
WQVlBDB+vEKJzIrTt+t0taN8WosZ5PkLYBoLfLwQF859HYSkEQeEegN0orWOaNp7m8CCFnQsdm2O
jLdAv/lqO1vhhxGlvV3lUFQ4Lgu/Y93qDy90GY9U9Z/m/YDswySVs/8UXzLkr+QsPSRjmbZQlDwa
F6DfKfUq2sBkHwhkk072NJ/0bdy+FYPlRwHsxLiZhqTJmWLjxgVkOwPUj3CMq4AAp2f7wXuYmEpb
0q+emCL51rpJ6aLF5kWpRkp5xSJ88Ki62KdNFI8mgg/Px/nxGRJjluFoCdAScmvVMMggst8doedF
qptGkmoQAeS5pMcVkkNZixRuG3ENFBW9ovyU/qM13Z3d0k95p6E2zkr9dvxXNmRIFqoDHKTi8Ur2
nsLYVoJr0abKnFFjR+L7yJDwwMsyUz8e+3TLhbcA0iUa8oiRDcBMsWJwMgGdHBhLMcALp5qStAd1
UtLruBXM0o11JnaxSgnZvG+yINlDH1gqf5cpZ3Z0Q7gOS6yS5J9Opkn0ooVMj7QO9Zu4lKnX4+3i
HKhGWVN5N0g4ZXquV/y4j/Qpmb541GOfTDMbKfKbKx1ubAhYLBleVeGzM1SkPx6CHLdHtNYZw+hw
W+4HqFNl1mp8lHIXtl3pNYxAT1acQCjYiFYd3kY5eM7gnbVOfJqCucGBNUTswSSNtipIsK9XejxU
Wxw0jkFz8SJzgejowXmVW0Y2ch/CQegLu35hmjIp56uH+cqICuT12U/FZF7hyY3CA/V0MlwmsxN/
j9BpfLy8tibzCeVnkXnjHSrsVFcXtvKbtgq/+USKxrA9/ZIx3h7JWPFgLNu0eesPX16mkayg/fs3
YomhCzp+JHw6Vy1jQ1uCzPaVw6W/hwWid5YtYiLPrnkeDGUu+S9CuzjK4fdnXZY+/PPKxFZIpLtf
VW/dOhHM6hQ+qcQho9B9ZsszTiHUMYBg9xc7t9Y1awjACR3MIr/vgFxk9DL7qWJwtVQZLb34g/qw
bhGFwvaqH7z2j3NQnM04Jk6mDfurIFJYz+RQcY3kAEUw8VSgc9kI0ZWfj36H1AYBOwq+V3BV99HZ
Lkw3BtnWoyqdVp8dm2qFsiARoFR8k6zU0WrsGVYRNYbTfWf3KODLOecnlDToPBfJZnH5vsgyf5qe
yhLpBnZensL9biR4zYApuH6tQhX/6LF3KzyvJE6pWIIAzKleVqNfQ4it9SUn1SABEtHv5zO4gWc/
9zoeOQ5xUGwSZxFICB1PQq+T53IFaLQym+krNBICQYInxfgoEna2xyPfvst9QdYzmFKFEYmqfMEp
wjdhNYmpSq6W+hXuQdRRunCrjC+scPU0c5zgNor4tNLJF6OBhMe3KjpjpBSQGCRRL7PshSnOJDFo
G42pWhCPuNIqpYQw5nKhd69kYejfeMRLwGYZrSbetPM5L6TJCv4Ku6Aqna3ECs+ZB/qwhWy/TiQv
BIk3SowjaI85XonT/Rieqj63fl0+6ZQmONn6beq1ZcX+jewaYNAIM8myD2j3FrR4fmmTUEARGyU1
IHLSnlEA07pnF8mBR0rlzCBklOq4yVCifqLmYx1elJL+v9Ub6HkRM3MinEYlN+oN3fvW77ItiTZs
hVyFCw6NcZuADJ/tJbtwLi5p48upg0EaFgrLre+FRlKkzqRzJb+yofswQ3UZFUBhBpD6yZzZ1f79
9PNQV9Oiz6ip2ejoh90R0LGLF8gVwyep1uxDrE8aELzptkvwAbY+JsczI/9lYosii0wBAx3o0iHr
rC18yJiSG+eM29XwpbVYdDxkTt1qmwpmIkMug89hEmuezM16aQOT26OICb/gVUlbdcFY2xTG0B6i
IhuvNkYeLVufC81jmtPchoma4MbtPk35BF2PTznUTl0N4U046pTskmpVC2GmKdMWXDCAFBNy0ZJD
rWHXu6WeAKSmLQDJJAT0Q7MaHY26rIbqZRPOy+V0/83FFEVwq+cT5F+6mDecPG5mg82oSneeyzZs
WFYRylsty4MPipPudz0lRaed+NQ4/p/rqz8lwK4LgY0aocqrY7t0eUSG+7cwV7IFuGB0FF9ztEDh
GTwwBqaRIk3X1q8ktuCMmNXZggWUfzuG0sphNrDDTXkPUDCsNUoJpYvM5UDNVT4UZ4g8TimX0xPZ
6mRciOi2aa+XDajWPe+PMIYCMULAWxiKVZONYCjTGgIK00xPkYMUirGSWzjZUXBU7s3y2T6nvWEE
HWw2jfVottKQkbE04d5cowaQgQnjHzgtx9cWtPRE7sq/LGmOa2pxTGWOVWSUd3KLaYnitLLKG4/v
sAPG0LKyJ9Xw7LLQNzHJfaXbMN/hGqtPl+mfZBvCCmAYG9Y1lfM2ejIiB7AG2hxyKBh6mtQ5wuWh
oWz8ZNoZwcjTTYyI/54rtcVEhaHeRmGQiq59gFIh+OF7Tb4GTnHhBN76NUMc9+MtJAQ/rWd89En6
T9kCXpMLBO9r3Fr8KA2RslK6aR6c3KsEH/CRLOxM/YvvGX/La5/PmQIy5r4c0fteraySb3/gALTR
uNaEuEVH86bZs8rQPwWzb2QEcvG3CVO68X0FvEHIuyjy4LeTfO//FDLa5TiAKciEsc/F007KEjpd
qS+X4MIuHuWNZyCRutz06PujCKuTi8cxkuHg9BMqm6Fw+EDn15hSHV2FOESFwjAbHSRU+ZmhXJmf
7avi7JHhggJpHHFLeMQSxZDz3lPKcfcrb/KFLo0MikMFRGLE/o5rCZ1QFFZc8UbQn77bLIuxAFJs
yV1dz8QhUlBpLsUrKo6Lqa5nPemXl3sOv05x/g/FfiAmWTr+em+uKt3XphV0aOvGcuo0tHqU1R+V
f4KVuIPb4LAUsbrOf2leuw+SeFzs23wPvO6bbhazRJ+BQCsDquMzjFDzQejqLBS0XX8DEuCBtPi3
xAs/vTyYqOPSlav6cHzza/oAD+GCH/x1OqWYs08o9H3m4Y+m/S/4L1WIXVyROykuznOovkP16O3e
sYRVssEEyfzacmRu7ZfpbYVouhySE9k+7SnlffuhYgmDDpsxEy4F9MxVseeGCPH0y4mxFzr9DfFJ
Md8APljHZlKtZZqhV4SpAfGIRDMQ1lzHI3JILj/3DsRlcGv+wLIw54rllKic5zo9gtJEbtUqrrLe
N1tP2+DMy0A4ToaenxgJecT21ja9w3xy1M9JOYzP4Dyd1our8Ap5KZRT3/6jJaduQH5wh3H4ICo0
kFmqKQ3fBroANMdKtKadzMULFySuO2X6XSS9ay5CFqxAeQQX+xLxcRS37QsEVW+UCQ4vYihTUluK
snijuWkoktRK5GFR6Ig5bxBNDFDHBgVgWU4Uxm5HH4+EauDMTHBOEQfTbTL921j9agS5jmJi9MmV
hNn0+/1aWKwo6T/SPJmDIOYhjtxu/UJ44DA1vjWaeBZaq+3QtS9hgap9vHHQrpyU0dX9whg+K47h
a0+8Zc41lN/8rWZJ1kQ+9kJfi3jkYeX9cL52Rc+rmAmK8v4kjvzBOBKB8dfvZdXr9UtWxW3KU7/N
eIs6DY3/CDQo6vZ3M1IVhvThQplzgSST7me7avtx4Lrc83N9kiRgGfzvu8UgPLZdDZA08K8kqGEg
qUCgdat5SbXaow0+2FTkNLbwmlbbde5yLrFfIE4ZgtDchjCc/WTAN67ZuHX3oBRcx16pGE8bNBFZ
JNUon0zodbByVx0TXTXBNlhb1j4j2EtOT+5RyEVVliraf+hvI20TjwHeJMd5pnPwxBlDN8Nmf25d
YTZU9XWRG6X/5xd/7SJblOo2U2YmY7ANPxKoHrWiAOPf0KCWkbBu2S/xQY20C/mHAiJekiLIEREl
zW2RFVz0mz3FtE2Wx0fvKmBCFQUedcW/uRf32yVyKoJZqQ23K58YyMm5d9tanbdv+28FXeqdhX/K
RK8KQ7WGqFSAJRY5ZKxmYTEFmmhzuUOYkCOh1oxoVRzTc92Y+C2a73+ZA6sDQDTnD99weMp4G/g2
fMaJpUDrJ/xWzW0hzjX9s7a5x3TxI7/uWtyxyEIwjnfwWB9/dLhl9O8mJXRo+HidTGyhjvyAUG1T
lP/8LJ4pVjSiM1/uCPjS6kB2CfAUKeQOyUHnAJH6sUeHMYScvUduk4cP/Q9Tt3/mBPN6c7xrbHS+
0Y3KfmERpbnqEH79V0bIdHotDoYYQ07nafye80QoaojH0GsofUYmyzVQRCkDkw0Bn7eIV5fhTvKM
AUZi10Hl+M1j5crEhWPIfr904spr9cN3jhm2B7F/tGhxfq/0Gla1DZnrsIlGnHAFU26diTNNcCBU
kJht44mWhKTTkeNw//WeJIrq9KvnzoNlkqeow8eISeeL00Qxt1JN1AC+f7b225Vl13+4S/dZQt3p
vNK7k7W1sPrS3rMysBsHJOiuoIhqpRYmpUgEldCaMWWE9RCOYQ6kJiBvrgVp3tV5HRJhE9SqeFkU
4QpwWKBPvrbmLyFrdPn6RBFq5wb3EPKQW69cbyJaRI2Oq+rNnXSjHPfxtWNrr9sYnW/8+/3PoV85
gV1ZhlO1DR7rR6PuqTP+CNSlqORN4YGYZRx+0ktdjBFM2ccfDSAh0AAi8af3mZN7O3QDM2gRZ1JJ
9ZhE0SWK2GJktpv24mYwCUo9jDGUvw/T0PPOIM3oF9E0Pxq1ZvZVtpD5xzaIZhx9RNFSx1o1t/0J
oYuGHEQmBtyGCXaohjNnYb0mH1fTJPxWmNsGKokDeZ8+5XPZp2c1pNKN0FUJZT2Xg3IITFvtTpQN
K7rOlR7uKnGP06hlwE6oEyppC6pqS7WA84OKw0RuRq1BulEN9Biv2GE6/pbxEFW4j/kOS7JGtlPE
ll9FVsDEcscEjqs60Xp4p5hBJZbg9lP5GAf1ffc1MxATYrcYga60JXTZ22MR5yikr32GXpNI2Sau
1G0FZrbAGLAFM9DF54eUWfHfud2lOIGDAPJTeqh5WcKcrVjcR0vtovicBIE92CgE9VlHQ8uVc1B+
KCdGWxIA9f91LOOQWAh8boN8zIAhpz/BuxdMwU8PWascJAKikFywLTcNWPthItZ27FIh50MEUH9J
4I+pxDVoo4R9ho6Dt5bqyW5+Z/21c0wOJPl3rFXzYBt0kYw64CrDyVX8ZpK9TjTQVBcBlYU7Y6k5
FOxgK/faQGD1GDLUnNNenkF/IWIbhKRgEFXjAH8w53v5NgVooso/g6ZFtMo//UwGbe3lkDT0FnY4
O24TyfrpoqJVYiRybKOpEVTlOXe92+0aP+SjqCHPIbf9GqvfrSchRS/TFaKYLrz7SntYQiNp6BoU
1aWnqNpkpgHz779DevBTd83JqGt94mJh6b/U3XH96Rw9m7kQpPRWxJCRCchRwHOdZU18T91R1SJu
JSFid3v5NrYmfXhCzAEMHIl5nPMQZKqixixUsJnBKTtg/PrUxINC0o8A3EWakr8Wg8cdrow6xl3a
Sfg6wXCrIm+Y2zbSDAIvZtOSWdyZNILkuzbCnPuRlNq4hU+jAVUFch3Oi4Nro+V39u7uzAoioHTx
DBqIWBaoFeDPuNThaK13+ZPuMWhaG5BhFNOwtj3O3z2oodKMUg8i8HW7Dve0qROGlbckhFb4dpBK
eHbmzMncMAwAZ4uuAAFBFn8YFwMR3R99RUYjvxEsI5BMpJyrHcWGt//1S/bXqOR/9XKE20myx2sC
dsSTjrZVY9AU5PrRBs5vjtHk1Vhwa9QAmUGzhpKZRSJAUyXKO9vfGMf0sfYlXFuI/i0XrItVlP+1
nM51cB1sNDYRVhPlmVH43q0pbTW9Ilt9Rf+0KGoeaTV8Dhs0cVHsyYMSDooEGHxhGHWZEIpvZWlz
iZqiR4/RVPMxOmDyukkXlhGFNCl+HxDw8b5IUizQ5ixj9zv0whx+y6nhq/NyE7iDk5Rb50rWmkOY
MMKJz52b2mWtYlRYc98S2zBOgcX4YnhrDy7EfmAPh5O4LdVtZs7DwaO7efKGNupAqaB1gkrIhbU0
OoI0KJwymtrvhmkzb0HMllJv+ayTNx2qnxBstwsp6NqMkBG7Lx6KKeKEz8f1buu11QHet4/+t73M
9VTriZs3BRuUK4RxJNvQp+lLyBRU9hIyUAXQahPeOvlFDMi2KObEZoufDkCveIdz+CVoc1dyS5z4
9eaGkzgyBFaaEdqUcw8Nlx3/q7SNwe8655+k8ZsOQM3+SpG0AhcLB3sIQSUGa08J68JhkRe4tXLW
oCJqMgCaCTbEBlbwM9aHcXi/Uk3QytGNJvYPHusP4lOVqqjiOd796FK4ri9FlgJG5bk2l9FpRyI5
/EuNxKq/4aF1ENjHruiLtI8IG2YfO8D8n1oZDG2gxs+TfO2CyRUiH2oDw2XA4TvFU5AVH9ZgAKA3
gChK3kdVvg37cA4LbQmg7N9nStIykip5rcjZcbIEwixOFSk4HZJAV5hFv57vIo6zs2HBkLFwHrxm
AbtFZK2iOo19FowstrXL2WBAjKApeBzY5rq7vb8F8ff2vfJfUnJa1Ota02z7qmjOnYLmsZ34mCGq
pW4fjtyfWkM6n5Tmenwny5Kyb2zBk5u+gLlDvlmzfhM5PqBuTTyVULunil2S45PJZmtrrOW4x5XC
8JghSxlnRykhXp7QHbT4vrEFkv34G/TKHroK2uiJvOGuleyn6/VKG5so4Z4SQKCAdqBOhp7lTHxI
P/nEGUgrDe/Uj0fbU27U0yDc/Xz5Ut4cviFimf/i732zqA7DsCb5v8zlVO9kxqxLXus2KzEj5CvC
2OHMrKWjQYRbi0Aq65puhOF5b1BD4LNaRG226qImzmCW3yFLxHjs849izbW+ZvYeDjBMK7i4oxrb
Cl/ZuZ4OS0EUEZytmZqrTpZeR38xc6GYrVdahVOD1/UkcRinQsCBwqS9Jv0al4yePxnYgv5DzY1F
eDtEPwOSSbBmsK5A7On+9Odd5Njizsx+htTe6nqdLQSq+5lm1e1ZkTmzugciEeJqaPbyjq7wZVDM
hGpeu0o7a0GCU4AKEjw/Ivu9btw59ngY50PHBd7xIP1mAaZNKA92MVA/71dfNj+AV7kfxfSlP48D
vpEyDPuosI3jqwCcXCxXwM1ZftJI0NMtQtpw/czNy3hZcaHTVqgs1xy+bYaPAoOnkPqu+QkuFfGA
R+TpJbDGaGKT+piDWc/5hxj3uFMppvvS9wzp1A2SMxwtWdTMHjTQ2QuPx2rlBbqamLmkvTL4AI7N
gr24s6wOCUgrebCIhmnscPvK4LmqbRs7/JjIhz1ShnIDlj2wBODh4Kid+g70CBRrLtLN35SpscBm
0P3g1QAZvUj7fbWfVeMQwqEHM5tuopavP5aukr+YgBKttoVsoHLJpr6pJ8pSHSlHbtS+C5XW6sQf
WgDrpI7wkYHk5P4JzSKmficMWoAM9PSo/Ei4tGhb4pW+FfseIU+N8aEBNkJo5v9u8wVaq+0+lKKz
jFin7EFGSfh+MsKy7xwxwy7w+fxfM2G6c/NMeEAFrFp0JIrLU/W2Ov8KaQlJ2keikGIe0xhwiIh6
6ffCmLLC8cQA+ldEaM4u4wvHvGgE7Mgh2fA5lJW+J56T66sxOBBaSazb3F+qWTF0Q9N09cD+8ado
kBAfSZGXnhmGwkrvPE86SyBo5nHTqUkcjQO0LPOCl6+VJX+/BQqRfJUWwlRnSmDSfjH55kH++LM5
+ZNT1aL5DTu7zQeXcSuKdT0QfOOaaYAi/rChbmcIO2b7MzBzU7sgrMYqjngEPKa2IUwLZYmaTWZI
tde4/YLOUUjaAEDJ3PAAvyCV5ZLg/fI25AH8aRlMiEc9XhyN30uUg3fC4RfQtJdZLf5cXvLXm5v1
goenMFqYza2QRDwMUvTzeJUIbyTqa6VOHUvG9rWJZwbhgh+j7pgnaNViqVCknNz0RFEdWHyacc2x
WvHEgfLpRVCsUE3UU0G2HonIhUxWarucnG1/spU0rhXn8kvXc9RWpt2Dtma8u0k/vWJjtvSJlvv9
D8zY0jL95PyWY3BjnPK1UzFS7qkbdMLXjkqX0q+rHv3SiA864j6DbK3PKx+ZUGbd+fqdEZp1ziqB
SnukqH+ESIWpYJ6cBWJg/9TZi+6NaD1aupyRlOLxAxZ0qBDVY7X5LzjwNhFru1xcsOGlwj0E2qbG
sh/4PZjpMKiDaIkAC41zH38cLHT8pGy5wtEgyVI5fFDIA5U/pzbza9K+BrvC7DdHmQ+fHDamjO97
rp5sUS868TKpcSKIyKK3Ao7MdctXg5s/h9AB2BJibYQSm0zJQx+ijFew7Q3+mHCYxdK9N2qYpSxo
ZWnKlf4xRzkDyDBjD1jFVnGkApkXebh3/yFr6TOlKewPlywdi15aF/4PJxvd5MAQJjZjpE/OwLlL
z0YXkxoXm/XHDTx2CzSEUerLdod8GinbGm4EghNbxbe7rHiC/jVeV/WDaDT/cj+ueA1VUsWzA73g
e1W7Pz8awpac50GzVS7P8i1xnR/yC2lmfz3ucAmjLNs5hITrqukKwJymugJboNSua6JNaq54AlpR
kjaMBPcCmejADKUsiTTZH3eThLP3+JOcO78hkHyLWz7IeYQf6G6BVJZo9mcfHdcz0yu5clq/yRxK
STvjlO/xL0/Vfx0uvvWDdAFqP3tH/a8PbJMj1Cq68bAniv1lNc8hVxZXZGvpRijSr3LNuMVj1SUz
No8KyhuI0HvyHJTMG1PEuwlnS1+vprrsLx+gMZNkiclmkngpO3sGtEI7CMPDyc+Xun8OGqhS0FNd
4ktvip4X8TKNOOal/uDCtZG4S2pOT4EKBcGnohuMbY8PDq6bjdBaQN7Tv7mRXMCqchL+HkO72HPV
M/+zpVa5nxI5xURzYRmgcRJdkOd5WZUjUJktwWXg2FmlKfMaTue6mMVhWMeW3seWYZIEmpbWobJv
fNhsBWxRnuR2G6KW/8BhEHPGP+4q88SjNvCKTE3Na62Xk/vRpL6rGOPnehGy1fKJKJMzzocWqkBl
OTcLAZxix9HMeOsFbIhSLeaGn5WaU2blUFfuhXx+DJRictcU3isRWDBgMhpBTMb8mceY0Lfborep
lVb/Iq4dMdHmLKlIrthbvkLeJ2XEswvaP+QW+cUF842ZqpuDnNjVmx1bhrnKDeUko7kKnQUWu7jM
D6uY0olmxKB3jZhqJuDyEhctiek3k1j2ar4/7beY+E6BhLMAbL7aQ77hACNYKN4UEfmNv65gnEww
DKEGq0opRbkTqJonyXgyIz1rv9ae9qhpkivAPCpccgRwClo9yo2rJ0im1RavPGaWn0CccfBWEyUd
/XZoSLEeipfsraCI7rf3lsAc0qyGctBKiQ6ekqhVo+pX0mTeNaZy9esngA5f3PQLqQzNdf+obGCe
1MHRpUIXBYrRnrSTejI5jARQwLgzfNgLI5jSL6YXjovQKYm69G4WG3qVZqZimIXx90PWBJjR77pG
sOtLP01UZgSo36S3ujVYrmEfs9KZn7MD5Dr3jvmmDhA+k04oijxh6Ub8iFC1niahQcJ2UOEfVGBo
oQN3A6M7lmowN64H/0oMhYsFLxQSZ7NU0dU/8wGNIAnh7cQswzxewK9pPrWKZI0I6aJCkHjhn1CN
0cOEUdqFfZnG+HuYjwrtB508hUdPL2Mb787AmuoCRwamsrkuNToLrVh1eECCXAJsV+k5pH3xU85u
hir6gMdnOW6jEEfYBOvfCjNM7K4Loenx+CLD6KflHfOEonJHpsL/VIxHohr9I1lq7gfbs3RXjpbU
9QG8CiZrn7MUV3sUYlB8wmCEPHQ1T2wWkphjX2PZLAkzaEAmGw+hc7AnCKHpqX2lhwB8pTPHxjVT
85NvGrpYKv1wXuIeCLl6D7PkmJxK+LkHMi+0DbdD0NpaqZLCxmQY2ocY4PXg7xP06GvtgUenURHA
ep+rGLQPbtF+iC1sIKk2iqEDCvmI653kHlLC9gMAhfoQ91y1y0XVrQYo400luoJYQ6uNPZjGaGwo
1CGDfkZbjoWaCEu/sZO2osJtM1+w3nhxY21SlD4DvFzFSs3WOFsvrNgtonbBCC1MUf191yYTDIC9
Hxj2R2IJ4RPYcX6DetgBD7lHpgvoqvE2njRXM6hM52ZSeMfqpqeQw/W21egsO1zB7+91D4z+Ggnt
G0qnTzZHuVc3ZRzRj2FdD4cSAUunjri1ucLCszko+nVrOexHEPfwNAY0r2+JtabUOK1N1WIj0FjP
cFKgHREPi9NT5IhSI8YWzAJUFOamuC9sUvHaVhEVQAFb5ULH+PK3vIUrTSEJZPzuU97AogCOhSlp
9DmB09TZYWONulDl27UibRZD9u9Ecq90GN96nqrUCXKxlYbhZP23jJRAuIGP4QLxXAy7Nau3Xbvl
k93/DpLUjG0ZwbkpSDBQSkMnuPB94DC4QZAWR2BBnxwUr/E5eQFlaOUZxSjIAKP2Lp/VKSSAjBWa
m9elchTwIbuV7vBH6rHzyZEzE+m0OWzSJbGpNju9ioEJvQhM0QnSUATiG+kjeJfuMrEfxQ3yYqVF
TLIruv+saiqQVo5DLlwxqbUztCip1FYErU/PGufv7uZwNDdPZnpjg/3dfGeKkPQX7HCBUYjQBP1D
bSalxGSVg/KbGy1LndzK6EO+mQ/TbqZHQt75/kjL8LMjyAEpm1W76dbBTe7jqdOWx70AHZPZtldy
agoYqm4JPJaz2O6eGQOFMqToPQ/K/zlsfdSbnA+jeyYKdXRpRf/YewM2MZzr8QbEq8Zjqyl8gJ5+
B7PtRYZdAIXPf3Zr/K/zv7p5msWoYOH6BuYerXzEtjeeVpnZ3iedKzZmM7c9xHDfjl0wIAOumr8b
eC/rAjWm3v1Da6MJNNXgg4/BOnpAwZhLQO/3e7Y/SqrBi6HW22aynBh5flbkaX/U7ERK7N1IDbCB
ECgP+9P2yUhUEQd4OPpHSt2PzStWGBBfElRCjLFbEC6E0fEXloj/dM8MUm42Pl6eA3wQS+qi7H8K
xFtDRk+kyl9UCivagap1pd2uSMs2iJTQwp6IwF2FDP8wJMYWTbohWBN901sYizwasC4LyO7faGSQ
qxbwTUmGhIN26Bam83/9r3uMKnMMBSA6QIdzfILOrHgzAe41WcZFk+iT51yzDKUS8kkslGhCIlhQ
5Ts7L2yTETtB2Jo/stmNG7W/Etpief9Tq/vFseVRz9208/uj+ShlRJuRFmvWGZphgTBWMqmgb8jO
JA4VmaePv4HftDLGOAkXY96lKX4TXjOOKYyjvE5UZ1tbXwQ40ImCBNegI610r/kIN1sOz4YH9cvX
39eOKRXyqvjThKvl9HincWD/Bg9hgp6NM02upC+fgZHxWdZwKfcqEXqf1XGZjYm6MobCiX1XWFMI
mnuBqQu9Uzb5kB0Ziwd5c0n+5eMAEmomF2/3CsfSbTOB/X1TQUMXc18oBiV57pQHJkvcL5ckd50z
58amV4G1upDnsdjTNFPYdJdoU8Bt3R660f70qfiY+AUbRervX4GcAdj0j1+cIL64ji9nV+nF5A6c
HgJ45k2WxVOIatWQkAZX5hEWtkf8Wjr9qE+63NnQrU1z1Cno6lgpp+J8wCxf4GoiV5crnFzNK2Tp
cslbBUiMneuuTkHml3yteKyAy/ZLmmS0jijZNE/oh4hH/XRF3k/4XuDrCEVdJF4qf07GPQTeRMNq
/VMiuLz7ow39EzZDyUT/k8Y6J++Fs16mdsIXeDFozqZP7U8Ent/qiZ8uckISr1tTWHwfdGllWUJV
hZO91H/ws5AlvlZ0Xd5AcVGeZaj48Fz5m3t0fN1Q3ZCNiuz6laU7E5aVmZosOBRtw5Fi41iPmlUS
29fNemxdrGC0eUYaE3a/t3Sym4wHI6GfJ+efj96lV+0xmLz8aEwjz7AUHIshjixq2LlbAqjPzovc
GDCZlHAFuiLwsiKafFOFUl3bdaVlUAD9RYTp3QceRjf0GKrtXfnxyvpVWHF1bNsIfqNtDtee5yMB
Yt38UTdxtomHLkugZoiEMTvGOElKvYAUmiOwVfwhQoHBDzLH3FIdc5DlsIODxqmYukS2HfwhYrWE
PvRCv5vzs9m0y7/qBoR3U2GncYFywHjE4YqEljFnM626xBdNjV/sbGyYwt1I/OHT+Xr3AEiVxBUR
vjoe9Rkab/FMacoRoThwYoPfLRyzlV9Swe72/zqInEl9YIeaUYe4nLAXGkoYLHVRw+PevVkyHLFt
Y7XI+3aokN8Z0dB1/mddXDHLn4odqaTqxYfg2CaSugsozojfmkZBO1Ccfm50vM7Kt1z0dReZCxwz
i/q6EpAqp+b4VUQdjwePzBgthJ1ZfT5S4XZ/2d28BQKzE3SK9KEb0I2IyVJSElz/NwcKc4wOZ8fm
eaQB8fP6jaX2Q3cgtWq2wEDDZSy5/FP4uZxQ6Nnld01gVBl+/6blwLZuYxNw1PqWumXemGlNjNzS
lGBrp6YvFirJItcpP9Mhxiit/64yMHJRGEfG+5zaFK6wSPwo6tL6rqn1Epivu6udIgC3H8bZfrHL
BXWtFXIMCelsGBsthSZgw71i1sj3t3EC2Ce3tBO4D2nuhWqm6oPlvgTs88czy62vi/Iuy49TLwSl
wPscduT+6KyJPHCMkFXFtGL+v8843cdfCeKt7vaIx2Cx4jeKsPQ2/AmDtF7p4SznTX+9QmdhR42s
hSp5Dp5gwvSj0Y/2ysleiOaT2T48Gndvg+Tw/cH7do2WD0onRNEq3umDBfmhDr19UVmLjyIfdXHg
8DqS3bjSK1yHA89xN6bN04HkXN+76i3enz2nb576IMtcHWGxupmcqBUZLuVAljZDeKaxIU3CEiZ8
YTUOBhKhX5THkJaugbVoepVCSGqExRp1uQwiLh3UX1eIU92o92TQSgSKcS20/aUDnGy/tXwyX/4h
yqXmDRL5zEqTJke+mJKcwFUAoCngn/dmCVJRtLpVLVgsYoKo5Y3Nq2Is8Q0m2gGO4VaCVid5tApc
AHNyzNLVsRXxoMJNcfYICGvU+Ew/aU+Wypkl/jnpoDiUaFmElILjlDaw7UtHEsUTBv8PVTkE+Iw9
W3lPMaJ/mdw3toTEHTab8whIiM4F3f46z/fjUs/zf6/USRXqryPsGIZtgU7LzrGH56f2N9YycC9w
HPJviSy2ywQc+WfFA11210I3KUuAZwIQq4ORl+pTOtKhcwVEcBe5sqjr5j1rLZVMlGAD0cywM4K1
okhk7misySdkh9E8h2n+doQR25nmZr3clOr9hWTuRkUZaiweYG7p8g6ww9qccblDkW/t6fBTRIi5
NrXjCYkFxKPeh313BdEjMBGUPBX4xKAn6MsJ0tSJUckOpMdvBRh4W/zMsmWdJWasQOm8EsiPMUuQ
VxOIc0ElpuZm2GhqbDXlH9v/iG8WC1laL5zZX7bKOR/jXUYK/eJcrP+1wnIzbx8by4qZfJKMeIXs
SqfAFDhQuX/WpydmnFnOUOUourivXa2VZaBBPTsd4/hf0xqV460IdCup1eEyX/Wf7bg3UWYjQrKq
4xienqy/9yzuLPcZICKzqGH4fmT9pGA1yYmf5MsKw0Jl+khxFSiVoPGABPkhRmhLbNyDVrfJkjfZ
7wVTDnKhN6TcKHfnNXZrkxrBj3qxblceNBR4GW37MbtfiHVdql9eifKs/+6FO92Oo280w3utIHQ3
lLXu+anT3xpIDAGi4AnyXnoPxn8Flk9OfkBrp91QBj5UyvHhMqnZSpOHUGSXYJRpsakk4ENykWG/
wZn/JCI5EqcZehSxNpnhA7R/heEJm4rZxzVp3lwraENxIWyJypjPtJCCILnKzAIutzdrjcgnjJxI
3BhgbkrbnHtpq3TKb6KKvvCtGQBjiWxpCa7/HAJglNkf/lamyTasX5otOPz1FzDHHc4C2tVRyQai
fsph3klkKngaRr5clUCU3VD7RVk0JqPzlKzB/p1g9Pt29u9lIC7KNGHaproMgvG8eDH9XNqC/fat
RbFXl1e808P3/6PGmY4WLrmzWMLDBgvV0wO51l6F++Sk6kk+rrzy3uX+mgXt/UX1DQo5W0OBiQtF
xkXUnDMhwud+2kY3KxJs3Aa/+TToMhX5Wd5H47yKGo53odo4mJYYTt/4WQyFPqGa2aJPOvF/yv3F
KwyTfl/3OOitXfGHtcFmcs3XUPMixAiqrt0uqDNYNJ85XemQpma7biKopDKuPtTCwIiWl54myR2Z
1XgEMWoPVT3VrGRD+xj42alTOv3IRkPDbd+I8M8YSH1h9oKGsRJBFZOFYRrPF8Z0ouZu1ooymoc0
4rlJ2pmi+L5z0dqLqg01mI92nIDb1GAJCMyRWZ0bXPdBvO+LKVCJC0xMu/s2k1/F8aOsBIV/8qL3
aaGZThGkqDT02oNMwx9VwUqth14c/wlmN62Soh2EHsscbzeOWKXuV1XUmdVXJ58iRgrycVDmPZox
iSxJ6A/9WhqRaRlEz9r06M11c/mYaerJyvhGlaA9uAXPczpaAqa8P6Y5brnb2B8UGhO54SmRGP2X
hSEsXzR0d9btaP7fKqJ9TLZXHV/bmfKmbg+vEqBOmLpbhVoi0f/vyjHi77XRAd3+687HtWeN68+V
FaR69w+rNk2JJvXfxSR5Fgeet8Trxhn5daoWylBS3Iyd/Gj3VtdbiDTlHKQuaxlUJXE0lSqO1yAR
ig0tibXNAWjkddtH96Y5xu1h1G4PQe/Ure2eTV1iG2mFsMEfPuMxzA2l37bq2rgermh0qxam7TGZ
c2vHO+otvlTTuge5maFAmkrOdSjN726eWQaJ96TTesbfAHxJoNuingzeDAGPQZTTLL4IDP5i+8M5
y4Yut98rTtWM2YDj/uBgwe7m4E7e9IyXTqkfOHgUGJSjqcodnmJur11m1MSP6ZVUabZxtob1A5q8
+kyXcSnff/ENFB0yS5qn0EdOPTRnfzdS6v5N2jJbmauWcHGZ79qhhM0hN9Uw1OPNHPnNWLbE/IYF
uqLXQV3vV65YkAqmh0lXI32K8BOMvmwyDeWOiSrdkiPYZUpZYYvAjIOc0PatMhoekcYHxjqvtzsf
XAMQ2kG6mx+TLxHPGEuHbESl3vl6NMvvSM3KSh8qwvm+N5CsKBlfxbbWhXzJVeJCOBwjv98mas5i
oXWmYGzJSKo9wEY7L9n3O69U1EFmRqfWnIZrz/N31pbVlBiNkgRFYMFzYidQnO2jABcqhgc2s4rb
p+0qiYG1cnQ3UC3z/ulAqj7qEP4j9eITM7g6pR3VYZQWO3JpMxJjlfkQNUF6CkWJHCKfu4EJYYWR
MZhFfSs0YS76K2UHWP+K83Ximpq/CQ2rPUY9eA5YJIi6wPbt6926D0MWGt2q3ceW4yDf72cP5V3H
tbUvHls/ldUWw7aID12oSXzXxWaQ1JRxKq8zwgXUz8I+1VSVxVdnRQXDWI/Axu4ZeTMbE4eB7prc
FVgYkBCBtSG6LUno2ePuz0KCs+QSCEQDee8f20r8ksJfsTz1xmeaBGPbLnDjzajfOfFadawuLmez
ihhz+axYSi7fT7817ofTnCWFSE2ZUq/CAsJfd0Z1CubyrvNgd32aitcuUm+lfiPQRBEoQsrs6N3I
2uLIvQBXlZ/6cfB/7F5iyXhTGuAo3luN4amk30y7SBR/hql1+ASsyseP88ETPJ19Z5yZkPOj/io9
KMC1i28Eg+xLm3kcMo1g+M9XZGpUl3bYc7tnTV+x6vKAuzo54EkhsnZvlMpFWowYGbAzDieowrIo
2dGLyWWErfTZKIr7bFpJgOU97W9H1DT5u8Xi67rxQDygahEX3bSf/UyBoiS2hHK9ONtbVKyOn9vT
tdCKgtncLshDhM1hsIsUMp/UTdAlOR0eF6aEYX3VnoV7BSnxPLwbv9eH/AG/5E7Tmnr98vG4zzSj
V1nQzZuJGRN6Va2jOxHjKYpvZURXqaMRxYln6duR4zJucu96uec7LWxOpFt+rKf/ScNL5J4V4X6G
ZIwjnRz7k0qFo1JY3h9Ph/5JrhlubyezkhHS/MHSLH8Q8JFaJZSnIXniD6/OEML7RQ5swFdNKZ3c
mf2M22Qp7HCgWeyiKYpkGyQGnI8bw176fxF6bZxsw9aMgFS/Uerv1mydk5//sPNdAhPX1b0zEKxP
wnlVIzfCbm0wNQh7oocEAI0bsBXtr10X3OPCTWGbku9dEvFXPxOqmUiYK/uJAK4h+ZBbPOQPl3er
OTzlo/oSBFjJgQS9fLWylfaeVqlMa89hDpji/yPUerPGAS9/apyeVAgD08sJQppFX4XMLOE0KR1h
xqu8kB6Wc9l/OF4AS9KRg8ZCE6euFnCk+X4zhSiBHlJH3j8SDH9dHc7HJ8NHUG6pEBr8Z+FojsMm
1JX3jp2gx/H2H6B3i5Ad1MyHvD5XdWhn3nLfgYcSif3yeGuotHnxQS7kB7xBkiCvUoJaL/oIT90U
ZU/QRNa0gvGnUlXew/yHYL34sAAoYezEoIwo9cFUFNs8FACsyvxgdc/2+VvzZsWXKjUo8xGEnibk
40udK2ZroU1yMK8OBXtQgFKivj1O7UmWPhG772271NcqpKfo7WbyMzeVrNNVBrMp33BRybhTnstS
ggNGNW/z//Y1OVtbYltnFftv7jd0Tf0ajzd4YAVw8fbc3G5fvwjKHWyPydSgd1XWf23AHZ5SCYeV
bY86XZZeJCai+mUuAiaHxRH9KUf5Dg+l+D+Srx9keO6cUO129ma6w/lluSlR48lmgkw1HKRTowQO
qBdydBvsAkXmF41QPy7TyZ1P2odDFeMk7TR4fywaLT5q2Yn3JRnt930r/0i4CTN/2KDOae4ECrQw
mMr0LHYwTYK3hPOTonvz6ro/2gArix3e3QYJRWCEEz6YrDXN0cyGVlIhFv6YMQyF4Wb36I8Vhpzw
wdsEI2G7B3YvF28kGV1yKoC4cu0gQQHeH2lupaHagUK++w/8OvkA+ZfCOJS/WWK6dJx+K9etvmc8
vrRteWMKsTC7L9ZcqJgRris4kyAR8tG26p/AglW1t68J4kKrGQ2g6Vrr0dwe2xiuOLFgdqo8pJs8
Jvle3YkV0zHXlp5/TbuFGyimJOtttrwZFkKcHVK/eJEOMuxYZgKGOvsy1jRonAfVcJqI8DogSZJ+
TR4ws7icLV3KM2tljyOVGMd6tPxrz8VD8IuC82qocLtbTco+bM9HDKttY2NPqfQXep/Ti2LmJStt
2hEKcE4biGwkr8F21r+tdUabtPgNBKvtbkgrL1sDj2+v6LhqV1fsjd+jGEwUlrLltD4ZyVYhOumI
IHEHBQrB/QfhTYynYcM31sJqM9FtvipEHvbrBWIdY8QuZ+l/47jKx//K/P651Fl+LX9FZ2Uae/bc
aKXZtCVVZqYGkBAFc8BzEnnSr1HtfcyXx67W599WAVYNu7PjiddCroGuH/7SACjfhztiYWnxiShx
ZtI9yt5vv6wrscnXUz/NI8F9HVnUJj2dqosFJlm0JFwna6DIEzduuCxtKBQ9GFOdHSTungNeQHC6
ldDAE2AGLxVRraY8+YUtT13yGLdf/mKybX+/HaeLD2mOAJZWytjMTFIPGlh1S6Dezut7zjHJgxBG
uhgfjAntHI7gy+yQc7VaB/X+RHkFEDNy17/jxUne0NtYTr0/W8tlDdif1nBwaFoyGuctAg6fOc9k
4zAUFTAgByDwYclrQcPGsOXj0B7Jh2OvmgP2kbpzsxd6bQfds8daa7gJXKvRu9v5BAIFdCFWbcpu
Ut9W7aR3owDz8AkJaSftWw8WX0eShkTfwyUpp1jNP0nhEZ6t7PDHb7dbB6kUTBoz17n7gPT6slWK
OpAZehqWAaBNJmomYIIpxSiEkBZLYMQdyhIxgYBWqP2MHw+Y11ZOpnuB/B2xUmCQ6gzFndJzZxL5
YLZVKM8+/dzN594ErQ8Z4SfLInAKYr0f1XGjbR+QIEwBajah+nLRC3i4SDOLKoytpbfJglk6wqm7
HKn3ZpxMvHeSrDIBjr9+/iDVjAtPbfFyHCymXI4V/SnVyRnPfWk9th28CilfRxhXLCgx5GMwL+e5
dn4CNSMBVkEwSBiD2WsDgDFMdY6y9bxmJqgZR2FwD3S8xd/o8daimDGX0AYvPyFA/9Hri6nmmA97
hMBwh5RentB8pa276y/dLNnLFUNLds4Lrsfr2apffPqhLXLXMKqeaCTQ7gcZf2L+j9Ey55EqWtcm
Y/G1lC9c/E7TNRy/HH51yCOirouv3IR26qMg1MOiyD4ax0ochqWXcFS8lOLN5cv6G8Lqa7JmYvNJ
zzdP8yEDIkk0Zp5zXzXiH9kh6ntQ62n9/JhExJfu1FCJl7YqxgYfTqMitldeCpMJbFmqrbUq1vQd
BZKmMwpw0/pPcqosgRkAt0fJP4phFzJj7himJg35EMVmII5TXc7g+hAlAlwqDT4FcBI4aQ83HQO5
Ukzx7ZMrtFi19ejhDW//+dNxlvArtBvF/WbKTiOVBXvbOWT0okdkOic/WvDbEiRicoUPeczkThaT
lw9Au0ffVCDklG9+Ou/qr8flHTuywZo1UI8pXnB2Ur4XTL7RArgB9iecoQavgagmNqiepUhTOgOL
H4wZhR3Iw4bIfnwY1O4/ZD1AqZhAzcTnfE839lCmMI8itm8fYNThAM/AQ/5roFMOU5TsGR2PczjR
uvs6cx04jdwR3VEwMgDHneFeoqPHc3nY5dbUcoO8e8lPXLLRS+zFBJvAbX+LWugs8zoszpMS142S
SEdnG9UzW8AiBfYlXl5n5zBUsQ62wOp+MDywl2Q8NGotPi16ElbUqQKFVcWkbJabvjHZMdfeJbfL
dB22oWh/wmUCVnBTxP95Qs354p8k60SrLrhV5IuBluZpyOmGUBpFwVs9bLBG8PbRRfokkOkEGWXP
7Z2FYtwoEV1+w5NQfuw25B04PFfmb8JzpGjQPIBxjfy57wrZYbQfQ0wKXivbBjjTZmvFbgjZYcO9
AjpmyX7TPAXBuMJic69GbmlfPtYIKXQbxX3dAtZ0WOuOEvH2yw5CVN9BDcMcTEC25mR6v6UZLTPf
7Kcm1V4N2ySxuTjTvL6u3F9bhdoaFjnzn+/ZekxUtILuIpWQmNNvflSOjfZkh/XDOX9ZqYCV2nue
1NwDmQ+uCZNF/cKH44R69bibjrW1Ua+DMRP30ZnsiJcPCnz1Zk8wRgcUElG82DlqtPAyBk4eN/2z
BAb/75tU9wTc2UvxPUszYkUJA73UXPubbryDPW48S8wjns12Dluqpyp+Bn0Zi17I5JDXnew2oSFf
fyGPDPUf2MR+c4NtCKAqQyH1QInBW6qNrYqUFjDGVyG5WslVPJodrqPPRNB4/KOfSgr3SquzhejR
T821dbB0d0xGfdt+dm3+m8xwWLC7NNCDKnqqxCwIjAsG+P/IhVfN2jlG3yrSO+0VOtNDLvadAKaF
96u4y50ccjuGSbZtJGXCUOl7NpmoeL532LyKmrpVGtMsqIseySNIzCcv2H7/suzb4LzVO/KRa2r6
r/Zbx3dvhoJch4LszThjryxttbniGnv+8fBTPgENE9Ndf0SPHgMT8BtFutoeIrsn5vYocsHhs/gA
SvYDWkcHpqfT1i9RbPInnHqanGq13h/pWLd8RPd241Ghv+iJ67Rei5AN1fWxyyRF7pIFnl2re+Je
jzsTSWhQfOQDAjVXrNjdv9e7LodJVW5BLhAFrppQwMdjSjSdib+cs0t65zT+VbNX6/nP9MEFM10o
NPpiu9D9a8bG52Ng9ENO13ZewHJfrgZW9dkc+b3X+Jp5P+McpePtZIWW0sfe8wGXFlujF/w+u2e9
YYlRGLThLaiW+yQ0e9STWF+ZDOtJgxAkDHDJaLG5QthNMLdPsObq21WHPg1xSK6zBzDYzugIfsUN
dcZGJt6o9MPcuM4+QRnAoorufCSR1qS5BK/D1Dycd48z4SyHJfrvPfL7r+zdl5jR1j8nN7RL/iQB
nX3Ze5Elk+kLcQSYjotxOA6aeduFgEZiuE7FEBDFQf1ymTyJEOpz1WUAJLhPGsKNzqgaGhOiF9aR
XRorfH2n9k33ZC0+xGNNnxXpfjDMysoEsABW5VPcUhyOhRvnQTF+SbRXEiEvJBhMWKbqumN3pUHF
CsH/f6EYfZ2CSNwVCkwdTVupbOFBC/4BeLvG0TgJrZ2kFbjjT3J7OTUYdLKMpguZxWBikz20+4uZ
Yg+d4wQbxjCYiRBJmS5aG/XkwXrQBn7VdQK5+Zfz995I9PX6jfohm2CgtNuJbKljDXiMjQNgPcc4
XpiPFX/1TkWGUQmFDgVOsDd4+A4zRU8ZK3tQBTzARzVCZnagsL0rwMSkCROSi65qrg8dwlUVR2lb
BmsSbhO4yCgI/T5sNZ//JvhjQg6VtSGJO8RCsiVplbe2TC+/w16JhHxV0K3GGH2TzyWGE9dGj0zO
phSdCVaNGHuvcsqwqGMrbeujPTEL3eiY+TsVUySu91NpOb8VDNVRG0gvTdFnkoQ4CJVcJYJFGaHy
GUEfygXv87I6x9JRXTJqGChZRzE4fiRvNlSLglB9cpc3QMqfwzOXardeHLI/tYHebhoelgSfy2ID
HH5q5QTxGx/4/f2OH4zFRvF64ghmU9zSv7+Fb5GsolKkkhF/82D+VUc3WeJzIu/mspYvXRfen/uX
h4ibAes1hHLZv5fVtCAV2baOk1zxsK3bpfta3pxFN4fei9RF8g9zu8L/0biAFkngaSRZ4h8Q/lde
H3rtXT3SRipZ+PR+h2D9NgV0+aVCD5kRCxPGU3r8ueWqxtQOGv5gLRoNGp6Oufe4kYe5O9A2Tbkn
fO8NSUqN1fGjyPN+EjAMbvChZAp12TMiSvoWGoykdjIVamc+s7YRysK77C9hNEmgU9ov80mXYYew
l1iIm7bbQDb7pT4/lCEXLle40/QSsNa06rJNhwqkW0HT552Yf3BTyvfE904XID6QUgaEZdynmuYx
EZ2apbKcuGPhjb1mKEu9TolVa1o2FZjmDXpE91Jf/sVx2r4taCB0InfIikGsuZ9Gf1o8b2l0HS4J
nKAjNgJP7XOPG2Z06dYPJyC7lIYupsmq8fQ6Xh7XsTzeCBsaVGUbIohOLzvLrm9ur+hRTRv+VfRa
848IM0TXuI0X3IoZLdryY29B4ab/9yCgFx6GyvbRgt9n+2yadDZy9hxw86nB7OeGruT5VQOYeBee
hymfkWpoMsU+3Xukf7w3B6tN1Q1lExrVIqnRlEP1Wd0/5DAOZtiibu92YxBj0WQd56Tb3p9D/jam
fb4JEtQ1BBp7wi8M2FkpVRvJ4d+2wpBv2fF/R+xR7EzHDQci6awT3Pf4JVjVCIaps1Fgkc69jwv7
8vbxu8CRRwUBd6ULIBlrPc84k4Ji0CRdkcXgr5yemQqJF81OGkC1LuHTquXzgQg1EK0+5VDwV5G6
hYSsBkcpJpWaXVK+4pao+XpVOB7ho1mACq2J5dOrNUVUOBuaLblG8Mic7pbN3uJl3kmOwFvpG56y
gNTdDzZGzTV0FlkKEYM294MVyqnT+QL+OAVmXPpYW2V8TtgTbvLm9m8x5ytU1WwORbviCq50TI5r
BGGfobXPKaPDtPPbLdbQ/5c4owPOBxZPwMFSgawlZGmsC6lof6DbpdoPXQq6TBa1tARa8ay4LjEU
gpdUNzKrhiI7zLEaCODb86UI6dsMtxvueL9nomnzcBKAuwEhHHlmvfp1iTX4ksuUmwwI9nez8ARA
wMKxwCzrJySHmKz+d+N18JcL5rdZdGoMzCjPYhns0HeXFJzuur7YCRtRT2gOeKPVeeHmXGECIJR4
X9/dtpn4w095zcaRcMYCRcpQ+WnjiiXTeEGjGIfbuxjB0C47FB2OKiLxBDtMyqW7+wmkjhvxUAT1
zRZ9SLSSsBIi5cRplB/3v1hAa0FATpUuC4D+sak1KUl9yrNhflJuLWg0kaUOo1W0sXsAjsLpTTqx
km9hNrrUySW/ieuiXsgw+mEEEQ9uj19B0g4f6/CKmrMv9taj2s4eKg98x/M5AnOEqHCa3Pls1i76
4gszO9HDHnPJf5naAqmlGCHJlybniV8qX4sSygq3uq236qx/04pYzxg6kj7XDQi6H+x0u87Vhb04
mLjR0d+W9YTaMw/iFmAtzn9Gs0jQwwYtz+wBYZPeimWRzQgsTGl8Ry4/yuZRAL5qAx5LjSCJsS0+
shQ48Zh0Ukw3Uu+/SQwXWiQepmNk1Uut6w1p31qsigOejOGqUtOuEiw4rXIl6t7nx25z+gSPHhjQ
/LFEdc96H/Q2j0DA4xsgvRz63TC6UPbDlgDFtz3r5CL2OFmEX2WH908wxl/22Jquzw1etc2328gF
UOvTAwNJSryqEqKY6OXcpTPSdhCbjyjJOhEi94WyDLc04pRza6iN7Bwargk+auat8h9btySdLOd3
f8vBCeSBwEdoIa1ROyKo30qTBr+FHRIRJzox+mPXWd5Bs0Xii8AdiRSRzJYc8U14Wij9pv0E+hqY
mbLU2oMNdXqdawZ66z99ilvOA9Ch3cbnE0Lbj3a8MMSyPXHKIp/5E4uLMbMm6xqlh9TfrnS+3/Kr
Nrru7wUOGSKPb7lY/Q6HE2Y/QPHDoNYCDAM34Sz4GMPHJZ760dsdLARXvUfh934XXyLMWUo8GZCj
7hKwq+etIpFHo2kbFc3coFW8CmT9ajeUb/Jy6K5jOHjUhShdy9JGtmp545C9o0AZDeQDkfN7nLyv
B6g1GYD0ZogCAbCR+sqZ7R+f/RXGrAlWEOQ5FdvUsouKuKAZm88SgH4Bzis6o4NhSfOfSm4rWLYE
QgQdVPMuFAwImlRdLd4vudPQR/tyR8tRD4G1jaNCgAuqazJAtMSTjjiooNYasOgqXv87ktt1Ix65
P82xy8Kn8B00KizlXTJCDWhjoqTX+dvaXygElWkU+085vhE7emWZZY+2kokHVAOm/2jTXQwN4yCR
hBOKaWH/7XTF4GgwGkUsQjYVikO/4jkHH3OJedEB00F8PC/lcR6JzjUBSg/+TlqpBRFz8D8Axb5o
ejVSqj1TTZz1PUoNcGFcqpf/898xfBDdARKdOcHgw9Fs34ogowkXmXiAmY13VvgFFtLEKxYsW9kq
pKUQW/oTJChU+pWVIbVKHxc64hSSMJlZUggkXJy5yhb0XEg5s5KXt1Mvvwm4ZxwJoBDPN1XfeWT9
P4wJanvfQs2+8qgPPvLW3V5fRoG0Nn6oYL80tofMwyij15UrD+wOYUri+78fjyX7dYem7z8eqh6a
9Eowg+RPXajAbBAUr7R86An+TyxchJPV4hQnQX8Jw4F9k8lnVPhlBlMYdRI+mfuJ+jqfPn5LoUql
AVqvb963HypYxTCSC9XqDcjy1kCmIlAZx+a7VmStBi1nKnX/MaDpOyB5NI57a5S7J1H1FN20dKrQ
tLGwk1czChSlFPeyloky2byFiFXtxuhgZaM3EcXq9i21xp7UgYgU6v6jXCAKFhA0gy5D3kSReHhh
ifDjvRWDP6LrEsbERYVr6ZZUCJ4z9/nXSaDNSsxjoqpLchJCHEscUetrCpxoCa8dS3je9659PDlw
DGPrPcMCHhgjyjo/2HFJDkhfJ7C3TIIgaV66vegC5Os7eEOJWWF1GMSlgvQPmzuDU3JZuU9NsdB3
C/TJZc3GfhH0QV0nWCbgKEduaT4mC8H4Mu9NT0nsYFx0SR3w2ZoiS7u8UU77YHtNKYuyCYp6UOTH
W/mQCvVqSq7c8Yf3Sbb3vlEIhazIUdFN9xFY386v/uGS7LOfnPLYEgr6uu698hp5MlfrB1URDts4
/U1b07hAVTmG8f/nhZH8L3gEq4o/eIxF8HoS2H23TyRxMbXJo+92U0ZHLUL6WROyrl+SY2TapOcF
jBBh/FHQLnNMFHsrabpTERnx37Mnq4KH272uqGrZH0BArtF15byJeD3LtCdC5/pvJvSOk3D8H5CE
S+0P8tQnQhhFHP4LJli5NdW5fFu4gWLEeQUeMSpvjWx1vnduE+dyx4tdBFZinXvahJYUggCbe1b7
E+soDlhDhn9wk+BKuszpqmo7n8qmVsKiOOi71biYkvwW2yYfrgevL4iLZ5EbFoEyBO6mI9EuwS/A
TnE+Uo+/qLbZn/y8ydeTd4m1a9jA1rIx5aUmDGUFpI4LD3qru8bTmxtLYgp1iJF/oqD3g6317Q3R
dC0bshIupwoXOt33Lryk3BcBcP+GQlXTjmLUwgldTSJJSJkqmnCMKgk3azGbvvkfIDP3HW0x7LtF
cNCM6SDQLj2hNLx2Am0Yryqpa2/+mCGSjbjbgYLmBlQ3aJO3YFn2c3oa4tiCGrdkHGBq7LaJ0Xal
Z2DEHo1notPsqR79/zVCFulJke+UXEDZVb2It6atjAff1buJW1jMI8BhLPzFk+0DZp4TlVDDdZRT
/O/q7B2zuPZqgxJqXXFGDDj24OaakFkZ6BMboXSO+JTd4WbGrtWIL05uZt6mYf3G/TiuwkUBPYfM
vDAn81mylaXq/vTqbD7tthcUQC33uZNHjqmqsc69SxbR0zK5fR9P3WJX3dec4e26rCDaRHSXUBl8
MW6wKbreMIKBMv1lvpGUYADO/rOQXbaUATSNXH+yaXgY3dU1R3uIyVF79969rz1vlG231GStLDiG
bSxR0k4zuBfdzDJgc5B6kHb6I4yUxBy5kZbXVK4m/72IUrBWYnjbiEihhY+4BfgV9LLa+1bcVGqu
+YDyAk/9ofeQh8RawMzPnaO2e4NCvmurh0mfN1sLvfWNnMliwujN9d66Knw+UydoBPnQxQom49+T
nDaOGxxsHcB0E8GAmRCCIVEK3xaddEZ/H12xt+t/bbPWRxKyccEY27kAyc7pXU1cpGKSlLqllvts
ffMct4xoNj+9OT+/1GRhCR7aqC6qtiPQcij92mUDvb1QUnZxmLwsbFgNAZgpd9BsGsOumPfAqLAh
9JOLaLAD3yBRDLE3aAEbrvAn6FjaudqZM/o+wTjd5jqpDD3q7/oM2Vc8y04ORhdTO7c4hGpCd4pB
5WePEmIJXlECvJIwTkw4DsZEH+t3MUzd7Dghcrbmd/HmqfPiagdD52Ql0R31usFT/BWipWY98qHc
7901eF3qebhBbaW+tgCXi6VVQjv4GMRBkYDfruJSJHNraBo1tw5N/8tOelkVmdq+R9aZx0p1Gemm
2YbXEXmWYsSF/Fc7jvH67mrpoqm8ezO4A86cRGJxndh5mUgUehdoqNwj8clFgvIym/Km0BmscnxY
cjHcCvu+sMqKlpSRfLSuYE74OBdwCrUTCEBOOZvZgC1nGdjeHbtGcqh1cxY6xGKc0xPJBm6FPRF6
2h+lsT0YyStfutum5ttPgqMxeHAP5ABJEAqf7s146Tpaa0M6HqhzsD7Dm2aje2rjBSTFK89fUq/m
KC7g3I8ToGcQD9Q1csdIXiloX2dLFH3Kr1UiLIlusf2wbZfeMu0TyqTLT2kl3uPlSgvUXYAKFgyc
P0zp9o40LOeyXCu/Le4F3i69h43fpTIZ6v0FcVN6AQq+R/dei66mDYHYGE6Xfh4NoELY/KUsK6QO
vTBcn1t6mYpXWooHjASqlODa8xtpQ+6MNoYTzvGrqAA26k8aO+B38kDuTAhU5MlT6YWl2acved55
bwgiqNIQHekcKOW6/Z+pgyMpLskC+cZKgk007ve4qG9xyyInyj/9zI07lqT+37RdI0EfhO4DYHzi
v2U7dBoRJpZMkZWMx2A/yYX6OkNH31YeT92mFJ+0WB4u6UcCaOzjAtp6Fi/qGswOSXw6yWPhKm6d
tudpl0rGLGyze2kfjCg8SgOYnBhMDt/h5+voWCUVR5y2kvLrk/P8hPlRl11HW+S1uKcg/TRR6930
Ts/Im2Dyi0ItCXYRby03YZM/T+hv/LOhYX91AKHYdLNs9zpGn+bjwLKV811Zj3pRBWWeqiHymGd6
5Xp3CvJoFKpJ+IpW68/ZLTIhJA/PqGVQ4+0ZgTG9MrfjUqXTkmEKDq8VMkARq2LZYemdmhTUGypX
Ul4ZEZq3nYcqxzOnprZzcNpM949luC6gamXqqShsO1AqxNTD7R5XexjisZWmBOKQ1ZUyGXgiq9uU
FsKnGYJnxFLOrkYpJecafZ/hkGxu4Kw8E2LSabP3W6weSAwKDTzCZNoFDIQt1wnIZ30a7WcK8+K2
IfgJ1qWM45HmnDtSD43qBvd4Mh84MP/DYVuyx5GTFJ8GX2UagJ7GMqDsuQ2RYiOTaZI5/GO9kM5x
0/F1R5FwsKgdpkENA41lly5NcF7635nMAvQk8nL2N9BbM8sS8hqNo990VGdBCtEIbHMXnUXnMDa2
mf0IWpDUZhdXIPgp5dY+BylAM6oH7NIt4uJIqv+esBcOL2Kj5YFwGmemm/RNJQib9bv20BzAnocm
bOY0JxlytnKuUdujysjZWiw9qUZnUmDE4KabHemU5aZtKHtkqhBoZg1ObBKdoPIqJ3oD27Wdtw2b
tqceuUsDivpRLoJNidWgg4MuhWoK/9bVJsqY63tXKtkJ4ebM6+XZ/HlkQogz/HvWXF4i+RrDq4TN
7QSk3P2UQTUrpHrHX/A/AtsNF60NgauUV1bSMNtqOZ8sKc/8H8EDoLBvM+rsSoB2JdlPUTuLXYqH
no542CY9EeYWxq44/bLa1m9/1jj3QUAXSuqJKQkAW/cOzSTPadw+6ajiVU7HXwCz4tFqpZT9gKax
KypetUlTOQDqvyVJ21QXTQ4VxzUs1AFR5F/MJmup1Aq3Sk7bSuO01gV9TK3kydXyud2uaYwjcmxH
V84pnUzRs5YN4ympdEebX8TPgccvx0b3W7293UbMkFSZuNa4DFHv+10eu9YbUmA4pZrboRy/dLRg
sMW8OSfoLp/Xw58u7ri0a6q42zuoLQ2ZMRR4Ri990U+4nuhvP94W1dH6H0+lU4gAB5lbVA8sVkeK
V3eedwoGD/EU89ggSOEOMXccLgQoVjw+oxjUz+IY8ZDrYvwT7zVLHydQEPBo1jrC9AvY2s6qu9Op
PzcBfsVifCXUiWF3gf2fqiSaK3alvJXTLGQzLQh5VuvXuAdSL+4jV9IfCAXoazokt3ohOfKV+71C
LGC305p+wO4jGiNnws9osBzyFiyFWiFdA2xwjQiNGbA2NzbalK/5nrHSAzOo3bj1axWuRuxA6bD+
PU+dqdcNvGoKGIh7KjJm75d5eJLu9N1+wR5lgOlFQ7LM/oUBD3d94DzZYmuW0oY9fhojxs7KtCUk
GWoTWFqkHZRDWVXNkad9aFbnVb7KDvwI5Mrr9xRlJt3IfeOVRw4QCyc23nSGSW5ZoTw1sVs9WAEb
9PJzP20WbmnPUjZvgIuIAghE7wOFbZgIwcz8uh+EMIW6R0gbtXt47nIvX6BRs9ol3QvHZeGcTw3k
H/YBb9FrcLGqK3qM3UyvXYAkBYzDE67zsanqcaBm3McDlXtq3RV/qgHVqJDm2CxnW0MNL7ipR2oq
Sf24ffupdek3uOo07tQYP7If5MT7YnIQKEfG3vrJerwsLa1no8MGKcx0SK8Ab+zwOWTytwbN8XmK
q/0vuJxgHCH6hzk0XmHzft2trSJeH4MWsCc2WiLFRil+tneSuX1q/klwg09d/9hc6UDCSkNANVJV
eTHIH6Xrda+hoGuuEe3hvwJFjhUywo4R6ArXiRcsqNlnQh2ddPUVEZOWsBQ9Aif4k7xTuQLKn675
x1iorVjlwgDgharEuhLoatuROis3VqkiVtvfFwh7IpkBt4AF3vuOihO6C45DbZuV3m2tHst1VrfY
FrtxKbN6AkMWBNd17JrQiNbHIuX5su3WLjqtE88CWi6mr/EChJKwqN8JOtW9qx39mj+Ut6uIZb7Y
q82ziI6KxzWbbmTODXMf77EMFJKW+j3BDGeZmRyizaDqYwRjhdBjwywN7rx0d1fNZj5NB9SX45P4
Pi3+pASVf5OetjdhmEtbAnC8ZZQHbzAiLHF/u2dQsEe1Db7mG592rbCkRut/KIBWBjdC87KuXsbP
/uyxIdIgsRIIS1We+aLTe+sxff2vKxEvAp3lf2K3YB6l/3YkHQfW35BtcuoBYvgs4QI3/NTyqKzD
mgrGOqjcMiyEQMs1LQbOV/mnvCWmOk45moH3lvI2m63Xch5rU5I9WmWZcmMDZSLKB1zb/eqpwEl9
Et1uwZhRUfNWAkOcRcUXH072P3vjVb8C68AZ6YnX0BTvbwDpJNtis5G7Y3Z2h4Put0cKKnEqsDap
TKdCVhr17R3hXISNadnbZoD7yu/tHDL9Cd22v9V58G4XriRjOVx+E7l8S592E5gdnH1EmuqnAOob
/F7iQYZraux2o/NhzTHZWMMupLjWyv/vGuoj04s19vUQ4VZe3SqWpxOFqNDzOzRM3BeZyGzMPfra
QpQtMAaH6hvgc/sQHuVu7HN2mA4iTkwiMsjtnancTgUhgvPblkGY/hlVXz23ExfoZEG63Iq2fQqa
8qqrSTWu+PdBH0HoLlguX6o+vyPB7HXQm/ZYhPX89jOdNwdH171wr9oLFdCtC5Kv05x5zE3wu8JN
3ZLpfyM5BqIee1CLFk0y7Ro42Y70gDyvfZK7KxzmJ6lp7qrcRF15O3lY588AVbOYwKkinebUCxLC
JWUG3fCI7Pu1btvuiGWMDkD0oDIi0pa9d6LahWtcE1XcFE8Z82uur24aXWpIIaC/lF1zGGFAqhlo
XEAzAtI7xWmIitnIJu1AFtYmBiebc8Bz9XwYVRcmBDDD64Ww4cH5DSSp7drGJogMZxdj6QEZE8KH
W8xIaVyGf/2o/YOvkfjDeIIVzFvbTT90Cjm2Qqg0d6UufSZnFCzoU6FjrCEdiHHQFlWIj67hrK9Q
jiGYAXSYaX/FyXflZkNXzEePFYOLaJDZA5RDTlsQS2UX642DtJbBfFYVu1/krSow6Ow+QGpOZF5P
tJNA2lEpL8/ePkPzT8MHfcRXtOg+ML3gbIMZN0mGVovx/Jh2ug8r54PBOSSaKR+VnHGBHvQ/v6/7
yAGkm4FbyAjvPozM5fzPZVu66A4Y3qRapVqtjyGnh4fiDDJo9X4UwTwsxUS7IsEhkQ5KFCYpo53S
OpyoQoAY8TFZjiQ3BxJyLOBjcZk11itdE9V6td6haUjSoEjtCAX1DT1O2/IkvSLTxKt+zvyfVrQE
TXdCANDHEQaBbr261rXFXvWUk82hgbx6B5pjhhaOYyx3esN5sQAwkYhXyZF/EuZ6chpMQvESxtsh
v797DV0Srz2z6m7+mXNH3dUUqrBaDrkCLa+qho9Za5kBn12GPWWos3ylrAil/RI9DhaMaHr/ME8g
iC0Un7Bh8MJ96CxsLJocmZqysdZc0HqRy7GpBj4zmvuVI3N3YaYsFUYDggsdw6WsHhpARe+Ak9Sj
TE8Sc7JHyk7OrrGONcQi+eUINDKH6k7sPLdl2z/7T9rcAadDvWJ3+wYaX5P4oNlDvTiNbVy2zIvL
kOeegIOmMnqOt+7HqWEBqwb5wTOqxXm4uo7JMhGZ40Egqa7tP6elv9itazOq8a8tRmOXPTsuzh0T
w6rxSuTRxwIj8Y5b49mOdaEOyV1vMMF262oWKdZ4XO4CNQ9HHMvYkQyVBGG43hizsI/gmurbq8w0
+f+aOZAg4pw6U8vUWLazKrF6lTrb7uOc2AZlbJAp430WmApVid17FiUDtPhNcDktudls1NkDaNrm
UCsdfTygGgmG02FrtJIfJ+Z7yBqepvAOab6zVM0HP4wP0fVBnr2AevST9/UPGbdxv1sI96IeHoDo
zjBpGbzdst+xu9Wdt0JT1RgtQ8G+Skx/tMoBQRHmI7IMoP2EQ4Q/313ZX4zEKGLLrww0+l/2Hkys
0f2foP9OpfVznff9VVpxxgHRYNYtfD5uoR9b0O48FzKkezQPI6zfXJbIol4vYgOTUwxHzTREEV/M
6qnK22tB8Du6muKqjg3n7PIxc9OhC/cGO4kjrZNTHL8YJen6KcQSuS29AtDwpCpgKf/i5rPYb6Lv
qRlGXFiLYXqKOX1cMqpY5cQP7Feom4Vo50ria0Mmng+OERPwLSoAUCmj48Xk9kHeSAj2ASasLxU1
iFWVatNbnLM2QVMGtDsf7FItsF471k7Ha/T0rEB/3jmpRVa8Q2GQCYxOMVEXrT5YpPPAmsaw2S1L
wLklEoz+ZAGB8ZgQmppv+0QwLkUjrVq+jAtjdymAVoQx1hDtWc+rGOvm/xlus+kOaHYgcQFHArCN
HwcqRCopuYjVK6mP82HEE0kLR0jze7eZ9k0wD60WWtyMuvH3j8Ccly9QTyBUY1dkwWyTh0D5v5A1
zFapC30ObVy2sFnlE43bUhs03SrdpF6fHICZFTb8d1+RcYbO/EKgYPFNN9Kg5EOKsRuCr6IM4Wm2
n18W1ZieARHSkL4tW9hESJJ0r57nlux3KlBBO0jpTdZSTy6xwLIObvxWe/1nazrYRb5E7GHxEiI7
48dRmgUriWxDo+WY6B4v+JzL5QlvQp/HBGoJf2cJoih8PHsf8+YJCSGrI4ElCMYsTfNsRHLxDkWb
i/oOOSHhsGV4TYopgtyucZe/JcXODuMns8KIv9Wt/nbr5dhaYgCycXaaetYi/pv2B41oy6tqaK85
E5wtmGMf6lIsO199PZZv/f5AFvJ1IEwyFGaUm6baQzsBA2M1EvdvF3kex0u4qlGYROWGptzSUe0G
G6qAEXVqOgvktiKzvKpryIyRTaWvxeE+bUmrhnmIKiq6w6R6TaaVtEVICCOaUMQV66C37+Ur22wu
nX9vY4tLxL2MMdrSclnXQMxI9d65DCyr9CDqt7LFDQtbl0R2Bo4Osi+u9ifO8DwkuExMZcCsz/DI
OOiAs2DFRMTGKLpMGfkdagrys+SPga7X82Gi5ttnX8sfdVlYB5tquBupQfxeNyP8rKnr5Kje1Wrh
NM9dQrJCzqjp8uf7OT6qLlsqnoyzkDupi9icxRlNzOvUUTR/gXo2fL+qQwx7H9s8OJVOzIbBW9Q2
zTIw+y2Wn9OWBPmoJjpBr9yGt+Q3t+Q4meCDDwSkWGnjOZMBZwHqhmSg9uCOOh7VMWFwymamyxXj
FLT6qYAynedPzAp+njuJRLVeq2vE47hZLf6bBk7t3rFKiJ06ATSmZ4cHb+Vcqz6GYEII/Bp5hjYd
lA+35CBrC2lzvQEXimLONsfysnnJ4BtjuQFW4o4Tdh8jefik5krG8f5VNAVG9xw/i4Gk4OzsvYs/
NfvcsZkKRDkZunXC+vnp7WhztDv/OSq9CrEM2oyNsZ1zbUibYAMlfXELKItqNe+qeyzGcpICwCxU
jLPapg1rxGBnb1XFLF3gjXM9hty5SNJjuk+gtbAqEhfbtL7bkISH56+6kyNRfpLS7IL3fdId0EQm
wB7cEdG5JLx+EAVtAccUc7fSmCAtpCvoy55DXU1nqP2wjE51dTJrS6Un32VZ0mZ1QtjPUHOd+GIQ
2QU+lUm0nDrKLhkNGdfQggBQKztPbnMa4DFJPmrL5pkDccxamV8MJqFosxNHJeiiJ9DLSKXoHx3D
CUNUWlydTFqLf8Bh7mNwR3H1a1ttBJr1dXAGY7HVGMqywRQHTHf/DfT6tiKQEAYqQoHpxyo7HGhh
LhhL3XlC6l5saLiYbA5mvdco9C2CExBzGAInsQMG0lFuH/57lVH3SpEuwfjhObLM3PNUn0IacqBs
sexbPSOeGFT8WsL5BsM33gRXeBhxInSAMRx+RJ2Rw+W6BDNCwKUi+j78NHm1lpE3YHQdBreJ8u3N
0UslNyiuUPUaz6NXSUNvYLs0hLk0DFHsz6R1qKu2O+d3ZoQVlsbEBxtAtA84mROWiyM/dKJSBza7
6zPP3xnhWCxApIs+LjIRLLIR4x64gsrY0GIpKqu7MJVXipbZ0zzBEOWsGLwVOZK4TCmlD0XhaMOn
R+GsfTPJWS0cjfXX3lOoAJs59xiEDB+5P/94un1iazu3yqDdEQO2Nlq1la/rZyKExKFDIGb47XIi
jSGJq492vV+iCUmDR+ixYzJvbwFZ8gFly2EiLtAP5Sygv9QhIxKAU8ztEEY9QF54nqd0mJmE3256
UmUJaobRdC0nG8moyOZoxoe/LDWZKk43SUeh3s18pBly3RveYAjyO5kCPIAn0SSY6kp4oImez4Tp
xAQguHaIweiDSVDfPsXwEkKEn64ZZOe7pOZhaIAK7xFd5OJzm7HvSXpP4dNW+97xQlVJnfKxxUwB
udLlY19vZoz4dIK8+3/LpdG/fWF6hzmmhllTt4SffA5VB/eDcmODgFv+8AAmi2COwndVulGmCbd8
f9D6eDODNKhRt9kuHft8pIG+NQTNpsftGwduVl9sGMiUk7kKzMXoIEewtQlKDqat2VQNwsAmT/NJ
17mDsSX0Gh8ClOCGoFlDEhdpM6yAsqYhFUx1j3Hga3nTRDEUspQFd6t8+UJmeSOyzCjWy6Qxu9rv
vGuNqmPNReWs4s7B4fzRatUnTTspiBQ2lrqnUNrRnyQaIXZR6WhsCjZ2ZWNuA4cpJ/oFGGLpOSW9
GjbCGmsEUKvba+CAQTEFKh3TnAYBT4iLbG5jBc1dM7wwOVADRtqNOVK6SMcc0Z6MuuzsM40pnEz8
2fxjZdKK0JGdw00+nq83tWf3OVLfTFfPkMXYxiIQKDVS/K5+i3J7cl2Kqr/ZTQC54gYP733TquW+
3gehITPTpdtQUBFy5W5Z1cJcmAcPbGv26HI408sNr91+eg07J8pPtLfoSJ4XmJtkH8/yTXvfBMDP
9QtIQ/i3XEDkQbigIWZluhOXWrzVvErnc5wkLleLUkEIshuz+eJlyg48dmq1LAluKsg5x5GXbses
BlXpBaxAJBlCIzkCtEjBlBPlB6Ze/nze0X/q19atD6+4m2Bzsrqo1fewlIkVjvgvV8HD8JTERCb/
yuRpimdWrUJYW60ngFkY53CZBfCT+oGI1Brd5/hMXbrSG5nG3Yk+SyTsjwHRqZM37L+YtqtAkYeq
MLO7saP/MP7x3vAFzbimFqpHvkINoFRwFVU3CmefFXlMOKb/RN41b0NrQAPX2qBh4d57uPzdTxPW
idkVmYTL/y5f44HCQErCywvDfUy7Ay3EKcGbulFIsDo9tMMDuuxPs0wYk7Q4oONYpAgzeu36/YTS
4Uy2aHEyrGZVD/Y/kNqXDBAyA7YQEcpUkeftSR09fluxEJmIATd/SHeVUkA5eUlwI1D/hHw6Vf+C
SdQXjJP3nx6pzW0spfptoRzJmN46/GBsXe61FNdc9UlyWps/tlhOq3qSlLiEHoMXuiZiUobjnX2W
wDYlPbHbTRrA/jvTwU45IXXhtQAq90Vuud7HAHrYWhN0R//TXDPvKTxE5Tnv4SdZsnl9TWz1w2ig
wgefTqKMoAmlVo0MyN/RFGKcXKxibADCu4Qlulwq0+l4pH+QvtUgkBXJv7FC399tzhlvagSJ5NMC
srNS8008VZ7qvQfQzeOeA+et3vz9+2e+Wh64u+QmbW+LdgWiKhrMLCVWEJKshz20kBHLHCu/70+d
JOKsrG3345B+wQ8D8DevjWljmIabUniUPVp5MxmTq/lVVf4dGDIwfJdEMv0PX64e+1CvZUcomQ2l
n/YNNr237lzwIwD4NaojccwxJKAxLg7UpTArC0SblJiAxnyB0P5kLYBocQu9D0Hgsyb6mZVat7sK
T7UNryKw0Soy2hz0L8kUDYZB/phLGHzmTEcjPYfM0hl6mOyx3KMMip+B+io836ZWCR2itEUklA/e
aaQh2kS1pye2xYadls+Pca+pq5TiEuLquMQPnA+VXS/5+NuwBI4Y44TO7qxG8x1xfEywcgWmdvoK
LLSJ1OcKgd9x2zhIloawZ3q2JCI8FC+3AKMbi2o8bvTy2CDe0tamxrjQlBQqUT1KgG45DhvEZ1U2
4ONe0W4QqYK9J2YFKjBXr3pOLMJIYtTpRDfjE7bl9q+H2vAF8nnZCCWEolMVkACgpTedAm3q5gDP
ClKHChn7/GOLjkn6J5aqZU0tIV4cliuE4f3ugLi8mHxj9mK21TFec3oBNfRdcgSoewksqDgyiqvL
EAWVyl8y6F6jUo86CsrJH6Pamd7x+Ltcj5wUQTUT0OT3OcZ0iy2FQR98zmoCi+nvPZC5tgDGLQ1r
aIF0kd9/8WwAmZXwLP0CRz3KiFHkcv1DiEZqAPG/3VHQTUkWgYenqYYFYvsLnmjTZJJng4+H5NdA
u548OkhHBGH51GyaX+Gr0oFprQW3UHSmh/i9liDfyYWXuTIJbuICSzN/8Hi6UKtKOG3pe/cFOOa1
bZsYjBulDPYxgG9NJ5ZqbLmPDf+CIJrULCptXn1b8HtEtqNnlqgy48U3qdVjzv5btv/kaVPBqnbk
oTHGrK+X6CpfRNJvHmmKM3VgirSjPzfmZb7H2RL6HVftAMu8nvfT62yXGqvocyd4K8Jb3WH4hQZT
KdKiUzh52fGPKzlhdNWYNYP/RUroZ6fSRpyZ09fj/5P+mVDkMqsgb2kf799Dssn/8/ZPOTmp1Xg5
vAITstOq9Fn8JsWjStSoE1r6lzJPL+yuwm5w0wpR82odPpLesYPfzxByTO7XTsPGaWby1MwnVz9f
71Gwu2kU2xey0k+LbD7Yywt32VNAvD0Cr6Nho+C+rMvoHl9J1J/HKmzyVow34t/mn18A1ZCA7l+n
OybWZsMMCtyTGMyqvawQ6mA4sDF6XpU/eaf14pMylf5IIxC18bNDja9j9HLXluSWLRH2ZKZtS9B1
7ujdc+f3BxB/H7Xe6HL/5ursRej3CnvP+tAlAiwlSx7w/I8qN/+YSJmR/Nml9hXWndqo8gbZQk8l
MlAZm1sZUmlhgzquI03EpcqJeSOFoPep0bGyH7MPoJL4MLrT7rgX2+uKmH+OTkLqKDOoNkQH6u4F
rsVoL3wDHrzViemd67wJNJTVLF3PZScWTyKrfWDJHGzE2NyKpV8D5VWfYT3drfJOINpqlsCBLEec
UzkA//qHxJAnMiifUAQxVEPVT8Lpb/QoQSVEs0q6TnXN4P1i0NfUkaTbUP4iEoaw07wapbFbd6YB
mGYYAqWU+M4RT2zJhCPxdFk+5i/xUgG1kDPjwwlhBx5oxncR5nqimJu7P7z+2ZrU4T6izavHYMr5
E2/kSxIG+R1rQsssiDT5AGqHyp9duh+xu9bg43vu4Z3U14Y3qyC4mMOOf0OvxaI7jlhC5FOfB9lW
TSDbdEzvbW8pgEuGA1rFTz8Rzk1ahCzwGdPXxsroS60iDmXs8P7r+rSyIIAUN8qTdrakGHKP4J8G
gxPXNg7KXhcsZYPJJBvBm+3JFDVlbyFq9iavOFu/1gqZyl5Xk3yYhaMRO+GVSVpuSbmqKyqbHWlU
DCTsrSlnmRxOSNcimfckplP7r5KjJrYh2+9qJgS/r0HbeuKbz1Re+WQr9VYbby2UDrjLOLAG1zAc
/qvy1iXuE9JKsMb/UxMmaYcC9IP3GahJlVkQjZEdq8qhb6UNka9KVr2zjEYGGT+xA45zXyuMuPHM
5sBgTZL+Dto8dv7aiPaMlufpF5fhqHv238xF0EiOKIJvYQDRAjLP/2F0nv0fZ+PiMwZKoTAyFo9T
ZG3swl8WV6qDQUTfjTq45BqPnnad86B8AA/0Iks2iFnV65YKOP2fsiivlXyLXeyKpjpgd2CD8BSB
BA9Grjy03C5uevpW0cma6H7u4TRJDUq7u2sdFVQBGiyr7lYCMLJ7vnOnhbszgOijS21465zIP3kb
SE4pYwUCJDd3SSSdfLm/jqFDA+KPAnPjlwZMOc8/Ivwq0USX9rgoLPWaTqEyH42tLqW2W94j7JSn
pxsAS6ufgIxwutt9H7oGrSuGLTWQTLHz6aZdiugTzkStyE64zyDa3fAl2MHF37L9fvrvnst7cHTg
Ga5EedxndaRstwzOrjjnagu1qOMxh06v9t1B2RWclXlo/3P8UjYEe7b3Cgf4Ypp7Yv2+yWlc5Esp
+H0hvsDxcwSTMiQmhOI+JsNqCvGMA7YelajkGLFgVttOPjx1tNPR8uheeOy/i6YRHe7FW+H9g43M
rld+Dsr1B3Gu3EC0lAWVm4yHI9kVnztfXJTtu0vats64rWz8ioQ7r8F5Wdy429oljKb/KaVI6GYp
CwJf1hYb8UjqL1K8oLVClIJ2Cta9mLD2QvQCQVz+HF8DyQHvKxjjWELY5EJtuExLxokjTHTzzrrH
IekwEmwTMvWHF0jWu0lpMQUTzKjOPfGfJO1zRZWVP0NCabLXE2p8d0o0LundA5YqiX/3OP/ZVbNx
XNF0Iwe+XOB2wSeLbKh4FJQCVn7ctRImxcUHaqEyjVFlsd+IXA3d54W70pmWfIcmQsVm180sQO30
eJCvZWdzjT0aOAMFr7m834IMPEEhONWsI2bcmbZBNdaNmy8Gr2hVl5c1UZ8AxGfvxsmOHzd7v2hH
zGNGqXS1SEoFX8AmSmRc5yarI8JJV3PjTxs/wHeqjfgkhCDf9w3NbJRizPVxo7CgnPoNat+Xjr5Q
pQU0pmtkoBFdcuFwrKjVW2IuZaCB9guq5pBvG+kSEz4MZ91JtLBMB0zJLwbuxWNFvj/wzry+8Jhl
OjinHhqEqD8XjHgR55lf92HZBnse9FRYI7HsDn80TZG2ZUISWySm/TMeWL84e1gtXuJ+Id3OL0Rv
cW0txoNWkevTPCtQTXAyoecwmDAdKqwVqwSqpx0C14YHhuuoqgdAGyV7k0F6RyGpxxWdyoo9l6gj
mfp/i/oi/UOCiJa6IszLu+vwrf+pO9XQB+C3mtEsXfLulGqZkHqsdVeE0rKXHAKK07ViQSdo2go/
frtN6h+BfqnZdNc2QrO2eAy5AQ9+qiaSt5UdzlZbv4FXjmziY8uHBbR7t1tww5MW7QDGprsxq/A6
Dhd13R3lLosHPXmbprx77nqpO29ywyZUPdSLY0FP4Z5bFLSMdXDIpNcUlE4/uGbhkVXyQV2q/0Sk
41CVav6CgBgotscSOwAvtdMFGVXvuw1U+8WZhTS1quTrxYv6tuue30he1sZ/mNae/XUExefgegNt
XrPG8uRRwwhVsNa51JNsG7a5+Rygmc5u/N/vu/Kgt8BKQUiC1J7CM2fEeTfXmY4LYncFWq316SW7
qKHk5X+apHF015hF17kyGkh51U5fLQN5oghPCcasZ9PUQ1T1aB3i4AHj7g9yhTvUOz3GYE7U/fNM
MFXoes/vzkc+JQHuqs7xPyGCAAIrOvRYix0/cq+JdxLWPwMhEz71qCZlGwQTFSpoOXvr2OCn4FBr
US+lV7Z/hW5nhJKIyxYvYG87Ffyok+zzF9jpRGTXNccQjklsfG8aLBKTzGOJAp45EHN0jAb9b2v8
jt8TZM8PW/LW1zXusAVnwypYmQpffHZNpfw1CgbSQnXcZ1v15WjgUNjm1GPJyODUQTkSSKFMTbQ+
qmIZNz5kJo80/j5eyuS2O50/7q/eNpgdfq3eS7rJR0GuA+YvPxldJfq5HNuApUSFMFYasaURUAO+
S3PrvUECEN6/LFHzSeKO0/HQCMGfnctuFSYueKHzaezDVJOELNuoHlfeupWfRD7n+z/T57A0KFLy
PPhC/ZIVN0USzc+9t6jY5zkXLT5ewxPgJDSFmYQ7ylPuyg9hkSHkGQVxSQxxsgBJhG9WbKsk8tmo
qwmsM2Hj8zwDK4MghUYGsa3SbE2apZice7DiGKw1EUqhJQXPPNRnaBQbVBUwWSqz/0TLdSSMBpzS
rjMQFS++E79RKGQ1H6Q4p9aRvieJWET7N6EO39osohOAU2pYKFzq8ml+LvPCXE6Bvhr1UuXKzI41
Qij2TLLuvFwgqOJwD+EEwZLhIvOvXBZIZ9mfpQfqThzAhh6LKr7gMn/FuATryKHf7Z8iIDCQzvyn
RsrzI+f8Zv2QICUaQb5m4VYX8ejEU7TJhif2f6cWbPWefF0RPEmzC1gmz4OmjckjN5s10JHsrUPo
LsXUP8Xe9WxbdA1ydOdIvlvHtdoB3GPhQBvkjrhvlpP4lmjA0F1LKFnSty0Bq9HX3/XTFtK2hHdC
sBPCtmfWLD5sPO/ts0QpVZNk/C15Eyb97327E0NuY/bhPKygP3LGCkJzxSC4zd3i9veH7L0JMKwr
JnUEJdIfOnjXjsfBDEiVBOFC8kvpMyXBIEZJGEd98HnHS0HP9pkmNPKRrnDNKWNM3sSO4+QSJH2s
NqS2wTTZ1s6tWzoJgR01v7nhHDmh80911ATLlrgxaQWzdCfLSdPh185wJxF2qTBdRFjTxnHW+fig
2D/ozFjG9ukGTyb6rcFU72nKxlbQbHT3rS57MfBQ5lgU+Fjday/8DuH+42mTDrQU8kGlYhX+JCQs
GeqJ9zJxe8beJHQp5//Mf/0bmevY+yfJ32xRYkt6nyzThi1F6KkUFVffLQ7/2XRNTAbJy0KNr0Bw
QJW0kFCHCVwau2REO8x+ZTrdOaOxAM9rnbxbqHn8RgEKTgAyg5TJirlIcVISmI2dDrsYK8n6VF5Z
rXjCCy4pkm9ebMgPlW8tzQPL/jiylVd7RAxiYkc+pPDBVmztxTdhZQfnI5qhjcKIo4WVRD1LOSJv
AxZeXKUtqHJF/S2B3Wq+LRKLx0vt/WpIgIhq242Pk/jZjQbrjPSEk1Qxvnybr4rcxx4Kd8FAli+o
q5q4Bm5JqCLOB7rfB9O6FjBZ9UbdZR70P/2M1lD5u67h1nn/y0O0MC3rWJvx3bua0IAa91rk5N9W
q7Khw+cHWJrgeZVUl8J2Om07uz3KQ83tj9SMtVoVe0S2rpqX8Jai6siIF5FBX8i0nPc5G4VcYZ0m
Nm3gfBfJIUhHrfIeNSeQq36Uv9mxGWdRsjUAMTdifJWoY3ndglBVuXnjItmSOVMWc9dbT4CZqGPk
GJw/euGJEbakUaMsgj6t5hfY1Xok6jZ8xQfBlI2fhE5/Bz45daoUHenmGGbuXoUtmcgS8oPNSgyV
F3HEYvQj4FVzXPQRY/DvJeBX7UWxAsYw/70vHKIzOfgxC5iiTyJOLV9ntLGH5Ga2QfZN2NOJgTrg
lMIEvRQH78wfK4XBJZqOgBI+Iq4bLF9DtzGioe0ZfiDGQesEnqY0GXKM4oS/C8hPcEigDi9AR+n/
BUty4tKs7MYoJC9EMRqG6lMQ5lZnDOowfMmuATmyC37cq/iRom+lRPtYCi7ylTcxylTTeWRy1mXF
m4SJDjsgD7hDgLEzeXjqkyxUejP6UU6HcmZgkC55qkhMegAkxqRyxaWr2ztAHtXIWhNc6ez8NVsI
xoRVAE0mL6yB52lWLiyLiIM+juONk9lIHyS6pP1a70A65/RYvhP6hKrZ/Ps1+B6PPdEdsBmGoVog
9zY6jU4EZ7uQ8Dl7Xw0lBMraPnskiHocJxwb5d4+tjgNgSt4Og080AuqGRSp3DvWeKYJBiHp33mD
4s7tHIciGGCQ0vYArQMfMbn/tFpGJZ9P8/Q/yeDF+QPhUovY9W78VlPum6rPtZtDluAi9XYFaj9z
/PtfoyvLRRHQ5UpEdE/isS7JFKsklblIJL/x2My3ZhfFn4gJSAS/pMu9LAjxpofhQSypEA+pa9/1
iUdp2vqAHeDF9rsDAcz8OS5uuL/fT8Xyrb9U+qC00JCRFN28xP53pSzcrNQBqy2ZL0ZdaCwFNc4f
9/9WCKwbzY6iWF9atE+J4D/L2yIORRNhjylm/iUFJIKacZXTvUP9IGboUC8BA8bIp3ED4eVBexJD
gicuDEn20GviSiFolK8U5d3mtp/OrZJZhTRO39t9PC09zVYlWvfzYsZP2jbub0a/MVaWtiq2QpIX
+vkonrkw7D5vYSwckHTHP2ZOo9IrsNSOI87BNqBVPV5X8LgjqgF4P1DOuGER1XA2hxE8xyqlAbaF
vP+ccnTUsUd1iKYas7giCzZDhOkalUehla0ilYp4J1LUG57qRubE4YGpzaMFa9hQquVRZ5oUJ404
+sdqVOavsJq2c6EJXRWspnu8X/rsqJYwHznK8NneJAliEuhrqCiH4zHcNH1aVCju14BJIr1IQu+G
mxkHO01HMBG0/Jpufg7oXhKvRtJOeKo+LRu7VVyDyOsDaiKkVPT8h3DrjHkG5k4IK1JMRCKXDz4P
y2HoJRK9PR1RGIY1KCduuLB1IMSwtRul3MEBy3NzVrpWw70e/91Fvrc6mj22IYGy6gQlAZyjQxMo
MPx51ooKKdLvp85+RY94ceV+tr/Xa6SW3qnt3Uodh8z27fo6VK1B47tydq8wr6gS7Kj6ybwmxbKN
LilMi4mctontbFrSNlVdQ96Y6vWsezMn0s755a8ltXaJf34DSo2WkAhi6DiRchqPALcDjIt92N81
yVGgS5BmdIpfqiclV3vUjcdmbGT/791L8B64jcBURHEYcww2f8IxqWP9/sQyu/HcuJ/y4XSUylXi
C+OmNHrULiBCxd/G5fCWgTuw8ujp1pOIkaW2t750ILyEERnQWJd8ALSHCllizaSweun2SjlB6159
Jtc+qK0oxwx6aLjiLszuafdqV0VPzBQbOycRIcdHoOwkR/NsHg2rL4/BcJC1urm+e+clDKaMVA7+
Pa7+TVq3DNvSq37Y6d9MuxHGopELuvS/9UysCo4g4yM53huKnPSKVwdV0ku/uX8yIZPLGzM+ufJi
hTS7p9ueLDhqSqyIWA6wVBWgXIzYR3bkmyFd0YDm69IP0Cyl8wSTOvtDsX1siMoNQaDyJTfTXIlG
+NSEOLSFqs939kdXIpxhrrQv7fKl32qjTDNtKaOSBCJNx4z1fDSUnV5VsIDmMfQ7Pj2P/wtoPX5i
JI9gLQWp28x0hscONkg/Fe9cWwCgmDLLssIJOpX19HX1VztqUcCBwH0A4GBo6irOt122mIlUYzsl
Sx9sndnuxzi4ssesJSdt0qdzivsFhxE4FcMmcMhDjS9MF3wdcXYsM8Ni/kgl+mqSYedUDO4M16LH
LV6NEW10JiEutIAUQ8wCBRS3N5zffLP6CyVWhJ9Hd9wGm4fnw1uP9D19hP9YpHuVRH5weSBpRi3L
FJkpotad+5JurNYtFM2Ghf3oGU8iIUThI00jrjOij0NnWWuePdwUhVH5ZirzdLWB9AvJvDq9w35V
XDumb54esKxiRRB07gfPoHWkQ8/JMHGhnVec7kx7/i71xE8fe52pgDGmou+T/hPOGbyB4xTXXAh1
Y1vBP54v+oOeqD5VPvtBnXnbmTRia0kLetXp7r0rSPL7GqrWK9SM4yCGoc1OVJoXOYMokdVQ3gyU
XotLohPjFmnvApbJBMqPKrEDoZPP2YYuX09gDyJsNlWIWXlOFN+KGS1MFH53VwBgIX2tjsHIG3F8
dMB51jkYDslMIYJkHLKecNnm72tkB7zaWJZ2NgPwhjNJPowv8TAmiVZKqP5BQbK+MDMGxFX/vwAq
jc3IFMuBEsVzh/KtSJ/qPkdv4ggFtp9dv9dxsjkMDjYX1P1npGUmbQlLy1il/biBY3iC+nEH4c/4
JHnnkxqcwT6ZTMSXZ+9L3+NrIGVi8scW9BQbpHB017Q3aGlA7pn/OpNBWjD0J4qe1ZDfMNE17yWc
UQb4vrtPlStQ4PWpZU6Cp6fXofxIBsjom0r+wXa+bD6MGmqonESVUKtfrm26RQp54Tqhaq4Wu2PY
U4w6DGwTR5hWjxrTgceMRCbV5aax9a4QzbsmGKuzPseqUo8jKAP2jX+KcTB3mqG1AFKHVet0d01F
kjlup+GbQ6lgIJ6wadJ8CFnXBH+nHkgkw9hW134ctpC4nap1tgxI1xJQcqmYFIqr88Nq8GLGFn7r
CABG18OFNFnAGgTiuE9Hk5bVETZ6h5OwXgPTwhrDczxxjpq2DkQpP/BYzkXi30QhKyN3kj9YDWP/
FfiYXUJkGCkcy4xvqgJrdLzhWWu645bOfN96wI3bqY0WyHRHVkBWdjbTo9niUGNN41N4hlccyv4m
waK87bWFXNRywChLVLXPHvD7G6w8RcaNzgb+NwZePuVsV9LB1SLupBMDHjLpd4nhVm2nepH1GNXH
6s+2750SDkDN9yNUIBG3RWKUXf3VW1UFORffhWNa2AUoYiG8N62mOayPlH69AtFnyBK+gQKHMQMa
gwnXvhdEQGBhGNtAP2XDukd0olDHl29ISlAkUDZIPfM58jVPByXdeapI56iFCixkE4zdokMxrXEZ
kg29CMXkTQv4ztafn0bJXkHvvOaik4/bXbJEmLUtesnPltNppZX1hJKCopAyarwpgKTYDNVekhsI
SAmxtAmxp/gkCc6NKHd7RGvHbnVFOXurG2Vh1oN+nPTBZLcq2OW4TNjVbxswOYppl3BKKYid3tCM
1s8svctQRSwIbpc/J8Y7vTbI5zICNWcH3UZE25Z2btyrTzDeS+dw3KhPUHqLW7JBX0K+nXef8J2L
0c+SCEP7qzs5waCLxkNcwzqo4hwhl5yrwv2pjplRrlAdPh2yJmSy+I8DGas6YgimiCbLoJyKD9zN
1Bf4eje0XgH5lqS297lGd9BPP5Sr/3OOX3cvBKG4UzXneSyzHkVvOrj1SQGuESvP7IcsbHdnkXv9
J/1H53cSes1Ci+6OBA331v/rQn0oMK+B/ZhXgxMnZwElNiAk/I783jBwbr0z5OxhMgfnBMnnwUmA
HQPyITaD2qoOZ2ouYiHPWNtKS9x5HmW4tfGuc2JOJMwydY4zUNuhoRCp4m0UvMMJNv8t4uQXp9cd
fY+nKf55ltU0jsWRSJ315qGuX36nQ+7PngoFpFpfnMqpCrkqS6l2h22vU08wVRD1IyLNq3I8WgyG
E5uJ4F6w/oRFhh1eFEUJRcRmYX8pXeFcgV3LRqGFHS8lfsKimwKtSFzm+DjA2NoCC7I/v8gxBN4q
qPAaK/ddhhApc3Nu9OZYUHsMutJlCddrGMDwtVxeWCGfAVSt/OB036MDqnot4nOEepTdFS+de7Fe
YdvYhgW1zwCQDFx64PTA41LWV1u/uSlhDbkezKa9HijPe4adYOJF153JBgOQRpq+VQCocnfDPNc3
x6B9Wnu+R7WJnUIbl4hts3LNed+Jf3x2joJz9q2mUL9OE+riiJfKSSlYPTyltFa2RXk7t/80dY00
feyt6bNSCwFy4IklfFydYiFx6Mi1CtOiscf06jP4zNuVzrDeIEdAZ4YJx6+r9qOZBEI654+TNXWP
Y/9OXIIO9XH9CUDx53Rz3eiF3VoTxAL6gFIz3gm2cC1fXG4S5okyqNqi8RrCYMMwpMWnT00UZvWH
DlZqordgrETn1WxvKzh+W0NmrtOreOjIVAuY62x7qalevEYOkttbyugS6NlcycEUDqSv0cOXnWQJ
uTDSNyoL7EAVgCR1rylF1eFE0FozfQQQkQ7LLvf0VO1nUG+icbygeA+c5EDvz950nW5ldy+lb3fz
jgPprSbF3YMCOzh9Fo/U8MJ8vSJcXcBl8o15InfwDcvfMIlndeb2HWV5KobUag25PaIKYeRidhXw
fKFTfB7U9C7aRaN/Mgux84r0nIQ/B6kB77W4l+esMWzf1reIbN+UdmZt6ES0tKqITDG44rqpulh4
1oWVak0oAKLrQAQ+UEs5K5NzhzbEOItwNgPAqEYAdJq1LakbWfMOfu2rGJx89U2P82f6xwf4CCzV
8C2s/0ioXU4fdFrUdgZdIl5sEXZpbDetT+66sXJhkKermH0azH+F8JcGiWHCFB9UYJ5u4Py/vv0U
HRN57Worj3e4dwlALQ7L43LeW/EkoxEbq6bTdaAXQGg3C4jeAjW8zEaS2Gtg0W6g09w48p3hhfRi
k1lEgamEBrTv6Z0FOaH4wCanedkRyWXaE0bani7vP1zzirGaIXzOySTwLohH0HeZgOEztbv/g5Cn
VygjcB9YEQN+Q4m2/556pNVjhhECN+aOpkMlsHeBvski29U4KuuLJpkskgfhC+FbbO6SoVM5XYuH
gbW6UtuHmdyXVhSqYyWe0fDWyNvAldYPiaOkH3uCjIc0p0OVkRmKNyOegGOHjB0uxcDKm/ehsIVq
c1lq4uqdnR1Wev98MHxPFZ2rM1u4H8oMrBULcUdi5q1dtQVc5ozy56iJdIYOT4vKlenKeZ9tgy9e
S5c6h8Dn0B6UrurbkH18UFQFDHxOrNsmCVfMnVBXKl7xy0bdxD5ffZdubPXyvhPkHwI1TAG90h2S
L0AIVz4UrB+4RCf+dpsqV5Riu4WCpIQwPhnICY5rdivsuNEcGef6QuvHdJBcpDQJbDfRmQz5UvFd
7upyMbmT5CTjfw0Wj0mn24S6FDt+sFdBtr9kETuzvS86ocXxCrjT70Am5F+H97Oj0KHxNQicvHZF
fDGazHF3X5OVy8rxEYzcWfQCY/Tso/mbaIPkp3PbeMUR/JN6P1OpylWf0Rm10dOXSkxUzeeRTbLG
0yZrX9TkT/N64EuTLhOsZTHo6L6KIyOoJBaxH/u0NJnNt3DMb6hv3YCrmrFAFQO1M2H24phYT6il
31RwAEY1bYa4DrpWiwGVhTQtSnUWl5m9oA1ZOUt/g6QgY+AnhAYPUh/9C61Q3snVI1t44xvxmo4h
QueZHeVaXOl6TuLxJxYq1GPRPLmXmgTWnvtH4IFSb1KV+JFByswWtkS5BXAC8jVfEXLsxPDFEhkx
bqBDx/3wiqZSyPHuFcQSnWWneFiKMbQvxxaqwQNKNw93FuXowuhMVWSK42sgtkjMGRRa30zBsxxv
1BDvy202jkvdyCkYBJXyas2jsaas5iALaoIS/38yZQb/dbKAKWdWcZuIQ6GquDGzcIiu6fNGPMLP
GL8XAghAApwq7s1ctY+8hYeQ+1PHNzk5oADSoXhzZJ6GCXZPpfmL0KGXyD8v5WzEyUtzKvvvoxnU
2bH5Dyz/Eq9hsmRssVZsP8dmsUFmIoAe7SVkUwHOOvBUJPaLy6kQZU8o/nfPJ2tda7SV2PJAmifl
ahz0ye+JPY7GFjd7C/m9gJa9hQ9DvJwikdvci2BkOY84T+tQU8cwDAunsIYRaYX3g5/0M6LpCPO1
L8zMJnqrEsVT2lr+2X6scA2isDjPfhpDZEn30FZr3LBavr/MfawQEEFHAhebTPKEEWrLmCAQ2ToT
j0/xUq3LNEUTI0+Kpr0bgM3A5QUDPxgXkEkSfE+9OYLmWawCzKW3f5WdfBl0LN+Tv8kpsL5qmUAM
XH7UZ3Y9cyd1hVVMuJnTU1QcMi6cEd9oB9uAQtkhkYuTVqkgfeoXZ4b/Oe6hjFspndqkOiikEGpN
CJ3ma+Ut/c4+4zqhbA51vY1al7JoievbsK0fOKjVrevvEzip7Xj2sQbV9a+b/WRqbqrRu+JwNwDM
/KrEyrJIBsiKXuaGs8blG0V7kPd5Zj1hKVWm4byKwHSRexqqxOQjsQRbLEkWjOkCxg3dxeAQ2qch
KYkrCCiuk5JSF+Mk27fCgXIo4sACQf5nU9Ja01UKkilKjMudgHEbQWcQQptnmEVQWEh7xMbl6y/P
mSE3Kn+7vQi89AzpIoufFvsYEk/KjGcyfZs9cF516Wsu8eTwcYjEkd9FloZlyKlyWew/i/LH1AIA
tP942DcA7TtTTeu8LzRkse+5BgPZOCwl3a4geDz1Ldtg4jUNL65FIcKWrnZiWJbzJMQ1mbeHL+fV
y5ylkGlJ/NYsEtBLZ7pb2PgrjerBDXDm3zGoT/QwcACUnli3qCbae6xav/uXRH/OHd8rHMYV19zp
KCxRe5XwUb1Knborww8qBtqKsQp7oAOWKA/jpxv8DP2M78eL9g4iCKXiqcxWV0+jXmPSjXL+u2hw
Poo9RSsuzoyi3SGWzDn9xZs+kpJ3iA7JghbBm1nHGdR3WXOqBioHar1UO1qAMaqVbibIR8JRzoe3
Vvc+I5xVOEJT+kQCubduQmqhxVehD0doDewk741jHJlr0y/HVFVgQTwF/x+7XXoL/iyvxRDkcXnc
neJrbpSUkeTJXCFjEcs7X651NpocAF8+IUyFD1vmJTIO1MauFRpcZcgzkxkWrWM3P64H34lfpps7
qD03D+g/wgKQMo52A6Syi7R5vSWLclmWy08v7b/fj2DJCJKQUWb7av5pIsrEMPexTYgpQiHLqA9W
y9KaJRyNj2PVMgC+/IDuX/L/0c8iot2wcona1FohS/TdovsDgLl/OnKhGh7ttvg00m7QKiVMFAgZ
oUs+QGqivBixrqdZCL4n45PbpAyQ8qs56ht6CkmgSTlOzyYWW0w39UqJMFt0UF9mdl+qXslSKSdq
Mo/fi5W6odjxted/rOFB655AyHJoKHmMU+T9Wij26I7Yxcdiyj8oiK/4LJCvFO2hCEqOfrVNRbnS
5f2nf5fzx5B9P7gpFxEhR/jlYY6tyBekChV7CDrdeJ/VvsQamIucy71nhyxE0LyYdthLPC92S2ri
1npRELiyLw6mY+/XSWCxqIY5zwZiKFNUevLnDqymQd6WG45ese0lYGAi/6c4Bri+L76vkR7ASdq/
rC1ZzBgZ0nlbQy3obOznj6QvapLgsoNOrCeap3zAG2S/WBYHZG9mJFgjlkwD7dVR/WuHSEi+KWKK
jwjG7kUru6EqmKp4pjuEj8haao85PmnXK8NCEINu7Fx0DcaC0qomPL12w6kvf2ws4gEuWmfa4rbH
+nWJMpdknKNa27adFOz0W5F9W0ahiom417Xk9OAaaO+E0zLHJ0ZGCzIPDAAz5JtgXxyzkkWEXbN8
CTJnGDH3AeixpR/rJlHF/QGF1ypM4KaRMN26kTjL1GjdC55dk90RMuh0iiOJZUiwBB4LFo19w8hs
PIQIDtJH91LqBLV4aIMr3ZCnWVr8k59xRC9/VwOnyA043JTXAEUvHDviNvqNUXaauJvPuIbgLgRj
lwQarT9LUxcg+GIFUv/9+ehNE9ny56WuwLfoEiXYaZGl8vkKh2uvlxcQlObTj6DG4P/mwktmet9I
uLDGwLitCgGfgo6I+iQ+yGD9C5ejn2N4i8diId8VZlnmpvjmzP/lO36w8DKTkIS1ot/IVteeP1R5
rFuKK6HHa7v4BPyZx6s17+GL81fmfE+oSVsNwrRDM3bFDnAqa46jQNTaPI9rwi9ehk3C5vCS/Vi2
PUB5lMPz+tzFcGo7S3v3Net5njmE1rkDVaz4EKh4OlqE+IAmk4SdaXy+S5oU03QunZcJpPcIvXKC
BxwkmGsENg7rFp41xpzOn9oM3Z19XVSL6k8M+KTBy0dU03uOXNDu0awD1XwNVuqgUjlNDYSfi4OA
dnAa66RoGCk3tbZXMCV1gaNypkcQ/EL7Vr5y1nvWe59KH6mQFcDbLoDvVwCEOazvCU4j4ogr8nx7
thLU4YlAlX+liDmVTqNTad64qDPb7ltOFH/MS/Sn3TGGvDaONoKd/iN3q0rXRIv10s3a4eWdj+J+
adorjbyFeMS8evlpeZVS5Boeh1KQfxtNjWdFqPkosqZWbG2tsQx5Afz0jKqlLa6odgoKxOsVFhBB
mBzNckv1h1ghH49YKeN/6vjXXiGlqqOJhX7Qagq30zYpDgL3uBQgbWO5jNdwBxAWPrR4wZdUZTcC
Ck67NcSqitidNcRsfLluRTA187lT91C5ss3+JREn70p+G5Z5Tu10cnVVjnrLieRTVQhJbQonJb3e
hxWDBzmr/atK72dqWnz5OANifHz7QBh/ooJQlc/eqA+6S/OSYXD5WmWM1sqQc1VQEWQ3rv7U8bKa
kT0oZZ8S7uD1cajI2bEMqr9doyxmUUWyAVACotmQvi9EPrOd3KbCiL15Mf45A5gPWCM4IVlYjtYi
iucpAyePjMlIFs2Gcjzson1stAGeJKXWVW2vk7m7dqDCLM7oLc4o63pwxXpwLODKDe5sX4tq6gGN
vjYQcqiyePszRmxBbq0qdOx8xWT4uNVtNijyU/yHSPLvqC/j3JTcSIikeW5oDRt6T/iwVXU4B69f
/X/wibbEjBVip+GyW3zs1VyMa4aEj/Q0r5J4HMxYPaYvOqTSzGUmpUkB5+1AW10cTcAHEqyG28Zo
LC2Wl6C34JoAhSMAV5NG2nXqh6GySOQT4LlVCrwdGQJscwK6iWEFqFzw1nzwtLC+1u7AXbcqvGHc
7/vTBLowPSpK24v9i8X4bcx+GGlRoiExi6ZrV/bm3w4hmH1D+SQyMtqj1HaiiUP0N+D/9ttti9fL
IOzLiOZevbtYk/+DwyBKAhwcBEbDH8JPCMC+2CQcpOkeAw+SNgTrWvEkBa2Bn8Gnw1fiu4PqgZyV
CNTnC4Oq4zTVPFXEVkhDTKEFWeIgMVvCnGs4WsUur2/uG8OLfTn8/MROVdnjnoks/5KkNsbOVrF6
uPj7twFhnoPh5B768YBlRdF2toqOYDbIh95gu/JizHMbUvMABrIoal5kC9SDqhK0YFji6MjtEOIj
6SjKQY+9k6EfbV9yuD8rt0aZsTzdkJ1SGsPH44O/5h7UXcqa28n/aLxoBfvHzArXmciA5v1VAxmV
VJ7sUGVCB2n+DK28Tlqi7We5n9RtMXnsbDOTyZw4Ch2beUhPrvKfNuwxD3T+rIlFF/FcHpd97p4k
lhk+h2B3P2mzgAe82j2CtwLXhx1Wuqtl5z6ugF51QRbt0sSVIekJYyt3ECSvN1e8RR/S0f5cz3SQ
qZPJ3q9l2V2Ts6ptHWcvXTjm07udfPhmG9SUeKAcxeUC7J/ZDysQBh4VKxvY/eHEo18KIlMxjJdk
sX1SAzsYC6u0YsG6OqmOq40Q1K3WaEO/RirjacIrpLZWiKqxLUH1T1ECw8yS7KATpHBkzzrDYPRG
+Dvb+tUd/cjWZmhG2/ZzFDlJOj6eFDuSYDIUM+0ew9hoKwG7MGzp/zYesMqUHw6ostX/5Qp/oPbv
MTZoYDx4TJdtFANVdkGSRm0476mv/29lnJiBbgGiykuMUDFcsvGUVwcxbPeE6dpSoJe/2DGDYuhD
mOmGZNqhIZWd4I1WYxxDA4cl4LZII3upMHzxQxE/oy8QqEwp9MMyc93EPb/yB2SMQeKf4ByMN8uI
HNOjyCbasiw6uKVfIf359dl7zucFmkjJUGdTq7OCNHZxZKqi5y11tEHROjlBARy4ebss9xf2XEEl
7HdC5bkV7JFk/eQEmfzWFR4gYDJuu3q2g3Oco2ic3IyAu6pQGCJ+06GxbEBguWw4tySROA5vyIs0
tCwyFlehyWkhAAxyW0SI5flrYvYAotG/3EOYwqRE8Gb1SMWeRjP8aqGhdKm0+zjCw1Xh4/jQ19np
VSJPOpNu42Y/0ggy+KAl5/kWT+K60UUAXwPwo0r/RVIl/ApAnx932RCoTdxRvvnr+ZLrV8kaTm+4
vI9KJJ1jfnnM2iJkkH1nxykj8swPBnaTPDQr/yWmONs2q8kDr7tglPEhPgt37F9I4QGZubNR7H/+
u8v0r7wZmMHx5Fmu96eziblCoL3ZkhRt2Hq9UXZSeKi4xIKMKcbFLFgDO91Sa6Z283bJACOZ87YW
AQk0B2dwmTMgIq9eF2A5+Q4Y3FLDvTsIWemCYNDSbs6yDWCJGy2XHdHRDGmpTUWsvvthHmE6IrIn
xdMtluw7tCIl+aYwYjJJrdDJTZNaxfeiBfqANDgbj/RoCrieoXtrXM5RjCVbb3KbFYWvPMH7x2jR
/T5n5LDF3WIEwkd/2u8bZWd8c5lVimmbv0OPdfUnybzER0aYgJeDRwdjIA3L+autvF9i5KJpDeiA
nLY7XmoS/B0LLSuQJVqjfRIxeTnL0kf3yLOWZNQecgkT9aHj4xTltj875Wx6eaJ5rmgVNtdv3fmi
bkm7KnrpT3udk6vHi25guLlwSIiEOKXaBVzifsxy4ooqxaQTq16B18HoygkYeGwtXT+ymAWuWiRj
Lg3tjlHpkZH9fPAKZ/hNzcERm+asEN2W+HekBgBAKs7QP+UPjNUcL6ABOWVYUJB5XS79a1Pdb7lb
vhuw21ryvSEl2gdi8/4s5fD7ymDwGI/mtA/AmYRRB0tE+Qve3B35seNcQorhEhPAI1FKFIduCrQH
/wQcrZ/c6VNDag4+p7zwpiaHwIvyeZCdjWsjgdC5SjQgKdXsnZJXYH/2L8aVdlApMnZiQiG2qKfC
E8J8okN96YAgn5C1e/EL6zIm77s/jDj34WR4XfzryfosZI+SUR+nqTHXOsSbuo+DkjVByYphEQEZ
uPppl8gtx+Z5u3UuNcQeEeDMmvi0gPD76H69mcAPTULt4l1vQqdubrmHDwtGvMJ162QDbQep7xIP
+nUadSunxxX6GOmcvTLTQWnlkbAYUk3Nw+uMCuPRXjWRddGJkDb7DqH9eZLcMboyppj8j7NCCFCY
DpaFPk4PRVcbAPB22kfZzIVhThvqpvA0Q6kIuwoLI1+BfnZaP08LGCWodz2Md8AxNIbpQdY9gnAa
/N3E2ILEZLJIyKtGjl67mdm+oGWgBIxaTfNz9K0GQ4zP6yWw4gA1GePNonKkK+R9ccV/9EsNJmCA
Nl9o9xc1y+vYNPEQ17EPlhWELZXYEeZAt/qjv3T7AvwrF5KljQCEGjdEsJsUO2MVHXAvf6HRDBW9
9mCOxAfSRcY4r0m5EEMFMaCk+MH4NAVRLSupMd8i0SxjnBqtyTprNU7kPmKXftI8XkHdC7Lc7VyG
bv6WPDEc7wlJGq3ChacQXh3o9/mfmTDFceoNFtGfEvqX1RWu9PMW2KmdiYnJP7q1RCn6Uu3Dp11V
FTmPpVsHPf9boCnRBWPD2NzUuGIP1SLM56lOuRiYga5hg4WKEvaGvQ9waZxblcTcM15Q1X5kSEAv
JL2s69dyj5TBRdr3AY4PMombKcXHMBjZ8PeV9+JW7Lg+9IqtvzHYWqYvu0//kJQE9ObMNUT+IczR
eRB7PJXob3Ta0VIreadPJ8o9z0xmGDPxUCeClDtOwS9bbAajrHpDQ6emZoNqDIkVqhnXWlSb6M78
/ta9sjTow5PVoQ2wj9Kr6Lu5pQDKP7Hu4wKNMs3E0R3TWdbM1sikb1Dmd695qSMQIVK5ffgJ+ycU
ALUyYFmhGNWC0CgzpjSzMTPALQPn+xvQSgD4pHVzExg/uaor3LjToCK4TOMDYQH51qJIcqzzBeV3
qfdxt4s9fvDNRw5HC2aWeXaN5xjdQ31Vqgq1pRwQyxna6ZvYJRh63nscXursiGpYsy6cSwnt6pCh
VmX0/WK03+w4wwagdje1v+LfxsJSXQigvUJufbwhBX1bO8qjN2F44VxIItiLiLyQdBaosb3BAYn7
nexFU7xfJnvsJGZWiB7ksJSoDTtRlySWbrjbaTUJFixz9C06j8fmecQ1/bGLDP8vQEvyi22gYTaY
7PgDt9jUSjhKqkeNY0BXwMWDn64xB96v7KZtFWYvsbX7IyhgGREDV5txsmLRikSBhpu4OiJzg29b
quD0J3PHTp6x4k7VjvAPc8i9ACJjorncLAcn69HAiGMJA1xgfGma7Kv6xIh81PxMPZPZPdmoAadB
edioOLYqiRBSMJH08gmtQRcSA7DcfYBLEQ3zs5glQ+W8Wfu4vFcQKANBXSJX4xcYck/GV5ZBhJFw
T8EIliJT8p3MDhtejVzKRU0HO1R25QEzq1hUChGL3rkAQKdXLUjk9Fji6BqlahHcyebgUir0oX4n
2vEHUEbGWo8k99S6GA6IXdokX81Bey0gk2k9d0SosSwHLjYnFLn/wp/s2CZWCw889+aaA+LwyCNA
3dUY5EvbeMg/hZNGrO5aif7eM19rkVzL+YZXyRtv9zKPELjRL/IiC4+9Ffhu0rWIiMPPiE2NbLM9
r2QOhaGrdkffNf69EVWGjmYxknbN/DgXSsEKqdWUMt2bSBdd2lvwZy7fPIVaFhrPKb7wfBs1deJe
7UXfGin+BWAey7Gt02yJVeis2jvn1Dv6kzxWRjfIlsn8tiH2nJJio04hBophl29sg9MSUl1iWT63
9132Optasuj1l1xiBAB3yTCbYdTT7ZmprjwC3KHY8pgzu9QZ3k3LiWsyk0MU4x+M0dmJ1XkUs+3B
yYfwBqN90KzrGD0cauk4FwTXDvvdVaIKsy8hJIwVTd4UgdbRQ/fQDJKVmfjZghWs/yGxOk92zAVd
96yjxMORyDKip3dbIDF8dfF3VmflzjDP7NSTN3mIjjmP8skP+ikfIGr5wdATytsNvp4gS9S/TJWV
xZHE5iSQRrxg2mv8zqN65dtLGHez0i6MYdxXXyKcAGAtCUeCenc+XmTmD5d7IxrUOPaY7JphovL5
jQMfzN/xYLte4NqMUxR8OrGh+bWmhjYc8N+UaXgtTt5gtW5hX+WOzt6G/1zZR0RxoYEORolVZqbK
VAo48CdLjybl0csyQHkcfxaP6tB9mLebFxtprvxvQf6DIB4dx0/iW+cl5cgfdHmqPw+/iucOUKXd
SuRcDA6AzQAU/5Ha2wRfQ4tcVtVHeokYrWHQsa4LMNNFAvHxTaqxxxCuLD/MiBNYyKnMAPIYoiwq
eM0HhT4Nr0cY+yh14tpPDrDloR/4e6Bs0C2lLqFpTwoUZyJJkSbXM1afxtY8lY4yKhiU1rDE3gCV
hHpmc/sAiIaoZSVHLyYGoK8uQXzyqew1veWCvfNxV95UWpB1x6dii0KoED2gp1lX7t4+PS/3E0Tc
ucizdbqTVlJu58fFNrc+GlmOLRQRkL18yzOoRFh8PNZEm2Pe83vnAXHz4PbibKealThhC2hzw9gK
ZoMcefT2H0Ky2eKXJ7vsdJQNpdoelyZ891ConuLz7S1pnhGVn2MZ7p878T2AY8nZOTK+QYQV6fnC
osaqd9W4T+KdVGKGUhYopVFGtVlz2KJezbmd15prMeQtzT9NdfXga2uSMVyrgsB4KRKMWQkT6Y6u
bZnZ+mr/LvhqT12BkZ2slKgj93W/5yr/srhyFBNS3prT46L+tDNm+yPDVR9YHBy3GlYdjBtiatT1
9HGUdjUGaYhJZMRS9tXNDhM6bgEmHtwIXccvm7QG1Czk5NboEggwgaKzb50n9fFu5YDp61TZdo/G
4y8fyl/WfsWKqEG8PmR4hAETQgTemUxosikhCePS9up+o8ec0dX/8jWfwXR/E3TNQkPpz2TKPt/N
NngfsR2/HEMUiZJ6L5VZkg152eQMv0CAfahVUdE3G1Rf2RpfpOdyu/xOkX5jOf2woxvDiEAfGAuQ
2h5F/a724pgR2t6PtIVNg4r3G0srm60Ie41Bd9266sT2YbApTAH3bYi1gOWSO9NHEEdYvhvLbmnD
bn/g6if+j0RxJlcSbuMAY5QXAi4AfdF0AkWnK1mR5X1I347kxq8mZKsN+BXDw0dyLXI3NYxJOl7V
8tGsW8wvowZxM1lZXJbhI2kCpWk22tCqMX3XDj9DYc0RTWOeQq0syQg7t2D/7LerBiT2/n5CaVFc
RixDdTL4ac464Als7FhN09hf2ssmuVqBFqetEdeBQ/nwpng+ikHoGdyZUfFMK9nwYl77gyh60Dfm
UHHU8IGtQ7b33eSxtcF1AeSEkW732JCel4LAMBYAfgAOGzxErb3rlPco1sx5Bb6h0bk3o2WRliZh
svRiSKjSCi20K4GqKEgyn3GLnG9bb6Ri/vaBQ5yLqBE2baMGWwNmReSQAl/CM/2IYDq92ijdI/ec
1BYoLXzzVdQFnyRR6qSiFDhO7+7JmjBSLYyaZkgquWT0MF4gLX4D7kLAw38BAQoErrRhZsLPnc4g
A1M0XiIX6qKDzhltflW2yrbcZHGjr/U+meqRGvGEYPhHSdxo8qkYs8yxZPEcSm9Dne2fnotRuHPE
Xb4XjpwilVHS0ytfz+J+fVgaVzWGxVAOFd+4H6v+fF6YPS/hprIB3yT463XqjJ1RIkGnZsuNymU2
DA3HA+7f4hagZ/ncpE2jxhdI+oJBxEa18VlPQkStua4etlSINqCIq0DEEZhP5xurHnwNf5uZCJuf
uijyCg52Tt0gQRmX/J6SxvBPq1N0kD9h0g3Is7Cpq93Jm5Cmb400kk44SnNawVYFoZ+WBDsD+D+l
iUX4b8uZkQOGeLI2k0udOtLnXuITE8PSIse1DmXZJi2au3MyoOK4o1sbXb/+aMmoY4HV8QbjOOCJ
1+oCO85/H4Ur0jmTa/ZndteL+aL6IDa6OH1PwlPe4xt7r2pwI/UtWZhSu4EXYmw35WxA32wA1AEh
KYHNy+4/qhPCqrgOW/dazmzRnXolwziogxgCaI+VunYl1KCntqrjoSzq3mKWOpjNuYKVjg4tvhqv
sr8Eq7k8/Q3/U4TsYKTK5wMMml+092Hdp8toJ8OF4SKp0rX7hcVVUtMgptVIOn16eW+3M0A69nKk
f0sRxEGQdlUxE1VafrZQ/isKvgGxEWp/q0+0JFMf312LxC5UZwKDis58w0RD6XEloQbMZ84TRe27
04NEMpm13bkhOmhpw5V10uhSGIKCo0CbjrF5NgP6zZsv0ORtTYvdmWOuqZSQafXhDc6Fwik0ZKlG
5lXCkmDFltEth66JN+tSNy4lMMDEDWGfKGOskqQIB9ZDz6xStoxrjd2SqWznhwkLJK0IZP8vZ+3h
KL2Xi8qs3LfuANDuOyKvC4fW3S1qF3jFcSgjORDB571trvmo9qZRau5uK58nZRDfj4mH6/EOwYtn
4DRVE7GGXSFV9fSJ1Wzgr5eMdC0L2zroIyGvHnumeL+Ky9s4fuscjBmjRETxjNnIH0oJeGV2e1Hy
5dYLPZ2mw/3PV5qGkFqhaKuzSeJpjAFK6Ms8BfAuJzxQNyP90zdvCDZvNDEHz1W89logxZ6OYhDw
dIwDrfBJeebHroZFyzhSo9Ft9xBoBGdYCmxiJEDsSjY5E76/tj4L+zpCuLkKCxVI2792+LsCnmbt
lPWrOrbuJPjnG4WFPnN5rs6THR6Aqz4UORBH/tbO1prhL7pfx1LPKWOsGzKIiA5Qotlx4SvPID1M
gojVpFMP9ct06mlcPQQ4XD1fnd7zw9G8c/vctiwpR8+tcu/BRoZi5VJkee6yzTqwTG2NiHo+MzRE
NByKFR0oaJQLfa1M9Y+Y9SzdgDqeBeTKr5VpuTmPk3dOwQVGwrsE7NYbDmXpfbixAOcEUcZ6HcTN
aA1bCl51OQorLdMZ1UYA4xC0mToVv1a98g4ZIWKSXve7siLU+8vBSWMTfttzlBZ3UaE3Cce+OmFa
b7NOvgZh2n2D8H5yw9KFxrc3N58fyhrkVhhq+DnzmXOblRI+T4N44V3yOdiPiUuuz4CoBm4dwbPK
K0CZZCBilVkQLPq3WosytCGuF31dGcvJZwhYRQx+u4Ze7O1iC/OR24vLvzdNRuO2iis6OTelIT/V
Q54kgja3/rO2qF8tXN+8bcoUzw/Qi2HP5/tQ5hj3YBW9/k/KGw93uHmWNSbRN/bUrc7cc+yTyBJl
bu+63IFHT16y34Ndv2NUEmnB4jIOlwMATCLrNb4zbVIQCWU5SR1jvDZYvQ1Fsr2NYDRWA5mA+ENl
iu9j3tHsgGLfr4YJdOiyH80lPJc0TidghM84lCh3h+2M5EDc4erv79pO5/8KL/K4XBNtXClw87uF
IYjajsSpEL5kg6jaeWyId3Hw4sfJKwPbdCfAC5dI3dvrEa0WEFxAnJMDWfyXUqTtIC8jKmRwC9Uq
qD6PLfP3RcmR8s1QOZQbIhz06auIyQPno0kBCW+wohoOFEBJUyFqp1fGb3qcZ7r+jJttbaLg34Sx
ND1XYjaUUbkSSgmURNmfHp/Trl+yk8pN/CY1XtvdOcBr8SOoslffIC6RfYJ3ZHhU/r+3Zx17uiG4
mu/K3PM/m8Ym4c+IH6QzBijMGSoQ9bHRMhvG5oGVMRHV7eyxE+0xPCCY/hKrv9dXmvtAcvJJ7nSZ
C9vMWAI4k4yn3NNexLetf3wIHrI3mk0mz9P/3Wcayev9GFQ/vA3PYgiCZ2NDA8cfZg+3RAmWxmwd
vD/Iq3aE7a6xjV5NGgC11TrNlNP0flZOwagRh7+L/jcNZbY2HQ2eWtQDVYf2bIJDmmbQCSfufbDs
QsG1YbiWYiKuw0sgxgzsuaFcfK5mV/mctwucdkJ424nJ3vbKGHWHCYNUjwNhN2rqLrBofS37BqKl
bpyKsWeigZ8YYymf9Tyj42N7CZqfnc2NLEdSrjk2lJ5PqjnIR9VwY+SXCwG8seQj2dN3QIeL7eWG
6scsDZv0+FdfpGruoY9hdcdEFJMYkHSWXv8AZpEBLaJJF2BE8jjbPZWFL4xDS6kMFpRSTrFd0S03
rCOgc0Vx4bMIOor8ETSLpCsUIPEKZAmomphaNuI4B5elKcEyNTy3AYG1PF6pLQYKoWeUAzGEpCZX
/6goenqN5KvyF8Papx5PLSEsekKr+PLzpwUJW1+IIcCCmRPE1KJ47wyLsoE7iG8ovxr0oQI+bDwE
AOd1BvDQ+orP4bNv0iBHFtgb/vP7J1o7rJa7w1Vy/8r0S2v4Sl1R/7r3tXAatgC4NDTxlGM8SyrF
3ACsMp0azztAQ9KUhxsZJXy+eD+HK5CHQZrQwu5COEAKgM42yhFj/xR8MbgEIBSB5VTwwm9HNW0X
ppot8dOHtJtxmsh/yjSB4gbjF6YPxX4fK6/9I3VhXD3QyfoIX1MWmjQ4Ie3sSAodLT5ZFARDMX/z
GYkLFj4EY91cfqudHtqxu3VMk1E01DTx5S2uQBh9X2jSAU1sqidutPfVMA1lXU3OPLxuVX8f/Su+
jVbQVcFL7TysWHI1FmHHDTVHovHBQhWoGK1lb+0HTvDhyFsUVFPT9/ywNbXyrGObt/5M1mfIadgu
7R0hNx5WKw0k1a9iVUhnXVIzy+B9HdTF4+QQWdY8MbJMoNhNYuFWkWcGlw/GE4FIvpeksG8mPHP3
tzFxGtVYedvMi+aJGVWcB8N7eFhN9bB+AXKd9/qNfLD4WrsxFw4b+iHYqpSKkrZe0IODk47sUqLz
0QFMi+zXJXNgXDMlDvEbIbtBJCy4J8dLfI0sjH3CmjzrTaPHpuXo5C00pGxzOdEY7gf1LgyHSXLB
rQN8fU/AtV7bKhcAVj9ICDZnOoi7pcyLFQxfjU8FQ6wxbt1MHS05kfiVR6X33o+B/TAHewOsiDeH
DrHcz5tkMYmRkeA900pb+akKOA32w8wmHqleN/VyzThpf7b5J+2MwAPvzAhWS0vyDEioa5lEToKj
30AWIjXzHi+TvzL13IYDtxppaUk2l1k2VbO5CxScME6Fsyo6gzMNBrQM5AKdkYk3f4w0Mtig3h2/
NkxRl/lb9uq/Vlyiyb/JQ6boMDqOiTeo/z9OAkcfZrT8gbSKZCFZS0Nv4R6O6wI8+veUlfhuy5Ms
HTpIyhmrHocTRr2SVOdfhm8HEXritMxg9yIkicIqZAVK05RfWKxtk/JnqoYsPV+IyWMq7zrBTZ6l
x8qaxbWvUseo6TDFGVRLkq6xPtm/pWS0Krco2s5q7hsDENheiXDpa2V8dUgnfb8KSk11rDuGAnlU
l8UDbsWOqINf9wGxHYGR8nYAtHYyRave3+pod8PsO90j7IYn8555TbhHOaKNiYub4rQguw1jjI48
5LvTvG7hIAXnOxbwGprJY/3RLYQ+i+WIecp4wfHABUutiDe+G2xKbby7lo8WWyK9896NPMLbgIsK
NTdaYkRMEufiQ2w7LHSa2ANMTJeBTLJ1bz+k+8lekI1byJbSk5LdmXqukFgKjSAV9FZL9omGKdFw
3DMMPmoazZcwpvQz/yiiMZ/Mvj0IUwWMjp7SndsNTyeuY2HRgpOhd0V1BOpNC5KoRJCbFp0duzl+
040sCY/u3ybMEwt5NbBOMiyiS1dQPTU6ky2mHGT+IxdJdy+2RB0xUgqN31evWJgtbnda3RZu5bwl
qZoWwced9oh7vy0IdOpfS+mWVwwf/jxxla8livEQptOPgLyrPm8+60m/iAt/b1yOTTn5xclXcNqX
DwmYF6l7v+2cpmql9QLICVeTjh8iE67OODgaXYAM/nQYIUxoSINT8wNa/W0NtW6AUp1AZ8EqsO1G
a3vPLDg/L+QmrqtrfV/7zmFHIHCXugD0BDg5sUN6hWeLkj+AQe/97Wud4kaFJM00qyiKDIaQ4JIs
hH+e1r7VPHUO4zZG9Tqsffw7aJyfUKin+HrNjrtYaEo3FPk3CfS6bBppW9fWrPaO3YeNmkp68Rxt
wPJfkNIr2tvquEOy2V/8mHAJQ3boTV9qgaVlBoN3t5WFEbskjhHDx9YzPFT5qOYvv5MpUrYf2vBm
scX0FVH0FWQViaonUmcmCJdOIFl8y12AOWbrJS4i4t7r7wEOWxYthus84PViBQCqDY+qghBva/Wo
jzhPkg+MlQxcVydjla5Rkz3nCnsIRbgOSTJ0xetD/68OKTk3h3crBF/29TTn/KvvEsn5cGFHCoMv
dububraiz/XozOMiFo1AEGpL6BwwqaSknAZrfj7P1QwnwnI6pBitKYdbyjD0iy5i7TVdTfesMfFA
4zN3Hlxvm2WoMXTYHtxOYAIdGt1WuB3l0EZrlU8yw5lzK1hmuOcxuER9SaTV04Kf9jBzE2hiFD4p
NkhJW4qsGVnX6NebjVG9neCESjUTAc6mZQZMUnZV8utGOPdATNv88+2lIHLSD9F3gGwjHk9PL3vQ
pa+xMoUni0f3KJcu589en0x+f178/DbvEdsfsU3sbExe+1N/zZhZLhaQOre8snDUNNNwx2AZiwv9
pnbHwZc+Ncbyuu9E23eXdGlk/S2wcwLUkte8GiIIPmHhDB6ukStmz8s1SF5N4zOe+8IMoYKKrpd7
2NyJUPWtVI8lkyOZwcvQJSMedoFa9WzFkNMmQ2K7+ch8EXDrazlJg5Fvewv9/9IUTISBInuGPAts
arQ5FYbO82hE6vyTgrQiSqSLua4gi8P0Zy847SCudQ+yKEVTSCSfgCSEfhy1FKT0uD0aceJ3woLh
s4Hbg+TXKq2428oA9BJ61KqZlv0cJD6Quj2jX3LHkV67smobPgxa50achnxGp3poOMvW69ZdMdC8
7zAkQDkXTEGbRvFEI4eO+fQV6NnqFBMNZbbdJjVcfCDS77aMNmjaInwKP+rt6xtsS9w6s1nhjPpq
iYvfpQ1/I5QAVzYO1hp5eilmJMKzbFG3Ft9Ck7+5UqYQicafY184MdAselwda8LzOfX6TCNgFgCZ
jAQD1l6jsWlR4KsVXI+lGpO2W1hWl6Y7a7uDwYEUtrNWUzSXuRF7Voh45EtzJy/sdK0ol6SNtXbN
SPWpAqzUXU0Bd+T7MYNlGrUgrZoTdZJoY/zkz8lTb1I0+I1J6krEmbAqv7n7i3P+S35a0AAMNi19
zs2ShXhRW3sai1Q3QZrAIX8UbrGE2Ske3PbwvC4jZ2mToI4NPpxYpeQrBcUegEtENj9fxTZUpLyR
yH/0wY3dAA3e+WB/UwLPPXUjCMGcFeU2W1xs3YesRfFMSP+eDwag3LtQnOz5bZJuHyKaLCtB7ECN
dPGs3Fu8wJzww/YSQFYCUKNv6Q5Nz6st4Q7VQgA95MKax8u0Xur8Q9cPqEQXjBmIX1ZkdcywNxkq
twywxl2YWAHOkXvXNyfk8b6RiEfuhwQxbFFLZ15uG5rCJNpn54cLRBEY9GsyaXVkGj2CT9OUUexX
LHR1hYGk3ORhyIShJBoMwpRAHnpBYznL1NN7XItHq2SBq5Idd5fFaj/Awhvvc/lAt6yTxDf35AhR
edJXbX/fCEfENzeLU/ErGHD5XtsyQUzg+XlRZZcKt1P0F1zWS5ee47opqhVCNA/2CyXtX05iNR25
Ya3F9N/E326RFQ76ZtFKDzEg3o9XZrGn/HQtrCNcJ/GT+WZE7Xo4G9oFytLZhK8S9h+hADl2+DHb
0ZBlhL58xFAkys8mqo1gJf8cIu/fgyrmvak2OrVGp/Sez7RQFV9n+GPlTiUsb2qgaxvhVaII8lNO
2SkmOJG6QsRyEBJxkvP8sLulZ+6UoNhn0JbpvzR54ydmkDf9Q4je8Vg67/QmOXCYUdUIqNrKrw1R
fNIDY1DWGNEC5EZSC+UW5VcMoEZMgDdNg6kgMcOFzcaGM1XUuY/c9bt7RgtZMKsnCMJXAEbACDW5
yVFguyJpmkIzqPtdmCCqZjm9GnBelzFAELGnItdJviL5gbJIHtuZKj+xUl4u2oOiwDPsRWIzZcrk
gUSLnj5gv6/oM6JKP8CaQ/io4dNzC1YcnboHjmspgYXlLoOjNNozeJbS0Tb7iz4EhxRO2aqUJE6i
UuQyUL5Nl9DXKUgaW8gRdWSh6oJ4m8bQO78BnzRnc7JauhWAmztg8Y40aORJ7QjkgXHEypHd3aDU
SW3O3JVGifFwKeWR27UPKDOH5EXZZduuq7S1mr18Xx0sZjcUZzf8n/w1KwaXuUHg3KVp2uEz29Yy
tmgUiGTvThQv87yws8YZpuOKTCBIx+I1/1FDL3f6fPXeTyEkzZSpArPYPpSFRVjV7wsnWFzw4u2/
Qu57qiNyWNmep8CskcCJpKRZy3379V+Rgc4jmhUqhlKrGrBJd4EPUIaT6Y+4h+fvZjYMoN8uU0i0
PujLIpqo3sLtu1PUBwkBEqNSAzNV5qt2FkjwuFg55c+bWS/H+mfx6kMFG95nFNwLMhFT/Pnc4EV6
31/bOyRQA/TnuEnHPL79+r4fHRGQeeOarYI7/qtGOVyjFG/+oDwerJxDSUDmVnchM/EHGQtZx6ub
C7qyTdurvKFrLJLFXJxEbe6U8Tc41D9zncT0PYvYatd/tzMFkInDrKsNJMi7RQn9XDgFOFWArCDb
WdgO+Ms52i6Y1/DylcYOuM53HlIWkISjIFfsAGwp33WSa8/rjuhc3pih9DzZgUvMFMEB5DA8tS80
ID8pnKaBGm37mOyoBbpPgDQ+GrdQ46RdxbNl78DnHvibMNR0cxMRqypoSEdpZ4P4ocPjzclvwJXE
JEqZfkwd88gt40YKWczBtqCON+oT2ucHUp/ELVrzVMkdlIn1cpvz4mL0/ywyeb5xwWPU4/tJ0H3a
JQWJG4j/oywTh/PbWgzH+c6h32D/mW+oWIL7Y9flBbG1DGfEyc2Ljb2dvodAHPFc1iXYFoefgUC1
7SE1cj/K8uXzecLmaMWdTH2c41IsOrflp/GJeZpNbeXGIfOyLpFFs5g3oBftpL+M28Oo7Km8bMB/
rH1T55Oz2uD7xugQGblu3fDBvqdDxi7W6zYSH7Q5sas4YE/ZkYZPqxrEtjCEfPZdPt0IvZzZ9ESr
4vRdFR5f/BdPEzJwUwURXyWTPPXWs1x0TKSGau0+uCRU6YDjLRIbd7NxeM1DZ5CzUnKUiZa7ARxG
0xQOJqjgcyMrLIOEKuRe42fqK+YWMMn9T57+H5zKRauZefBUd+5+iw0q6nSZMbvj+gGZA/tiybcx
PYuo8rif/ccExw29ffxMr3lebWOxgk6E5r7gtesiF6C17cpRTViWMPNRSwkLz/HhsWwPpkLP6Zvl
h5psQsdUsGRVegG8CjAWEUyi6XlMVqVSyjFf+qyPjOVVSs1oiMO9jOBI6qRJCD2lCCe2UXKFsEIS
hXv9Q+m15Bj6NEN3mADlqJz/3Y3ylX/dEOIPehSKuqt7FTEQt6hC9EUd9Wty8Lh2oANMeLYgWNUy
LSB0f43+cG2c/387anuG/ARNDz584RPJ4DZ4IpY13Zf5cEJutK5TIlnZPEMWA3xWO1WkQ5npdLZV
B7jructqieq9OpUi+HvBEv6rKN4qubVlzkq89qTlyXm4LYhdWkIt6Ecj/jckYyXN3K97/zbiuupi
uIlnucReoIQOYkUh0+Q2zKZ66qMlh/5VcI/WjTYoJXj4hT6vsntXbc9IfHsHT7Pbd2rwcWAvnygm
MSGXwiRuLF4BNCNa9bbotmjQ3HQGV/kjCy6wU8D2prkG77tOmyaOVqQj/lLWd5LvViqQs4EtjrGu
i92WgM8SfD6lJre8x2nHlt0sZLhP63w3N4tl/F+mvKG/rS3dOMOiLzh+k/UrL6aIOP4ufRdvy196
ZbIZIdsow16a7cRdLPkKA1i+7N3JG11SVMk18wNYqoYZ1pu3ZZKTyICxMqn6Dk9jjBYliCWuMYKF
SQXSQ8mIaCqO2trMV/HRYPQYU8KXIlNeV6CIWaw2vCYFNCajGgeQrBI4albOhC1/BVyxLPer/3fm
NlQn5PGlQGuqhggGb7WJYTpGgGaKP7bMPWvLnMaabVJjwu82b3/9vCIxh9Qigdpgh67HAJt1LHJ2
9qcVP238o8rHlCjFODSAEysFUZ+hNFoSBbjSxMGZUHVRAb1KjEzi+2BkTcu4V4pt0ELmWjYU4liZ
I2mkTX8Qz09b7+EryFC1Q9ZDNWs1JzLicvCMx+kirzVFfz8xNOAksXL+J6OXuC3eD+eAa6xeepV+
uKGbHb6mgPgHpsBFa14CLcSqJMwwGVp14sGVtqAHlwPVK7Jb/nzpMnfctI9SxxK5LQ3CAbq+3djD
DSKMiWClH6nvQ/3uvpVSmivv422qFGhTUbgy1az9YFSf9LLlSKC4cLwZK8TT2Wk2LT574umXMdGW
G5EUfTzW9jO68dCvhK36SfTFCBLJlI+m3fCgYdT1EMWjm/jhOJmRDznSuNDf8EQCdAJE5eMDdhnN
o1CQ1eVgXtJenw/xRCxmVd05fDRFoww6KH6ersCm5YrcIrqDHLsY/KThE7wiQp+loNTIyTf2a27U
ZhLad1Th0VP6wfgqDimejAexUWtVeVRAMLSW8Lw+lGBdWunGEpg05OiVETY9wDzWAX62zgNgRtM1
7sjx3BvlxLmfpp5tLOsm3hrpMhR/gLbVKtgp90S0DCmW5KcVAycklKr54LzylNWFhCz7JG68x2QA
xReG4vFwu/qK8zb1C6NrlW7PcWnUdvF7x++SqxWOdhw6vIEz2doW5r5UqFSS3uCjKtOOhTHam1WF
Yb044b/mxcOAcsMgOxBCRkUfY++ccr5Jq7hUsjO37uBnj0iSgnKqL7mYympi6O+mtYXAAdaHNa3x
kHbaqr7Mqe3K8M/sP3xlSX+irSFMAYTIxzxPYZSgN4tABiOQ0eSXk2hRV5Wte8FPhPFAE4fof6JK
aKg6v6JYelqpyTEga4eE606c9S/nQqLUMQMJI/+6qrGIWvu0m0iABNBjG7RgkaSPEgQZIt60YoN1
E12A0Y0flzp5TFIpSjjA0VsPr3c4egf8VlAzp4ZmSmi2+08y8tdqtpYGEDSA3bQWWjziebKpjdcJ
/jebz9SajGDjRXrEb12nYOg4lmAlUsINw83cZBnw3RGJfnye48MWjf2uzly2QnA6IosUSyocjoGk
vhbD3SmpupUPUvM8AzaoQEpdLchCrLy5DSl3TXjMiT5pfrniOnSJX4Z1wtXKqFwL75RsZLaEjbBj
v5PybxhHk1yT5oVeWxDSigq+W4Lrw47G+jtY1k9HE/JRlbvaW02uDeS9iZ8RQKnp2PNXsvoBAcH8
PoihkgwuUzmoNu1kyKs7mya/S+vteJYyk+3lg8t97DVA0eR8MycWj7bscn+0GlLomDhZcubR2Sep
pUZWingNn/yqZ7e+737qYpxmpu4/+wPCRGsAGZA9QtzcD3Xj3YxtHKKWQIvGEPRSXX2igudgU1oy
llGhD4OMUDrqLA279rri81CoCVYUvEbalhETkvwptyBV5KNSPmPG2FjWcGycr0CGQT+zGNwcKc6o
+vFr8N03bwQCZVrp3ejPNJiqqG+lFWH+0f37Jmzu84wXiuKCtBn638evTV8bRPe8Ew9Xg9Fh6s6T
ZWzSFNWn0fGI33GbBusY5YvbOCeF5M13AK7k06Ky7cTYd7C4bQo5srJJh4nHKk/9m2Ch2EPIkwb4
lRd3ZOPJ6Jx8m7GJMgyLZq9TTAuFrCWEDRZyNW4x2WvmkZCPrrP6oxazFSZ3DgDOPbCqfY49El/3
UgQs+P2QX25Avt3Q9tOJr1L7z5/f14YIor7XjgHmRuAykSs6GPLWXK1mjpndLcvsnxdM+XLmZ7Hs
Og7P2y6z38OkykZw+ZSFG4xpZ9qC0N2JqJymT6rcncjfkfMAH7Xb6aPWsLiC90j90JFKFMEhnOEd
YfTuJru/ZfKZMKqDQ0GcxNH4vtRVNgtp0fc6Ngu3u/mUyBp3P5YYjNXLGDwPNxp9SiXjdGep9M2Z
wDZBmTOs8j4EJtKx2iOr1YnADTipCJOFOCmoe4tXGxcatWvHkYeyW1PETR0mQGjsZ9hS5ZjXSfqN
V9ue6UeyM0mNET77sD6Gi54oyrND2auauWLQiL4blaBfn8/KC32bAdOT+D8qOCxBv1WAwDgt36O5
E55L/lrpgZ0OQL2oy87g5GkTQ0oHCqyqxVR1Wbqe2IRQJNhj7BQZS33OnmvJwPbmwHn8BlpIOjlf
onn50cdXlEvtY1d81p5OxGUc1d4haJD8z30TEvjI5C+99I/vej0eRB2av7pdDD2PXjtMj+2qVDQd
9oEI3dP/cNwH9XVYSNFEjTVLOZyeD7g6j8iAjD8QssDU9eHQ2rhfZf6gz6SnRpoX38DdCgD1ZXNh
OrIYPrd6FxSToKaeboV4S+T5L9Un6jfFHoBYVVSPMPfIw8pZ9QfN1xLubPFMCwNBDyMs2vPXqHxG
3yHcw1aYpD5YHulEwh3TN0d7ZWFh2/Lkcn3r/WP6OtOeGRLOTL0C7p7Uyudihm0wEbTaazaOtNB0
zRLPBhiEwrmIufOSufdgu7lreJPjf9LaQRADqeOlJ6JQYtCycEHwLaFySJVcL4481smT5dvHkxYX
jef2IwSvf7IEHLYVD14U1u/TJOZkt7fUGO9Lj5ezDmb68Lsq0apC9hZ/zfy+y9Dd96HAFvEIm/IR
h9t8Bf7hNL6ZOjcmEuXPqEYjJ1uF7glfpKWvmghodwATNPHAmW3URFNKc6lqEOp1cK7Tux5ItfGL
KBObM8bCVzh/ve9ILpw28EXNvCvWRpMYf7jV3KwfaJ9p6FwaHTThg3R2qAY39EUVOHtpIAwjALhW
pSBOwI3jbRm2jQZ/Llz8+O49eFqyTxctg2MIcWUrxGRKDHYhLTA1PN14H+gLJrRGEeGS+Xh4G/RV
HctW8BFfyOhQ8OnyGKIJVAUM5kfSy4Rc+QrCJIEgOpB3Wdq+K3JMVhEdQSRer2KfWudmZz2S4suq
e0fjuZkXnQI1U4iOL6QGDZ72ZVsVzypgwvPPS7Xw7uzYBvm6Y7VcEBxzh5e/g5zk/3SyuDxsuuew
4sOWi1T7gRbIwponSrjisv99I97m/RLi2AS6Phu95AJqMMOX2uapz0qqj/yDpEsKCMiviZpUqaIH
qccw+iVD/SyR9uEM3tOfFYPE5k0TsdlOPIBbxXCA0CVqtplqd8yZSpEH6sI+nqM1ANYeiPbQM2GK
x4VilaaWxaM8f6Iaj+TBZZZ1c9U9pMbf04+RvQErtHxZ6Nh4042pBaxORfhf7B0OzhqaNH2eCcMi
CpgOwxl3WhcI5dzE5TanNl1bgwsAerjKV0Yc8Gpk9q1OYg9u8GKsNIrShriBsoS4SB0k2IzoyBtI
6rIWoD1jSklXE/WtXVLon9ZXFpx6uStxzsRkPLPLTSjaMajx0+ILHVrorrhGWVgIl69eINl9fvr2
9SYWx9Wt/3BqHmltOAeZ/Qo9+EmQ1HAkhXjs0OPYxGVVZxdAZ/deOgtsXDNgXIx69rpS9kcC7V4/
LLNAss9/zCU1ytwt0mRrqT1e91GdvYgSW4Toz7AW4PRBh+jweI9ijxkJlCede9ynO+uW/RpInf0N
MUnGgQZEiOK6Tp7Uk0Ey98Fjdf3ksI1MYxNpVq3r1xx6th8SMh0Jxzpfe8UsdcOzIF/z9m3mj7+F
eMoVeEt7R2lGJhb2KNYpu0217tPMfoWj4/9W3d4YJW4tXr5O23EohoAj5uPHQpaNggIOiMGfHcOH
QW/ehIz3eZrWoqBQ4YUNyg/QQAKR4jQqP94whyBaZiIAbHyPhHiAgZqH2LVgqbY8jroGfinMVJuI
rZVVaCuhLKwUqTJCr0+Ccnos59W2HSAArbu8rLkRjymMDl6CoGleWQASzeFoZIwefCywgJCcW3jL
e2xEvhiXl9Sny8c1YjWJKrMjT69j+MTEnXT4l12XHG6ZsMBKunT1kyfk/Uwi6rKz8rEyEt4UgTkh
WKY+Xy3uDGyf/927SnQ9pzWDqKiadaf62KdXTjm3/Rv/QbuBw2O/xUpFgmRZBcklCl0k+y8rFVNe
qEbMaUGwLHzkgfPc2vverctSaPsL/+lxoRjnBhwrvx6foUnM2uf2wyvvI/jYI4BUfEER40OWEGGP
Ujlp8jUASpIzPL29czKSEMD+BCuckoh8B594glSf5UZOZRSZ53l87z4j2ntuSSW+tpcTUTj7Ljia
ymlqAMF9NL48LVcVosNS5pI9OiVmAQiCtVUxjnGBDL9YMsHu5tvrV4vOfqxFAXVJQP0CeJkUbfPd
lfPwdw0eZpRnF8wWfG1vmRaI69GR5IFFjHbdrjQWxrZ16WWg4Iq0YEVePhlFF3c1ty4W3BLbSn9b
X+N8EnMZ3opLSYJkg6f60h/TJzTMzONfIzobns4z0IQgI4amhHilr6R9hPbP3yEHXQLNfxbMR9fw
uCLAcbejYedn2B4INTHm5Y5diZa94a11z92Zn9aFh88KwHnkSNgrAfsE4KoQGYGcRAQdqurS72pB
YCNbloqCDjGXRS+4c4bOia/x8x65ANjBvoFQVPax9btedhgttgkdIaKLjY5KyMLUEDhaejvnxYBy
zZ/+wpKDKxRJM30tnnBwkiQmWCLWx3RlyIRR6F8lKCP3r5548q+yctx2Kcri9dLHfvNGvyLLks4G
uZWjMwXWJCtGNi5O3+QpC2D7m1wmVuYAraKKcIFWiwLklcpX22HkeSe0p/rQOi17jYWrJ9yctvpH
WoDZKPB97dNff9inNffOpm0o4/JYrKoaFxRNPugiJt7i82V1oiA50iZlTxJ7+elXtjfPzVqb6Rxw
MoGFcK2e/9Hj79K25dzdZgHqCcf1zRUuTEj4WVlKRUD4/luXXBxFnisiSsze6L+GXg5OoL/nHXdZ
2qQf0wtCy6EZd1h4wGgUceQwMcpcUACQgCNslkReFrXWY7wcpk6Tsu4YE/XOWN7WBdny9rZeWez1
zOK8hWLIGrPxh1LYU0f3qbnECPbmp4Xur6zsan/ZUkyfE0aMTg1e/mFre+JbyEexORcCnyqajKob
90AYS0EFOtjggNaLrjCWZER62TKpeqLfUKoXkfrdrwDjerpSgKbxnMh0st4BAXl5ECshRkBAOfXJ
VbdwR+d11UCOIzmEd5tbFQRVEI3TH1TAOTW+vKiyMOK3CfZgM0dZFv1GmN5S5Rez2MTjnVrXtAWj
FR7+KH/dHclcsrRz0hGrVfnJgjzNk13g9ABXjdhopFRpjk1fq0KVUuhAA8FPsLZ360RguFtKDSgV
PZYkDCbtrnC3mxssGSwHTq2hTsDKBBE3pWzKbfe5Q8+EblGKpN4QIIatiqF4RMDpaZ24RzYdnvUf
mYjdaJoQC/jSD0Dj+cnShC3P2w6HKMvkinAwN3BQmiHIfDOpmbY55+Qyj33ilCaR9ZMiNPAJ1YrO
hPjxSipumPsAFdOUeDPCcOUBvELAtuwMMdy8kUNkkpyM0cGbru25AtWCqcdRhfUK7s2qEBbgZaxz
hYOZnvxm/m6Qn+EP0PLMQzxa8OldFLb+OSP866TX9vQrNincrsqgyu+bMvAAnZiWAh5jDRlDZvBR
6jtE8ASdbq6ZdPQ5x8411fYLQIgffT6k+xEz6bpU6pTDOOXfixemAa7orTfQxVx/E7E0qWtdpmwi
lvYoplF52C0yjnHbKtuI7PraasqcDOI+PyFtMJ0W8420zV33gaGjYa/tyqIQB9qPsxFc/GvQC4+Y
0wu+AyV8qbDLegr8woNMhsGKALRW8Q8dffmiqns1JO+eF7QomlNesYRIb4H4xbvKRCEqkWs+djb+
CkNlW9G5Z24vTBX0jflbQ/BRyJnKYOZSlcigBP1juHPQZJKOftJd3c2zIRBNfdiLnP8wB2UtlNz1
NZSjHmdWyswLJg6xCWezcH6sSXD4eF+ADw5zeC3/X+clJA+LTAa5uj69nT4nnQ/no4FqsNkMyoDt
+pE98dhe0xlzzPo38hNuMH/79J6j25yl+H3gYdz2/uJgcR5GR7s3OxFgvtaINkPya5eZMe1sMU5L
e9Cm486svWcdRbaIO8z4PbLHpMxBu29WzokbfisJguLtOi8eHsvhFj34V9HP3f5J2IbkJr3afuIe
1vKhES4ynF2RO/wCFY9LhUtLpzDUBuQR6n1kBtwQSussoAqGHkveZxiHsg+IQkNTN4xEbzz+pR7w
8N7+2E1iIB9p4oI7bbpkUpT6G/xTsHJO3AMlXXsae/lkLpbOPvNueZDJHzkm0piu+YJu/W6Rq9hd
TBk4xj4FwPPQXcDA+nLur0p1xseqQ73DR4BkO3rY0GsOgjTEhfdJpKxgcT5zDeuN3pygHEK5m1Mh
FDO3NFLxjBpobJPgdTCQhWGPz4AYrQMoQqDeFxAatFxOJv3VhPlFMkVrtOWBU5Wxef6Ui1v46QNV
Z3J84enn8rp27RpYMhoJZ7wLHhdw4Z7G1cgOZZ2SyfuqMOKWvgvft88dXsVWRGJDJNvunfweAz6D
li8RzSSGjyfP3dB+l/C5TPO4ZzlblTN37mC5fC56KAm7MeKTU6bMyZZuNgAUTICrulUONdUMjANY
/WBAu52/Jfw9cl2hhtxlgqsYWbVOOhwxXdq97sAziWdfu1ftdOKlv8wjYh2B21l1y6tAhHyQPok6
+dHxCQvvpTQX5C/5QPsd6VHA0zs0Ku2BC2oQkH5OmYv3JTVHS/hmunxOLFNCykBDIabOJez/KM2x
H4Li1ejUAgx/3zIsKIEWSMaoGke85YceQ61suKeQQC7foQRg3ldWCL4fFmFD0fLfcY0X47nCJsGo
LOB1eWGXco9qkNsogaJjWo2g13ho0TMxEzLTGuT9Lov+n4oOQEP0gWuhpi+Ws2zh98nhYKxaTSEb
U+InLMhFusjx2wibTE6fqObt8BeRJbcNaJC0ckTJgkmGPuycimoZL/gmMpQ2dhvN54sskewIG9i+
t6GTgv+85UjnWJHPaS9lemdkm00MWaZPhZOkkLXQ9liqT10Kc39NR3CQixSm79UczGN3n3EYoBrs
w9kMNwdbDg0tN49lltA7DRQMmo9kRr4Ja3xX5+7H996XIIOGbGB199AEpyTggVcPkfVeGABSNwGN
NnVZdN956ZRtX5mKi9vrynzxvM03o/n0OgqEoz7+p239RsYuiFM/mvRx0RV85MvKyIDFui0lSOYu
sm5ZikH5sxcPb7/TSZohEeIkUCJMZI72n/tmx5duL61bA6IZTQtJJhp4M6X2bQOJ2Lo4QQoa59b3
a0iddn4r6vhB27MFHAx16tx44reVBEVb4iDSWEVEeu3ChkOETlnEjI955gR69hCxB/R2avzmB2/h
wgM1sM1rJ2OZVFLhhtN5R3OvDnjOeNbOKWWZ2R3FlYV0EErwGfdPRLFKnZF/VMfEkBbsjjXaHdWr
UaEn+pVVbPj4Z2/SWGukUtzRgZDSpzJeg/n+3kzkbebG1Udp/0nUUX32Ko/GqqbFS1bi/VMnr/Rq
ef2g3lgQCUzE01zQcpSTO1+tGkkBg5emcNkdF1hqY27XDjeqdXmH2kAi/sCGTGez5AgVpKBUAAfa
eqirR5arnW7GLiAmKvyoQ/MkXwwQQyLeZ4OgTZ2EiZrsIOS7kGJetDiPPlD7vWBixYuEnJtRYeKV
0TL22onmd8rh6MwY0Nl3lMGdm7728OrfGMtYQofY78o8T0NCwDBvh7l+NxU6pa4sEZSzdDPOtY3Z
XGm1e+wmKQuHRy8dQeSxhXeknoucNFzQ/JiOsTNBZqTJcpzantY4HmQGESDY0fHWMcbIyHIF+Td2
A9MdBZR9scNzcSx3MpSg7bnuyWHKyrJUt2mGs3zmxk5UOfrATLBgyYyCMCUhqtDPITCwx/Js80KD
hBZiz+BGqCg1lgOvI8xcsPgUDBjJefXA+wrOBZI4uL7+zNfzQDNtqQtjgvSuXQUnXAfzeXQV4Vqg
aHpDijQyg0VYWmO6LpmIkiafpiaChJd8fJROZJtSTG4FHdsVdY38GUfTAB6oun8EZVv5ZsEwd4kR
0+IKlUhP054IO9UMg1lv7KTzkBy2lkuULhdL8Xhmu5GxduxL8+ZYIGPzmwyLNdZnA3AX0frOijhQ
EwgtrUd/hLsbYFvqJnoWV1lIs2v7J+xXwiCQTTM+URgSEgpQJncBc+1DcxWeXWGo+aP7V7WWcT8O
I6kOq/+VP5S8O1jOow0rGzhjjXm39+pp5GoVkmWD4PyO2B2b4DVd2PCPZIGvFWfanQWLlC83eJHl
7uiicl/sLCBWRYE4Nrd2v+vIfk2AyZfVGq+lYrWrJLpghQN276+s8SZ3oCYZCR3dpUIE6yUwmJAD
P1eua86C+VxvuE5gO+PO6orzykZZFof49Y8ot1HwEO/XdzZH1MKd9XQWZurdHrkRcKeDOpSCvRtQ
f4hYyouNlWoKUn7HZEWjJlFHHY0esWxarOCjd4CzLFZMGiFX95s/oI3F+6L1BfcbqJkcz2fzKByY
IDJGdy2fj/6Dnxi/pSH0wazrt+2RjxM5ySEMJhnA6JeRAOffOYqcY660jut0ndu32oxqTzbecMM3
l6mrdT/MUhLyisb5xUlIktXtSQ0cs43QlAR2tEKDCRXAOgbG0hFBfR/QVkeBifZnlnqFlGStdg6g
Ve4N4tkZI6XH77qHV441m5TpF+VvULRb6c3mAFptIHBZLELBwFdsVOlM+zTVy98IjDJMQ5LKRyae
hr6WHlIUNgz76gZhR/zOhQpd+FvV5LkvVXHQDsXUU6GVrm2PCzyK8xKkyCFHbvk9CnPXkAM+wDEK
wFU1UgeL2h4VKJCszpQL7kWyVf4/BrWIuC1J4tvXXuc9ofepkeClAaUx8xyG2g0QLR/MWV3dGjo1
S3Q8gVO14nIbwenAEOIL2ZwdFDgx9T+A85y+MfvrwUzSXV+jtCyVpBUMHvwlCAlQ7zuEAfVVLICH
CSKeiCWxxmX5ahzZseyPH4xYhNI8Wbgw/tfNjJEFmlxm3x2nr+h5GTwTzwJtvw+eLoSAiV4Sgaeh
zY5RtP52yusWKjNqja4QpFvyuwjy4mld83KoxapC50KdCZkBdTFJNmIiEGEC1cfgnCQGBf6d7UJp
609Ge1+bEYsz+olC/JnviP5h2AV7PjRv/gN5wRK7KJ3RKCm09I67fw6koQWm5WGSABGxynEcIUlU
XptrjmCkmdgjGmEKIL0jxiQHpGH9uH+7LBF8Uhhi1Te8XJ+fMYPJkcKJVwTmlX4oWlWY1r70mX5L
ZBgfJ6Vty5fkjpiLmN1OH+5UbZYD1PQnAvA53bBZpCoIiO90eN0jZLbrV/H3yihAju2kYEGmw6d6
DGs5tlSukVDP+8OkH+CnZv7/YmmrJt8v0frc/9buSi7M/Zhe6C9liit69K5YzHowLKqnwb6Bgqy0
hDvzq3mWVQPcyC8h7Ng2OV46pfVofTFK82FSAC+o2Z63M6IwnA5YS0JWQSgionBai0PJTrY7C8ey
h+Rh6UU/yjueocSJoFAnRqjE1eoIyQp+Rj5SwnwNxuYHFwPZ2Ry3DoPhM091S919GPAO5Xm8wzhb
kSXFNiTU9sjdd+Wf4Kfikx8Fh9C2kfKZi/tesfTWPpB401Q02B9YHpSAF1XH/CCVECgjqeS092Mp
9MjYUo5CBofBKdWYDiqAQXgG98Zvbr3AdjsjbLnXSwOoh6yS/bHLEveMdjIFuBtuCOURIdc2s+hK
dwveiHWsO63xtTk4HIqE2wB7zH4kL1kbse8Q3kfDX7QOV5ktIUL64/mTbpsrAbrEf2W5lGwZXy/d
30MxRHS98u2kc9jXhhWIrNxrOXx/++cU5sDMWoMl25G81TyDYjuIJd0BjaJeyBieHY8GN/EHyHTq
5yXSQZjWW1DoD0Rm1Q/dlZ6pwMbJKtuCO/FdLPcfZzm+EPyJvu9p8deXkxV3Ai0mDLvx6NXd5oDX
HseMPJwNvEYhVVsoGYiIYxVAl/nfwjdtt4Yijp72lnwSfp3sqQh9DBHHCfHXdKTVlcmYAVSKatuE
SUslP4cAZ5D3w3AWVh0jvvfZv0YYsHHvAtoMKklWuDAnBZ2bYOKNerm8YPFzzWTT2NscyjkLPX4q
YOowwCRKbDR8lVi2vljAWyx0XKVFCFNTAlpRHCaQhgrVjBkmNVUu0IaCz9qV7YOCf0/WXTuDnldo
SPAxa9QtpzHDzVV1d+4ncHd1vZiN3GmfPEec+FxIN9KDq5Rp0r7gF3+b+qfjQ68rQrBn23FpCYFZ
wOHtGdDzwsBDH82wdekhGYUzWSdMbrxNhgfzu7YaDehLQrgHkfnb7UeO2DPMMW+aKpO5A4Yr2+VG
kSJtQuCmBYObczV9NRHD3QH4yY0ESRQ23hGbQbyXJuJ2hGAuFI5SwRtLJAY6qSJOBETlolKIRyYC
PRLbDZ6wc0oblJS+sgSXTR9Hr0V4RELasCnpuxzpRfe5rGYcGx5K3sQtNm2EZWvXVbyOV4dEqOLV
XiJOYPpygsh8pzTvO3OCixpUCG5PjIGO/ByHQ6Bii20CVR/7o3arLoXEWs1QD0ciABofzH/UmM2k
kv8kukfuUoxmllLKTn+VIcEKOUQ4ksb8f3L+hZh3QVqdnua/8sa2w8ByR9nHxTkZqSUG4Qq+GIMv
DD4+DQZegzdkaf6yqjhoCiGHf8kL/8+fi7jg6Xga19XI2EQDr1G2zaxxy2+rJJv9YBn0x3AsfPbx
wakb0QZQ1X6Zaf9jdYgCbIIIlKlpJeYvuoJIe5CVf/LqR+vRJ6aitqJ5hVlOo64UytmKY1ptvzoh
GEz6YkUSt8fyy0cqI6auRgHFnhlw2rzXicW6PmETBOMadE3+fTqA18ZnjDfY5vAdgphPkPnWuG4E
hE8+QKQkj3GubwJwoivoamhLZoAMZlltLUokkuAJHhp3cI8BwB6RYNCOmMWbl2oAZ0QJ5rkShQwc
IleXeyUZbhNONikpAo3bZRlVoIrNfswaifeyXlIzSyQ+8WK/s7UTdp+TFHsYzaIjmPd5AgCgA7U7
Q1+JQ+DBjnGvVp9mOWAEyb/TjVLxyulOrEc61A2VzwnOgzAJPiLP9BOmu+WwZzGpa6EVE4gNASWf
T6Jv8YVSN7+RItidpMAxysNhbaskpp7UzE07mZf07e+gUdZzRqI4aEnsku6Ho/gevlh9Quhzb2o0
q5PSNroJaWFkhYIg4nHnisIpG6k0qnN88xD0UNGMhb4LMFK7Jwsk4dgHAqWgpf1KPHFfc/a3Hmlw
V+yktQD+Cur36PNbrvxF5qflWwzxwDOcW3LjuQX+fksic+7gdnIpKRQ2k0sMvwCfXdJZkjQ9/DJ0
S9WG2ipf0Li7jozLM3B8NaXd5CAC+/XxDMoU+suT5qYzI/q+8c0sQ+g6haydG2BTIOMS8I7ZSH22
gJJEaN1hhcBNl6LO8NtI3eNKd8BQx8eOqRPbv1/jf3+mRbmXIKld/SJzTq92Wm+ToPW7Kcd2ziTr
IEFtcGQJTz/vjXghbJHNwcMa/HoAUVB8RDEuLgpZiMzmBerYHDRh0kNe1E3OxifhQJ9Cz/YUabmU
j7/8maKJNu4zfKOod282zjtbNUucwkeyWjhr3vl7v1Z1biPSQTFGHhF0uwlltC5/0k3FNy5yI47O
8DZzWikhkie8gMwwfMbAU7ilo/UsFeyIGSgBiuHStCv9KgRjUkaog7H9dIR+1IoApbkEAF+V6AQA
sDmYcfNslECCO5ycm9xYjXh0h/mPezivN3SmCsMovcFzY1L6SaRfuIYBVasHLeZyhMyXTaLzLWHS
/I0YV6zamd9PuerbZmY1Lk2nY9v4etqfHTdtUcoTMYVIeUSsmBZg2yHQc6dOmBdoDdrKMabjzH/w
FOpFFaNQk81pHBf3rAjXKVxn1SGiWZtbA+hJeEyc4Ut6qIfN7L65n5gJb9AD944x2jEi45C8bjFT
DGFvgl0hghckajzyx6PV4J0AcnysuNnRu7X+hM9jtuyApO3skfWz7DoZCQQ9FO3qDiT1sWqhPTnc
nBqE1rVtRsWa0Nu6F2S/GPVCjf90frtuYPIv4Pv+/Zxl5S7PvTbUTgviCohvO4h30ug+uJwivLMe
R7KDVI0bYYfSkggFgYFCyjRncv/W7DN9LtO4LZPX/5T/1Zz+KpytbsOQFmRqg9yOQsePgokgf9+Y
iTN/+520sR12pFt+9kS5F6GR2o0/irqC1XdUQ5FhCA/Hn1ggsu0s3jOpzk/9sVbkYMfJPmRW2Or1
61tfmJ3Zxf8OwBPBidE+vwC1d6iO3tScTm/Fm5E78csOKc+axgT35Iap2+isktwCS/wraJ55UL6L
GcEjUMxTJZnHIyRKw6ptiEzlsGmkJ0AdOXkjNVafHuvT66qU3aK/aAn6kNQSu0cuWnYX/EW4MmIx
7K1JcBIfLyvf90onPVMH3ay7yNhKxSucwSGBFYRRKRB/B9cPlKTtXK31h/djT7dSBACaxeswN8cW
5N/ZYx7i95KOjaHml9IX43hEZB91Ro/XsKer5hJbAdjSg//fDXjYx4O7X+gU5kfkU5IS1q4E2KzZ
gCVT7n6J90CRd858A6uiVdzaydLoWoQptMovv3hue/4tW7GAbfKeqLEgjS1bc5Jy/bElkHeoyBvh
S1LKniW7U8iN0ovMZswH9MAN+17VyoOzZtPrZJSWaTVeC6sVu/xhS5N2/Kd2lEFDq61jKXfqmWXs
XK29j2qMajK6WYSLrfid2EA/fm75xBFFA3uIYL+aLvS/1+F7H4oqmIP2q8zxZu3Z9jWXxndZqJez
GHs37ULGYEIfkl36W0hcvkC+CmnC5SLiC+x518mps1GOH/VH8mRa2DILz9OQsRc1+mW1tc978bbS
r+9U9Rs0kJmj6qZ4cxTAaUaoYv5pde1SExCgjOe502paeVyv4VYZidreAKOZMudnPjHe1TBFw3Hh
YJE4C60SsL4uG2NhK/CmCfnFw/dpfShG0S5BIAjsuvBRk+vag8RRT+rdJBUyy5rxA2p1LaHhNGei
vlHVw+P5xW6W9zzCjcAIaSiw8GK98Bd2kT/3xbbQDcPIa4HPfy71tktkK1GJLkcHz361uPdWIJ1p
8GMxItn0CmHLd3TmQfOiFwcX4dW+cXo+gfFx9mdOr7UY6/MKkuLSYviS/NAVsCaJcc3dq27doW4H
IWYA1EV1HSHFjFfoQ/p4dlbI+OqZnVNdadlafEsneStvHTWgpYcCn9ddbW0QYTPSkQ5dRuz1YGfm
ocwhAW3Oo/6ZiwpL2zuLttjJO8WzewYmCOySPUtTaicvhThm9bqso+Hv4WmIu2aPzmQGzorfAvtH
WKM/LAUPAuHoPYtHnVWB2V4bEqauQczq/aLakYTWW2T2q8lGUfUsf3QkL7OXuae+asyIXx6XxeFJ
jofspU05T2I+OuHO2+zcG5OcuNRdydqSsD2aJdtIzD7AuqM2wFcsCqZPp/geBpo0UFeUoQUfSUv4
vEjj6LcmkoxhF5+75gJcfbzAqqKcaGtiSDXEkzIxOAzIJ2QziiXbIQo5gPUbLafIbmhDnI0/iFiw
8ee28DdzyES85r+ARZ+kEB7XeJuDvuYOpgSNdJk89K9jLRKpnCB6sqG9GZqsaAeDhQiAV3AODzBL
wNw8JXpWspzwHAi8fZcUa0gWNHoLQ6XRn7MsCxq+TJQKX42sh3I7e5vfoQgsnGuk1q9vYzJ0OdM4
Anpjr7gEOax+yO9cmEj0gyurfmF3XBnTIK+AnfZ9Zd3P+xLC0TpZAzLzflu7gmSqgscdhuMK/jhB
/cqlJ8Rs6Ixu0wC1tMScUlXWOkd4DbuvdYE0E2dzk/6xf8MC94B58xLSeDb3B3/CTYaRPZ5epLgt
QtRvYK66acjJkVrWbB4+wBBwH6xb2qbztrVIS7iY4JWbqIpnKG7bH9pHluTOZ9MmsKF7P5zi3EGy
w4OjZQEvszKjL2x8wi3BW4hje3aDPwodzW/1D/CT4Z1ybGPyem0RvJ2CPqM4iaTLhuTuFNS+tAPm
sHg5VECvf5ZCrGyv/kPn0fQgxWhMVUj3OItY/Io3HKs5CiffInGY/FK2AAdRXbalZ/LP+50p8vIx
XYUSU/bwiPPqAF+JtWkayHHGCI8NIw4RHci+OE+a3aXYMaK1/FtAHUhkeR4kjLQ7JBujLD2SsAVC
CTNAGL8uysSkJxM2nACxypzWDW8Yh91TqE60S/KPAkXxJeLmmqby5iydpmApUUHgfxIwimlB+dfs
K1GcVkZMpfDeSMWliNrFiGnpuMrc36WIUxTTkYjOqTOIDIbM4PRL5pb9FJ6FMICTB8npmNa/LtaD
Z298CfigxJEbsKl6rKTecdVkbqBLRSHxEH6TviDmVaM3zT2+8ZZAvwNpKVQZgNJEKIKPkc1TLUmw
6h4mdFaa+i5hRoU1S/YAWFEkFXrnF6iZ8rT6aoR8j9oSyk+yE3Sr9+s09XTw9SLmzt9QS3O2cy5U
w8o+5IUKJK5TRGYAkQMf3Qrhg9L0J0eV6AY1cjRcZwjDByk+EhKWj2vOpvOmDZUCFxmKSb3d0IuO
ZgO5xE16fGhVFkNagsA0yeSEH7r9yZ3b3/w8pc30Zb4b8t2nWdPBCDJRJRgzBtqiF0vrN+CbSqjm
9N6LZ0ybR1Bm/cJStAtXwekcoO/rQstcZuRpgjBklLFxssbya00AxugvBct9128hzw8e2qF78mRB
AplSAn2Om6RDBJuVSSFrQx8V9AtTN0Mmwc6Dh5vG70KVijT34DRZhtv4O/xn4wEIBtMqMUq/RW9i
1Aeqn4WFZNPqR0Z6GV5jXA/egp/JbMfKUxDgT3wPo7ySxCneNqbyhm013IV8rlqQbx8pEczGdods
sJFX7delbFVgwBhgttx+QCweOLIKK1vXggbofrDCRMzXZSBNaUOxVLdF2BX2771EP2l+YoGpliGE
8Z9kRPwcIY7Eqw1TTbnShIwvb4INN7mYxziBqv/G/JYmnmHQv94yuFQLM7LdUuH8gP4ut/9n2Yxz
CO9aSoH92Nd1ntOhrcV14zRJYypVQquervVtutY0GaSiGH3L7pytmD1I6UTAHgVbf7slGmQ5Cbgi
QDqEzRbzPmkoTS9B7VZlnIBYqZIvy6+QsBBRQno3rTGUb4VubtqxNIkJoes6kWfZNvVJcMh2Slp/
AwWPTSRDMzWrasHY/tRZn4b/1P24T3KP2QEj7Bu1DZxDaIgEZEMb7ARsoSzVAqJJAiMuA0Rc15EU
Xz3sZBLXtNTLUx+BlzVFQSDSru7ZyZkqGLBMbGxrim2JW62vmHmjuTAQodhEjpa3ipSbvLAde8/y
67OYxuHC7rOi3uqsMPXXUVVr3JNKQ8mFcK6DqkHOOYbNpijcrDdIzuNniVsbCQ26aSpnzejsf6gC
jsXqGxG8nMF6rq1ktDBzswaqdE/WFxxxhDkUDiaTpAytFsMVdgOtMYlyg1mXVXf+FFDad8SugS2P
tPyL4MR1xWxv2bT7PeAclYyPZRBJBc4QoBRFarl/uEDlgJ2wz3WwRYnQmcqcBf8sFkXUBssTnr5v
7htUyul9SN3q2ZPl3iO3dAiTBGV9BLCMweBFeLH90lRy348vyTUYPaQkWBGgLKvNJxUkC40EXTCp
EaJiTwvpjr0SjMqRjr7jwWlalxGKza+pgVREMdlzMXJXCA9V7mcGxPKkMoUyLdxG8TC8+EyAYibo
XBlLaJYW6jslMHKofljCWVG2SV2sNTDNVP/DYAqYnx8OTXaWMXjDzJe/ADjLhZcw93eNOAsfxkcm
PI5TwBcsyoN3H6gHBlMNpU4rBQ0k4qaEEoIAIfXf3CC8ei8d7ju/y6q1Y3eSQS+jCsmiP4gPFGsX
Wh1kQlLQAiIidD9XKyrVvR41oL1NokdpDqGQZLO/cE/Azz7iObSMBbrLJ5Y0/EY/+/xIll2OSzWr
n3uHsVuZGqK+TSZUkQFAMaXffnYIlv/DU94g9KtZdYVlMZGcLlCYBYgKWN6XQZMfRB2eRA9OEmZB
OagPE5ttv76TQ+j2so3VxX6wwQNc5+46TfDskVo2AyURe7oOPQPu/OCPK1BInwYQhLq2SO0g8xU/
3GP3T/5ep3IQfkMGRJE7Rd2h2MR9hr1KJwWANv7r+HuXIX/4MC+HZWCNAFusPqLVs8eEigTMu2fe
5JdF5tsGC4gGLAyFBTpaLNA64Q3sxB/I3AFETavsDErkRl/nvOuKlE+DSINrO2F/NWsvH7XHbwGD
B+2zon3G0NcBWuDmpC+95ijC3uUNHpgjeCGubdXd+/+yMP2iVty3wT8t7nPKlNpN3/sFkPKVW50O
oAyzDjZTMpnhd+HTkfBUHTmeqDKFO5XNBcfb/wjY3IHmxtMVTM+EhpVcjfQg4FDfoSq+fRsqpCJV
D/PYv4jVnnAxfgiPzLYQ9XnRTGNsAE7y/2O/lOEdr7oOfmbV9jJpND02vYSAmwTKUOSqDaZmtjCY
FKPdIFGo+CAbf/ThIREOiuBOYYtTT2yK1DSSn6rkmJ8/eJM7efyyU2EFiRD2Hrox3z4qBJSxRzWy
Ngy23IeN/r2/DuqZGdW6/4kKR+CjJ0aLqKqkm3trpT7Xf0tGIvxuiYYGj0tEEgKchjsqjmagAkUq
fbJiecIdjkzTKI52fJN4PPQwE72TUiornCvN9j4qAjtDfzD4uM0XXGJu9PXNKacxzld59M7zCM0y
LCxoMl/y93jwORK6lJQd8dgRCcVjdf5qVHacSZ6QGTz2cbltuE3j2o3z63YQUo+C+tGfx57AGEq0
61Ld7eysNAqAhhqZZI2UcXzyHmcbnJuQt254bITw35MvHg9EjPma9kSZO7VJsRafvh2yEMUNB5Z6
CgPmYCgU2ariZfcP89YFS7JzeAaIPS82XjwaSbGRIutQw3r+nMRdGwQz+kNDTZDUJg3vLzuSSkg5
ohl2gEUgYeQLR9emfWX0xUgTN6uB6EWxPhXLRFQR/VNqMWdPJPMdwQkwd/pH5clMt/VCu+xVbhli
b0bBtmx4uM9XpbnJTiee8ITJmeI0lWXDEdDdYHUfp1gP18temeHGKuouPyPW1OyaZYcQn6ZwdLzx
cTaLiRyYPs8VaVoSjYQ+1BvQCl21mknp85vRMDPSeFryFGWtiEPDJjErmb8qTS9XcRkIH1Fr1lc8
A9NNsUiv5ZK/hZgOP2/UIeKXrlckZfPYKnzgKaEB2/iz+C2XZf4IC8d+gk8PQL1lUw02+G9EaKEN
JwyQWKf/ChpA9yGQnvMIim7dGNNQBmiUFdS8Fhj9ZRZGx3YdRw/fR2LqkxObnIa5hcq8OC8DPKaS
j0GANFjnxVYu+laxx8YHsAA0UWSq7wK9jNG/zJxETxSAoa44rIOjCwy6KbJFKh/ziRWOBwsHWyNf
YKMlAxXRBr7jtuqYS1YNOo3Ab8jFYWOPYpRDH9o2SStkQK550kNm2tX8Qow0f8L/MGiS4dcI4qoV
CFD8HCgaU60rdIgyoBxZjTm4SBT6dJ+k6rnclE1CUSOcV9zZIQBHaYTOgmvMSYtxrsJeH2wI16Wm
mAzClFmTVcrrJJPwiAO5ZgLtb42oAJxU1Ozu7NnDz1CCjFDj1glNJi1Lqf/hE1ichvZl8rrIH03m
MmJEcsxw+FXUvdbcXLMCDNVSRyDeoeqwrOS060HZph+gqxfbnkj5uk88b7hu7HoxsMsJjnBtvSIG
7LYNKBvD0QFTLC01x+ahSblfS89TpaEGxc274/Nuo+m7c11fiOzssT+vVmcCq3jdMtsQkkNvIOcW
o6RcyK+tGrYApC7X9XnDEO1u6GX8NS5r1m/QnqFm+bFm7T78xWPdfsEzx5yjtQiIm676XZRZSPFe
YpeGOxJQDxoKS2LaN09HyXVWoWxt/V8ZymWN3Vl7Ebud6N//+IVRyfwqnMRxYewzzlyaOqEyhnji
gAe46ziVBw/XaVLGqfO4atSQ5X214TPq7q9Sr299a1IjDhc6A3K5AX2tCSiITVh82mEz1QuYekLM
0pt7YUzcJgaPx1JVtzw12fQ/HMwyEEN7wFVJ0pwFlfiOWa1gs38PMGJKG8VZT8SMPlNt7E/FfpzB
oxDWZ3lHvg5h1cqekSPOa8VI/VFO7MF0MfYK4gEh+T5zLjJqtctPGnX9QBjui+hRle/xGc8bByJc
8M2MdIHX5XjietlaZee+jHBh/CLIG+mDaGZ3rxJ8nx87jleILIYxYKNTGYdha3hhrqVt3cdVno2I
mAehrhoEqAJViatx0/U67wf4EbEsJd4341TmYcJLBCWuC+IEu6Lq1DwkqLaDfB8gQ/I/L8ABK1cp
9pTbNBFw8zCgP54+4RavV6zKdeW8fNZsdL4SPTrLYEiRJRD+X20rf+yCHBbcAXVFXhij4bUeToSV
dJr97USw5Dxw6DDxE9o3RyOhgpTti9fJGtzKk3biyLytbnjqsqIPOnKGwGsZplpzxQV4Kxz5aV2G
JKGyY3Bl33TW0T1D36r4FVADx7Y63xhML7GOkmM5lOUZ9T9/Y6pVvJmNnrtqV0Xb1jAVlHzNnMUL
390z02DYwgUBsFCDB0cf3D1xDesA8BgHQHJitM1rk1GeGprZzv5kavpu9jGf+w0x9UXiJuImBg3+
RJQocaeGR/uVWWh9Vdb1kmPAFjVWtyVCh2+YPdT4RKuxLHMH262r+LiIkDeONRGQxpLBjcyMGamU
Fj+jVEampBXghDo21mSddn4nQlypK4EULNgaK5tZQaUcnMnX6LizHgX8tZwTmvru4CPw6oVA6VB0
JIfblwRN2BDcRNtOLjdKhiq7pYaqY4nA9if5VLfc9UKWBdhqnRdL/1ztTv/t5Ya5u5q/LVDOjGRv
45hNBLY4HWo2BUp5Ds/skuGTKMY2n94SDr22I0yrXUBAwIxctbccqgXa/Myu24M07Fa5caBbSn8w
p1Wz4w4O007uoZgb76gwnebad+bG3RwpV5cJkief3Qfyy6o96kT7Nrv2bS2S1KxwlJEZmkftg78m
u1SS2E9BgUIs9p2MBZ+c5WIi2n6LBSB5wgTehdigD3bS+LVnf8G8hDz0O23GyWeey/HRFAiK2Mik
a+cdDkg//JBO9IUrXI8Ls5mihIHTigueY4HGCaRHTVkI5LOGvc4ROhJMl+llTSL85KPNYwAEUVdJ
umq3+Komq2svH2C8zGXGHZCp0NIGxgspdQnv2UaTZmbDaARzN5z+ohI0V3OYG6bU+sa4LP3OfYSY
gB1rvOaHywUMzHriousTtePeEk0KhrcSW2Rdi9dzdvI2tP4R5bhQ7zAQjQjpsVQ9FZQBenR5ME/B
NbcATTfCsRqErlGzIIe133RhTYRnrUiuExxodSZbEwlMbvHRYVYA/BXEEutFo8ZQTEIpwOgNJll6
Emt0O8vfC0YYZi5jlqqro4Olub4mbHw0bzW//zyHPRsB4viAruADr62aWa3KHAen2q2hvJRgq9AG
5M9/6vm/5VrhKStQR40kw5q8fciSf9lrS3mtjcfKZ+Z4qNQig4OMh1rqUQH/t1uWkHW+4aEgFOYp
6Zt+3rZxh4thOkkOsf8bxf56BlpHDSh6ALgMf/fr1vWwimoYpkosuZjOZRtmHNusVP4kP9PJUFHX
2COUQ9Fw3Tn48nS1NHAjqvT4+xoOyUyJXCCL5QuvtSV4IralyCFV3aOVI6afaABrd6VFKxUNCXHm
OozkEWixUDR4kd9n7m25vUhhYcqzlzMnRKFrp7BHf2EGdMCMHM1olkaOrmg5cNBA+Vplt3d9pmQG
Gi13NG2TJ1El20qyjkI/P5xW6nQKokgark6v6B64oWOHVS5ZOgSTh1hN5phwojAa/Bma81a6QXt/
AsQltbU6RnkHqvtt6dcMAOCK2sJdgacCNFbolVO/0WEnyaweGtpB8CWsAaxaHiZmE+T1at1YYvaz
ZKtecM66GoT0d25Tk8a9hUtEyr3hxVamGcOytZzU3ZtVrRzLeRQJSIAAmwBq602sqeLD3XqCL9Zr
QhiVhBr1J5k/gR2mYBD0Si/k+KawzvvuU864fSLKznP8T4s+vL5XrpELGQ6sVVYvH8PKdtMcn2fe
A8yR2hwnJKCvYA5nzMDuN8vhvjFt28q7ijOjgJIerTCRFyxwnzlkGHBcuehp8qxXpQv/klWDCSFK
f+zBUchN9NqiJItAFyU4f3oFZ7DBuD4YJSbxt92gsyLI/JOJWYsI+I2miZDV/MIjCFeg8kvLBm+/
w4FSi1xkdht3Wptv7Us802vRQlVs8wc2WInqXoplLyHBijE7oqSxGAJXjvFV7Am7Y7UWe61oiXRU
cNiXGRAUW9nXyUt5BeiNNHTZInD5+V9vS84uYEiKwXDb72vAVlyjCtETxh0dIBIE13TOXNKIX1t9
ibhx+ddh2Q8840su3jccXHu3TOUmz0wFYOQ0Gx6xD4N5ZXIFs9s0ghy520vLqdYUnJR/Fc24jO0+
gKdQvWtKYlf/huAaf8X8D3w0HulnayNfUU6br5NUhSjvwWfyj6+T+XxgkxuNNF/ppZCq65rH0fXJ
aO3dKGnB/KnXi5lnbyV2RFZfmmuDem5e1UnUGI3qttQb9sNtG9KpEEjHPozpAvDPi/vNXFKwfp21
UQZVrqNk+HCFGHn0TP3v05biRDzX1v0jqD57IopznpV6waIYuY4VGoTbcCEeQRNtFF3S4GKyLUOz
NuNKW2R4vc6bxNDUqa2kIR+Io7Zl/BaophqBmfRXCPcKgAIyII19vL1W49J4LjGiknjyXwmT5R16
mtT+qoavTEz2qPsLC3yprVGMIuuYsnLi1VM4ASdB4cIJnU0tGdQBw2pWgfa8MRTIePp8q4GCl/O2
eBC3jOR6oRTTvZAREzWWsF9sQdVUKJZ98AO7si58dg6agvXuyFc1f+Yz9bu/UKFBA64lRcLOiKYH
BVS0koOrVKReRAuOVV04xIHKzMPov5whNpjh7yNKB5hRpxpePV/gbK0VfmU/70rKBQ+dU/WXfUVb
teO8l4KdeVnRO5rqTZcIygqdkrFpk9wPGpIStXMI0B0rZ5/fk+qdOfmw6gMbYzDROdxnTB9fZM5E
EDJXuK5Pjoct2Vlgp3hvi2ad8xF1rE/T9Gul+oLNCsfE+A3nl6efyoEn7BjXlEJDeDnfoOZC6NZ7
WpUKlHRvXtj1BBWuHSNujnvOGcRvlM6XK77oDpK1iAnBxQ4XC9CJY8v8hxwhk7VOai9QZHhkmqVI
KkeqwHoaww8oCGREN947tm70Iy3hGBfvv+kLXVEz5utXSpSYgyaumwpt7tVmx07zhHOR3zIJ37JE
yF0UhB1sb7pjKInQ5Kj3pqCitbq0lcn46kNi4YljDqBEX+M12w4gOV09qq48q31GGmRclikjDC41
XfC5x5qixkPYLZOs8HwhAWFVd32S09WUwFCO+W5eS8Ks8XBM9q73AHNAY8y1fQxC6Mu/2bpCHCEb
+NM5deCdoZp7B3FJoE8yfPXplZYMXq1yKVSw5Llv8qccDG4In2iEgHmEB3UX6KLZuSvVKP/Yn8xh
Vxv88OPzt/ylEGcM1iKU/7Jm7Q3YyYeJu8fVC7tFlb3MQGSsbyjg/ylykF+wxR1H0MWrB1mYivRy
tcAtwpQCh/tP9H/qrfeJrvd3uR9dGPGzk8QXYrN30MGjKtjJTAvGVx2qcMEgKbicjsmJyo+WBEre
E+UwltsDA04e8RmRxHBLujrfUmxlL2WkB80DizPXwkm085K99R56f0+rYrRFOnnCnhksWXy+dLXJ
FeBH29VYJ0qccy63cyXRGiEE0HkrZWT5JNBLFAx93nZKijrTuVk/JNQlZREloxkuxKLp1JX372NR
jF4zbqGsHmJQg5XrA0G8yIpFG1dd1EzxcdCI0jY5GuyTEtc0v8m2WvXG+8zNKEC5rZ7vXDxp8Q8i
Oyg4H9fkXJijGKjbvSWqhqBmoa6xeSUHpV6owzBJaub1jMYH+uSEiHEKJkS+TOddSFddWTFskA3L
EQzjYvMeVXahzIlCmKkC79fz5o58Ezn39WMgOIJuXVsDhs3RMcWfILbyRUR28ReZzQpg7IhM3hLO
d3PTaJiX4UVtBi3fhmOtIQNGbSm9+bp8dks3BjCPbBjxv7uw51HLB/QWlYAKkUdbzOUCse1GTrvw
MBoKepYn+yetD20e+kKqWwQfrzBAod/8vxuSqwD+I+ngUgOCe15FGdhRezFqf+LGPcKm4OANfzUb
yk0yix2LVwFkgsA+v+yq0y5+0zAA8p+vTfrB3Bdtv3/vxkxGGfMfUAYJstE5LRz8LFYYlAlRF57G
i2psXwz+M8f9X7lZ/hNMBMUBsj+/GfycwtPfclIr8Ok/N6ysV4oPOiyB3HXQv4A5MIu8stT6qgBX
cLPml3eoOb+7oGMiS+Gvz7RjgyVCaxccIP8Rdq4eO/icmZHbMSGm2xtHnwqzVtyUuHDW7AYtdSyK
QXwHarlFkREmXZH9rVTy9X/3tgZW6aBrx0G75BeQUpBMBO2vF1Px0FHkEtNT5cTVqvnmX0R7v7yb
1wXu26b/+y3sSVmLh9rlV8m136SFu3EfctwPNeibrNmf+Lmc5aq2oUa1xmRlqUUeZiK9y+uK6xU3
g5AR15qXFM7tmjTWn4EZ3l27aHyQFVpesjX01N+HdMqgr2a/36qaoUnqiTwddW25KFgdA9YDGyu5
8hxfChuhhGuuh13usBgy4AWu7y7ecsukKAsezhGHdxJB8/ZHfXgZlzH78myoYbDR0U5rrfdPMkjZ
wKIAw0fzLPwEG6LK/WecN5inNq3FRFNHz8JgVgPs/UL2faywczwGXaivrflBr5YOcVwjnklU6ZZN
XJB6Rekp0fhwRbXryOK7ukE2+mXDJtvfyQbLBSvx2i2HHxqZRYIeWXQi0EoYfCNeSzQzMK+BQNwh
Gt7corU8MwBULf+95dnGncPyM6xwbon7NbWqDEkpsADgFYazgYdgCeI3mWwdLwmgcNJaFWEG6cd+
7buWkFypet8G3ghRMa2bZYrLEFC7h+BdA5b56/eNXakkb+Ks9B3wqiGOXfFCKbo/uvSKQKqFeFaz
rTqu/9ZKGJXBqLeQQo8KlVF8jSONodJDbO3v7UFw7x28Tb0dg4LaNyoqTQ9GH8K89v/3NFyFiyu8
xvrIRGaX1VKTh3TfLj+TNAVI3Ynw2mkfRmc1JvQEA8DGqv34pOhQ27QgxuuX78hsVsJlKRntiqGX
NU1WLJjroShNKzB0u/1r0siG+3hTSN8WFXlXTeWbf0Lemqq7Gm6ZNhSvqss2EHepgffngmbl4yod
5Btj4e6PWU/ovgb/OIf/GWkLbESegUTJS1oDJ8NGrNQYnZHB1NE8EAzYm5WAKro7whBJ54upu9Zm
TipWQIoxugdTrD7F0qDL1aGrWmhGaAveTUQGfmjy43rNA6T732cXvbm2uSTpjgbs+pOL95+Nd6sm
cNtMUuwRg7PS9GB8BH2Xved4TvAVa3+c2FpnUZYbQwcnP9F45+4UoHu0U3Gbuw6ZvzfHrvJ6Mxi+
BIp/ITwkNVS1sdOoOn/zpXKNSALrnAjvwLr+wwKuyVE/D/XEARnztl8Z9Vv/uLVh656OBTr6F4TY
X46QkbyMFzyQ7LOMWMhYQRqJrCIdD3aNNUKy7pT5rZpMirHozJBqVVSRZP5eq4PDGDtBMRyce2/U
thOjgLufAwuBxhfQoJSLmv+APkWY2taHsFrc0oszwQZInnJRyIXYvr1HfNOZ1Y+v10VEmrbjZQs4
SB0FjGDdWKa7Ortr5dIsmWKTBbuFE2SU5qNxnGP7vM7baN6Ho7dBMmLf9omAduRBSyTanZ9zGtvS
HdCaVG7CE02LOuIews0algztndVC3vPK0csfMf+oqAEHvGcIebbzjSmQvDas7CXFtls442i26gsL
jV0hvYWIAK2EGMROC59pz34abXrFnepU/05gSuybqA6/sv7kh3oTIpzZIfaj6yBA6d6UeyANE8/X
v7xvCqlz3Sf+CuiBSUE8eTVFQfdAdF1N22RqAXdIf1CPchZun3or6gANAs9GwH/XUcwpnxMZHqmi
KBhjbZ+dBXzvwggJBCiHx2+B10vlXzpKU+pq7EJWTaj/5kkhxwYvEiHNEpSzFTM9gwwKvbI+BaEV
T2QoK9VyiMuQrJqCfI9rbN+ejqq/YEZ9mhkO1cBiFK72AW16J3Qse7TiOAdG20vlet2myDNRVgMQ
4mtAdc2o9D0CCG/QBLCrQ4qa3HNcfEzq4KmAaUL2Z8lR0yphAQNtcsu9dQPdqA27FI9IoYYth0ZH
9jFdB6CtMCyBkM5cw5nKcfVedLVk7I1hbADc7/37ymoFqkVGRuIW/BTgsU0JvjMJRePEP9LdN3LG
vVJ+P0eCzf4+gqNt4EPkxqH+szVX8si/fM63VVThS6K5SpAo1mdOzlaktlvh5MQugc2GDc/dKUVQ
RumeWjVKap+1cpw6Q0uqAXGAd49EnBsrStaqDsK4cMnG4uEUE6SDJm/CV/Lton+gpvhW3Yeq3BgY
aPeSjxcPJ1sxRcukTOkQOTUfsUGSMqPtnXRWMZQRga9Vwvnz7mWF/0IJvit2/pj8jLmsg7I4cxSE
titRVmOW+1ubwA2oJuPwNDLstJ+knJa+EgpVxaYCmgQxKApyhOFgkTbiHoEZal15i650rfiFwejX
LlZto8jcDWQ+2jbbCp26fi96F7l7Csq9BhAN/HOgJ52EedgAVUWoNJAx+znLpPIpN6TY661j0oKP
sbgI9soXRyunkYORxCfUQNloOfMUB2GdA+DruXVZwbHGZr+jiQI4gKQNcEgFsH8PjKsLoz5+FzwC
jR4OAVDYvUnSfSRHBFKV+GQ4h+7XLSXXxmS1a9TqS2aLVqqNORjLm0JGdmHUPYpDP6tca0Se9g1X
boy6RIU9a5fdjrHeM4auLVg1vRpX0BokTVaHBPfoJKfMHGo2iNQQLdQdgYyDMv2/BoPgUhwAalYX
Okd2g85FtiX0Kw4XFOuZZASzlhPUqHSuwH8RoXkFwrspx7XqLCTAjmqvAVf4nnhbrMLT1w8qUCy+
RQ0M0OyhiN8rJKMGs6md/U1wtR/g6yqmmYQRe2i8XlBMEETOIER0tYYFrm1oN5MQzOYFQhwczY8y
xrD7DbS8qEEdfob6uxV/JhMWYmzrZwoATJq/fLVDnaXtxymhsb0NU8uw8wm6sIMYxXWW1F7h/k7D
srpGjV37ZELVc0YtzJkwVVg/a21As1NMzKUpRe3l9c/ewTSAhhrB4d5Sl6n3fraGd3B3fmnzMvvo
fsdIVogw/acy9iJ4ztrDwf6SZl4rsmx4bCLT/N3xVm/P6yjyNtjEi45PS8B61g7U1+9XmZ46wKJI
MKxBEw8kzEv8w0iJrc1a8d2hjczs/GattUoO9RTtztu7oWk9e7EwIN2J3RrGPHfhvLGLZMAvJhiF
J8/k5aOngR5nu/w5Pjkp/IqnXNjCq9+bBkQAE0P1BCjaM46BmO9vMAyf0YcOz3Nmm5pkSKB93lvq
Lj9BUuTHVowCqM17af/Uy4bxKsGare/0f5UdlA3wyYkzCDG4gIisGBfcE2pHvleOSbiRQI7l4rPA
+2IG6O8WJZL8l6P6raU5IlU5uPvl7HhV7Ud20fVWvx6bjUb0eZOWJCdkgSdLoDFUFX9rENDy7djs
xwcBK9pug3GcWBn8hFWcTsSaJmZG0z2rGU7VMxZMvEpaWbMzE9RIB+vyVPZa/Ga2VBuBwa3/nMDM
ZvJF0R0kVqmIX2IbVpSg2BJ6/r8aIAj9Wtt9FSk2qz+Ud0EgFo/pnmGKHLlNbusttEnSKJFuoHXM
EglI/GxuohWGea7afNCTTahKqy5ZrlluqCuFcm0I1BJR0VEzIvuUB6qLQ5NLVqu+QPKlxch+7m1i
a2RPvMgrS5v9M5NbeZhg/Q6y9pVQIQ6zqHwGc6cOu0GSOEtvAFASku7e26/jCCBd6XwX7ZHNwCfm
Y7rJwvll9csVisj4CJYAXi4dexL0xHk1pF7fLnPDWts8gGACkmVY1AXIvu/BXQ3Co/iIbNHyLQBc
n/2vupCJVq7M3vIHjXO/xGX8NQIMo5LbnKQl48ZMLPDVCCZQWRejXZqcEI4qGZWbaNvZKyte3TsD
nGtF2tjPMaheTGCOswT01ViQ9QeekR4jYHyc/UwcMhHuT9FW/0REPxTCXRI1HdIEg5ve+aoYehPF
g9TL01kydOoGokwqI0ilFFnaNoPqa4G/77p2nZ9ptGn7YrbHZumczmEP/5dFKIJThRfy/0SzFeds
XC7CBDrhumQZ0Mb+Sdhdmx+hWXSIU6DnLBpy3EqODgHR4a5ooYNGKf2Tx0XIv6EFWPo2WQaMQHuE
dcxDcSMjTSPoySxsEGiEUaXsTV1mF5doYRvZzR8IM3ESpqpPJfOwzvKYlUqTAueSWHbzesQEx4rI
cPn2up8cW3rKoRsGJ3c2eXrZeJAAzokWL8B2d5FpwJadCftHn7GV1OdE6kwTnozbRrO0kvWRUy0i
vBV05v8fRlqcMm/iAf3Qfyi8TkdTmYyyaelNGS7jUDQrR2zuRJCapUZR9JA0mo5nlBldvNGekbHP
hpkY1J35Hswj3UItoy4bJTTIIFMgprig0OZPmag2wAMeu8MZq02KqUHx5hOk5jrkiz51OCx9NhcV
HBvM/or7XBO2rwzUZ4lmtJP3UThoKuJIJOBiquI0GtF7cXtAYiiC0YHMSrSy0UzJOz8QkTINJW3O
i3b7nm9ir6SlFobSS/vEEQjWCzSA6BNyZ0+qyOgiBhL0FGhqf8PAal9Xm62pvnJ2ZWisffBN2zwO
k1OyodOYViDCEsb+HPhVI0noJsxPhEliSpCT8wN8DWDowHdIxAwJGpX+zUauU60NCTjElV0F1LxN
rf156vU1pQ9Ca28uGxRJ45lHi/zBSJC5/2ANvPx4C2qdSe4mJkdBM8c/HHL7Zs5UweCktyAVXslQ
pdYywox5BcNYzoioKGfnzfwvt1DJiZWGZl3UqIScPr6qdA/TFWnOueJvgPca6G4YfzWyTF0sfT6m
FmTM1icIgPvq92Fto0imV03Mu2EpFelEgEM/12JkGBLe1ZBsOhAN/ydlXKIIsW3jz5vQCotRK0Rr
79s8HbQdrry7Tm57J+m9EZVxAuLqi9PcjL6ah+tWiHP4qbhAdRznh89tlN2mp9aeeN/AR+lUM/b/
kasfy9nmu7FNpOySuCzZOgoWKa8pkBjyIaQ3GS+C+kUT/rpIHhvkaSSdIIoxs39VlhJ/SaHvIsbh
pDs/A2UcHcbzWuKpOZ8nCkzCoD3a/TBderk2BCguo9X/Jr69FXIIk7czzo59C8eleTmK37M6bs5F
1R+BLjf8iS/A5tt55uV6i3PrMIEZC3xBEImFsds8lVIUP+uWGAey/+Su6U176MhkSkYMJCQpuVmW
BAaMJ0FXkqrLG16sFtSb9zgoUlMe01y9h7xN5sU5ZDnaUL3jcrvumZHz74pUt2rxwLVDLUZBqzoE
vr7SygiYANNG6WOqosuJGtP8PtPcMujCNCpReyD97DLkG4VCm29iC06qcgHyhhCULCW9fwK72cfM
SOCqonEnH15eRZNXMMpDRSvHNYwbgGmeKLgbhwubWPhlMl61RIvv1Xa3erF7ub9idrEnsDJjDK98
PCk03JlnqvfYTLQotoqYydRFhx1lwssZ+uycaBQOgy12QiJqrfGRzovqtx2lG4ozu0v7yjVPNEUa
GvoE6uxSKkRdzV577yi8hnC3mPFotWOMA7GtUCKh6k77AXC9IoGyi/Lr6lzDtlxe9n4pQm7CqAqQ
zUC7OqHjrR62XP8xeeRee4Uk6ootdRvvAYZ5SPuDKll9vSlzJTEKDtIcJqqSFtepwM81cpBBhBZb
yIvgQQmaTXXKG1OZ4HowduSW5ljjk2xueVCfc/PWTH6QRPiWsuF8mkBx1Buy2ebnwljCiVUzoSKM
YoFO6P1gDlq2PI3UYodre19AIHI7WXL2JeR6niqsjgHvEdc0f46xq08P7HDkCAmGpAOuP+QEWkjc
tPunOi0QU4Wd6RRYJ6Fq6/QWM0kM9eheJf+wgj6jshStwhG1BXoeLrQ7t4rpZNq+t/MffAAktIKd
eTLR+Mk42YiImuyGPnTs/uPolBKnTP0f1ieTRBwNkIjEQgwiaHsoi8xwhDVsqZ2sHf2j1qgE8HMb
1jmoD6EBk6/+1Az0Kp+ArlzvOfgRRv9nlVdeCQ1udQC30RQ3Ihr88Qtgiq5eiKIpp5FgQaCkl6+R
wG2q79uAiK11kuHklDKo+y37Ib9VTuMdQmES7ly0Lb7uba9xPy5+RCc9V0kCmkt6xReXnZL9f6mO
tDnlxVdYocWhBjx+z+Fn3gpctyO6s+Wf7QFCCOY/1S5pz1qhwWdKNE1d8xSAJopp25wjNt+UDJAX
Ey+0w2+HcFDWDm2sGJ6X/V69UyQH+2+yRlYxWECiQnfBhVOxb9p0UU2gDxsH11aJ7LTJY2Jn9xFL
qIzhKdgffFGpEPJxsZGakrKtYg0aKxjitUHbJP5ZEgMWthhPAPhvnekFMFvCUVPzT0r6sgPfZM1e
qqIi8gNyJd4KzpajzAryoi7quaXKwmp6eysjmz3xbtIC3GGsAu3GuLDFdOu5c2TuYAXTCqgv9Zzo
C68HrksiTjYD8ICnFxurQoKqsot3nq2OCT/bO19Lhk0KCTwBuoFFrdOYZc5BU8G9ZWdfvDTgFSIF
UOmFxalCVovIMc3BQvkat7sEnR0Mr5PE77TNGb9FF+SlZ2ZwawqIFKVt1HJlkiMtK7sSSoL+CI+0
fb0nEgnU2IcnTWo5wX5LQkHMMtjcmGqpzV9V8gAfVLQLgzl8lNjbucA/qWbo+N46NrkLDAvLh8hF
oPyVpzuXge8Ub1zyQ+QL9Jt1ZTVZVSXGznLKvuKlLuqguwbGI5mcR+JcwBzQJHEtpECTQR248IVZ
2UdQ6y+jo0iUFKOZ4OYcbjkSOpGI2SKLt/Kgg65KD5lRyElO/EJ3Vfd5NYM2lxf4WUhNwWXBYRsb
stVty2GyXTN8UWQJ64WG170pNJ9Lq/XF5bo3rrvNDCQTM7n6uYT6ffqLX97weFxTVqvYogEZwVZQ
PbBTVIfZnkVVO8A44neoz/Ec9pBIvxeiLai+Q9yIT2+kHj+K7qvPLLB31dZiKybWNOonCI0MsGaV
NV+PGMBPJRqcNoaSLeTWk4ptzQ3FHzEZ+4udIGu6j0QA2v9AjJUOGY0E3OWM+V0T3ewpqyO4I+nb
CiyWIx9HmBDQ/lbnpBPV/w7udcB/0c/aW2eM5nwV3rk4H10nUcqwYVML4++2/d093K2/iOUauStk
YzG88I/sGWnGe8NwpMswXKsXUIsVF5v6k7GtC8oBA3DRn8BeLKACIjmCWCfrGasJvXKoS3K+DRKl
fgABQ5ubOrbwaQc6DKfsjo5Yr/o1ws2So11omo87HTmttUivUFrsyH6NrV79iF6Ut9OOSmBaRanP
sir7vSobKb7SeQQSJFIOlt9aoWatZzIPle+L7C0zU6HbjZeeYBHTc4in/HlbJxubtKXaiDRumxC4
zm2C4Al9FTv3Ft/lN8PjJ/CDsblvW93k58YBu9V1+XbrZmTM1kR0QQCx/RUsqONoQ/ktZVKQDRvq
BppOdSjQzUQOlLisgIPlDOyn9ywLU3D8nn/4YpHYvFHeeFvrfNtQYSgJOpzcm4IjaBaHsAQ5RWt/
DtdxLKWhnNkTTCidEPHIJ04VKaFKOLeCGqFeh74VokBqUVyFmXGXfzkfVK+sdosckQCsXyXMyd9N
Pcw0MdIiHePnth9ZR4pP9fyQlZO5ETmo9xYvfQuktdfmDSNFF4OLMOBlA83mUwCUkE3RkM0sYhd3
pOrrDCBhIbfdhVWNXt7LpUnD0s75X2rd04stPCLyxZ0GpHgCZuF+bpU0tVRAIekNftpdSCLvq944
wzv9FI2+TxeOaHRWt54UJsFH82jYLdV1N6ECQP8i1JsIJZmdBo13nWLKFIi5R6pw2r+mWdrm6/ay
F8xjHsyFpvoWoYZ5x3Wl0LLsjFoFytiinsSPVZMpg3hrJUTyAOiXL5tzxbHQaf53x3oGxDR3pbxf
7gIT2De/ZQ786j90v7tljw49TyFRpAA8UmL/dgVPE57+JjcfP7zQVph+xmRzUiMUalzSKlmc+7g5
9BPTSF4RYbvtYSfb+9jcj0+SxQvHuTA0f523zq7mIF56YWpHqPSs0OE9PhV7bSzLjDmglgVX8ngE
TAl2zZX07VD4Acb1lNcQsWU9sBtHv/8W8YI4+2OIICzNhckLMmlSa1ND9NXQa4x49fX6+llw/syd
CJOMh6nUgmtbDQveUMqu5taOYDSqM3GEbj0z0/YLLqrydsT9XOVtA7MU4eJkCMJlS9PRh0+EFvcm
HtRuWDvKhRmfv93anM6RdnC+/0Tg33Oh3ScfmtLCXFw+euDUhrivDGfou+AUBR3d0u45oyw8Me1b
se+AJe82Z7+XVAPpdOHFmlHZ1RvxdPI4ZcFx42Ks/Utaci86Bg9UHXFn1cEb71ow0nqiXoB0tjSd
HEe0eYhGsf/dLcElm2/NXzT5TyFVA0PV0aASBA2R9FajFfBRjprogjugfDeF0MI980yFZL2Dd8AW
geow5E3Fk7NRhCkWNd31BTUAi2ARHE0DK7qNRaJE/QBaYsMCnxLvz6X8WXjG2XB6nbhoXc88JlOG
lgvFL2p4Brip03FKDPOMAR82pIw24fLhoxVVnfbFUkTibeosBxGAFVeC1NuCanvtS2N2i7JZUwj/
MGWSfnaaD0WYFaWnR9YIJ8TL/OCUD4IlXxszvLSNZ3mM2WRtRY25JxFE+fF2EgR8GoYJcLIe0knt
JpcY0mQ4TV+Tn26mU/KH1qvOdjF+smKvEvhdv64XMyohTHpr7GiKVN6tMsAQOEcOU/JnUaYeoBMu
Uo8bCVpHth9qn5W11xUu7UNiRko7ry+DivtR2sGb6FBt+ppkB4R/3Dwb0rsmk7T881xxzgun68JJ
jDzv8Y9FrL0e9ITEjgoK8+33BRtvhNeOxUBZy+G1fmWh84xOLtxxJ5Ldvq/KXwlG90HniTxGB+0t
A+SXoxbe+onDqnEx2cP7Enf+jf3HNBRmKZgzbc49XDq3nfFHRj5ZWMwR9J7bZ79P6L7aIGR5XtNu
MUrSzmVJgFE9EI1UQCawtraX2764XGX+XDHxkETo966JRgQAae6fRyQJJYAf1NKl7jPqT472/y+3
QQv4t5imyghuKHoNWnp8Vijz7Zw6yPwkIuYPYDili7NnJj4su1wySpdhTHahJUXcL8Mp9kIqH6x3
f+IuAUra3Dzm+bcfN/OqIHdSj8ebZnSyUlLu/jaRQQDlF5Rviwi5HiYM2j+PpYQgUyRCIMhvPj5d
siI4LCD4xyW2ttoATojwGWOjwukCTcZRZatzdI4eIVk0zSIcP+IMGsWvvJuLjxc8+70R94WAbCm3
l20cgB+zSaQwP6qFgiXJrbSsPem7VGtn6AO7N5KPsifblJhPQfkODUXz/ZDbcy5/sGbOuh10HsBC
bPwzyhH3j1AYRMq7I3aMP3XB3Xrykv21aaSHJIOq67apb7kUXLsNH9gZ+qJti5+HG142rqxFXSoc
HrQCSykYauooSeRj8Ri/cM9z2eFTZNctpsPZHqimlati5WfPaSU05RyCDG1ucGjITOMcBvxTh5/w
TWy9QnlyC1nNuSEFeHSpq8kB4g1fIhKWyZK6hiY41aloP6blVV7JXLxJKL4iFDi8bioC1SRFxBoE
bg2XGGCV9bW7Mx8CaHkMzqZXwhmNg8Dn4zH2bH5pza+CpHbyUCSxztLO+QgTWmkeJTGwF1CKiGwp
SdbdV2BZEhUGaABRrRna5nNpbrMSgB72DfYnIjJ8Xw9mhbn+gTEeS3mqLXzEP4Ox128FNR9/JlqO
ZMqLrC259tSh8vbtmQ9FiSrn/DhwdNuYZF1x1/XC9pEtXUqWFMdWLpGxh5kXvWtYHgj0HmQsAg5Z
VOaogSnzQZ8aAIdG6ZzFWMAmWERsWm/thL/2gywGZqE5xDmEXzj11iRUVPy1vB/IymjRD8mrX497
lfbDyTfiEttcuF1LJ1kpXUmD9Nx9W+RGk7QzSD6gZimbH4qEt0XwFnwlf6TOveVdbFXJrWptDmK9
WVGtf6R+NfQJ7wdg/Rd3cd1TXRX2RZ7YQ5hiARGNieLXlxhMM4kcXb1dPr3hFsStCoptpNPlLvOa
wQDVxk6ru9TNMbKRYdpP10spLotTGG+HxAfSNxHbjSDPev7O9DMipJGq14YCmvZOy4sVdonC9stH
b8l1wgjMTVE3exiLn0Z1mceHKKvTrm4j2dkPwh+KfZlbJ7Hb3i+8kiGFBamaAb8ifzhHBDX7lOH/
VVLX7zS84H1Z4230gPmEQynJHX/Hm5KuOQ1LPhwsdUfcfW3tDIh9uzA6b+za9wfiW/RgzEKW6aVI
zv88mevLy8ESifm3dthPwsmPmIRe0MKw4mVEmQNA+QomHKhQuA0lrq4CtpDn9/wOnlByE+C09RHr
GTjW0VfW62Pu+m3qf1YSYkCb4dYnN0eTdnqixBBU5mOPbCfYQnz+KpJQjhuhyDiUXy2MeGGL4o0u
/w8bL8s71XFUG/BmgyUHeERPx21IoSoSFLgwthNLynBbHY4GfxU+21j0TYnAqRCMBJ/toO/dED+x
aLoJZl0ITDclGrP+TsQg8YuiCewmKqhE+q6/0Rzn4evxshLlla+2mivuBi5Qy+2Hf2QWrn1De6j8
R6UuLXnkKPrDKlGgYWfGK2KU0bKQWQGgSywXhUsKvateGJRBpmXHWB1eOkfdu3YP8cA6d35PCHcO
V0bCikpTTwyFGZP2ynhYd6mirpomBwiW0qW+nT8a1VG+0AWc6M+XkAruBTf0phrchSGBnzYOO1z3
IvgBb+sEL5K4ve79d+JUJEvktLmS/1Kqhn56yjT0D+1JOgZDrrAiC0GERwcwkPvSm4AT5XFSooOQ
ciBV5SgltR+0pyLQsfskqqZy1Mp5d75p4HWyiTFr0LKHosgCPu4u91C199+6ko2Vw4qHGmd3qMQq
uwVIP3d09pRYLwZ0wBXTo/zrwWbYkMh4EmQSwu3hXJqT5YNelvmrLn7QZQyNNQzemPQGGieMpwTN
lL+25RuRfJACBWAi6PIMTecmJzgyTwc7RL5vK9UFLd73jE4+HCDTGXht4tUayOX6kUzQ8zrXp3kT
H6KZ8neIDJ+J8LwnPf3V11HdfLusEBF6WHbLPqYItfc9qB4h2DOhLGGWu0lR594bQf0C2fL3KU5U
6CBYdUMnUTFkwE4o9jZzUD6gSThtNHVS0Es99NEt7mWk9QDThCcRwCessbwUy7d54/i55WNHpXUv
/LSpi+dblaZjY5GphXq4ahQkQ6rHVLsAL9gTpoy0NKCC+tApu3T3sWiT7mqPtX2tLvJ1F0Jdu/Bl
aNMj8/rJgFJ1b9Q1pan0XRWh7jazwwJhUHCr196q4xKKUyjFjBEp3Royiuoi1Vcogk3PZ05R7Jr9
x0NQajhi8jsxn/Z2/SYN3UArnNcxmoHiGlceT+3g3gaiIA0rAAQjTES/M6oh80DMLsFf6tJLX+nh
rup0kK1TL+45S9fJx/e+ms6/4HATR0+4fCpGX5P3ZxREujnpJr3YFI9SUIeuIuK0PTESjGvucyNA
9PRG+Bx7+qLjuwte/riu4orkh5eIUqCqJcxxPE0Zd/hn1RzlpSK5mi2dj7m7yU3BDaGIxFUi/j3p
sw3rRGN64WLOPUITqlclsK7ozKtkqKMdEQ49UdnmM7hOudlatfoC/qgRjqRsMc+d82m2wbhYq4bz
roF2xtIYGu9DJtka9ITBGIvlNK+nx+roSYzZkedtMkTi60UIO3JZ5j53viEFWCx2fLIz6Vuwevqb
SuRDV2X0RHV/m0XdN3tyGuS3tkqnbrVUdwAs8GssdqdoAXOQS2N8aHXPdiOs2JoUSJr0mRapNmf6
rauPC1LrU7LgtrSOCHBs8m3b5dTV78Mhz/5mvqXGGWqOXmzEfFDDDqOk2gmSWP/1IRrMKOrtbJ+L
AJcFGyYZgUj1erVyVsu0vOuX0AyasB8T4YYXfanzLKiy+rd8ZB08fl9o9WItKanW1Qwesv/2lAR8
MjjCJDwg2dpppqT2msjDvmydiIbZSRvZmuE6m6oTVNXuo6JstYXucs+wrKv3STWy31zOLJTB54dX
w4gP6TN8AfO6pDREJOOwjFNYxNhgoRMSz+FzwQPPZp/iDC25fUKK0ivGgMtp7V9gyjJXU0t1TlV7
igugtl0OLG+6VvEluRcAm7hQaxedB7788ByU1HQuDvWYo5QkSdjS6H6UVQgSYAPjkyQV44h50P2P
cBYkJ5mS1rBjviOrh1gjwGOEmh06DtscfS2P5kt5lTTTLeubY8WXZE87eKG2qyVJTg5FjprDGNcK
Dpvx9ApBGSh1NvlWEeGz8b3s3nXcYJYaasXvFNbsJiWXtiR7FOrw5OCyYPOEfW/NyR9SYfLPxJvz
u2A1EPVj+F09YRxbOhtnsnjDGIqfKy/OytEbzfqQEJrFiTmDi9kthtSbF1PEXpDnYXIQfDA68Ymu
lOvAnzWxKVaz6C2JwwFOajXS1xCQFmhTiqq8IgAIOQUszgwD85i9HboLYMR7wQoDVUFplh33Nxwk
ico0S6vGZzVrnAq5RUgNC5a3TX4En22lzIlZ6tx5KrG7XeRdVPocVprLmk/tT0XJHuYkM/B9m7cP
nVqoIrB9vR7PIZNx/hH1OgOxGqdzku+yPOzwncpcVy1orgyEExML8T/wFbACW85eB/JlK8bEEMj7
zb/+/ilAvrotnsZ02avE6wt1gZDNSpPUprf/c8cqouHutlbl5qCBLqOJGy3wmhpDRMBfTHxYqQZ2
FMJmzPsV8LCJCx+PAZv36tiYAR85A71n6OhPGKse3rOexwfyvnSym4rSa4PTrq8isyE20TQNjmt+
pP4BznzDyfE5AmMq9it31qxQ5Mk283zY8qVMecgi/AQeYMTcuS3dJCx+R2X29wn6gXd7RIc25ZR1
YeYcTCr6JuQgjrDSjDSb9NKUu2xig/gIpSRoAULNKzG+tQcTYcPRj0ZEHhAgWKRSMsWQGeDra/kg
BoU+HuqlmpqsFQlB2GYXcTMUHjLFQ0eFy+ITrEbvT5Kaur/mby3Hhmi/pL4GIkdK+ZxiF/tsU8RF
piAJbzehxcaTb5Vbo2pDQsWpxMFMvlbu+ECeWnqG2rh26fwyzAXyEHF7dZ6wgvwIE8n6bVjKsBmK
cbrJSpKNFhYo27VhdyGbLz9CUdfOihysWOLqVMPoHMZcIL8FcDRhxQz2ONq0uqjzYdUFNISt/2km
k/QvgbLe3KMf8yTNpqWHYjr7MDcjGe5CU+QzZLS5kAJXNEdOp4VXdUhbBPXTLLGfbLn/FHh5iS9j
EPGtfVIvzI/YyClOxLVHSTv+pjbPftVKz55PeyK4iuVU4C0WbefbNwdP4E14rxeQdQEpIfRQ71q0
3h5qVCINe97E74xQSGRoDGlEceurQZjLyyTnMkQ9DmaUHJBFY2HZ7aOEYI1vcUapqodwa1SY5JjN
LMocCvg5AmYFHpi2zrHKD7rUYqHmNgsboB0FVAo/cnXZ9PlIOz13Tmc1drdo+OUfTwpRJPwWf2yN
s/AifLWxz8QFH/9HwZTk+cyWbGGaJLwoR/IrjEqzCO8c3mkdmB58bLdbBnrX1l9EqvggrmR4acFk
yt4/MUhuGOxWTQkSNO7rIscYwEySfke2r5Tky2TPWct6YQ4tojuUXvLCzFmd+gHdVYn73zMN++Tj
aDD+xxDKkUR8rC0oXPE12v9FU8OVq40+YjQyllq+8iUhDUuVi/hheF35/0zwaqJZaXvBrrDAMgJN
Yjax2j30gty57NOrnY1+KQY6y5pNgxcUFNhaanZXHOhEuRJUq0Gqq/7JyGLFrAoMFpduXbRWxATw
y5Q78qm+Gro/FhKd4+L4PVimpwOFY24quIdpdPd+m/Y2fT3DE8v10ZAPiMPBjgetni/Ve3eqQ+3m
cHkld5RMCD+eS+WMosvScNE8CFLW2lB6cU2IMVWpP2vo6ouWf0OnVtCAR9nC3CoVxdzMOn5VrpPU
xlnA1piHTvER8/5UPLG4+vwDc2dyLEPIPmtkfesS6jfRUm9C3sIEOdWYkWQD56fIarpsAGzNlBPW
pdsndKIXCYuOCslj23F/Cy1x0xHrFOAtFmp7T+cOat/dRwFGpNE42cjbjLDyc542dhG/vA/3y9qE
cSYrV7iflvoQbFeKg63hnenpa7UPG0DsO3DjmoIdd3Lfajt+J1r9fWcgNzO8cOZtTKR7peHZoKcc
XFKktofhbqKGtkkiilQ7jLsF8kxH9vI1R3ykTYzf5ss0GuUMorjnBUz7hNJ+jYec7klqvFArostC
Jt+ypsx0ZjyyKTgyu94btvOn6G9DCbh22qPjpmZ4/XMosu1NqI9R900d/1xH1+N/sGaWY6Xlscrt
AX+tM/MMFZJhOTbNngiAU/Ll70otwndupT++EEeeol0Vk1V4WH7UAAvarrgP5UZtPKP654H2C8Is
A17VcI06TGmY1P3Lny+Mor7an2Lvs2psLBIm71iNQMybdLlU2tBabiknI47TcFWlpwC3TJpfdN2D
AzPHc7FSKI8qhRGRFcWBQvHbnIFDxv5gZ4F2BZAdSp4WdrTWudOJWvRsZB+4U7RFQHWUPWqhbeZz
s7XkfO98M5vqmryuDFekjdneMHbjUdBfLcpHOV9550Tt/G7IWNjMev3VWEw6xa2pRKmvtcfpLYu+
k56Mw9+n5sgYwyzl4e3P2HgXsKiCyKDYMQCvJDJPwBoogaMY8s59XPBvku11zyGf2GexpEYVqZS4
0Y9GC9KoX4k3Y4vqOqUAteF7nddbXZUVx8WUhM6TmQVLgXFGbEOIzG4uNO5YZ24XsjBsh3NjuD9u
P9TpL5rSmdiy4YGuPKAaHsC6z7MgX1f69H/mVW/msgqrZW7JtfyUUJYEF8JqlrEnFcMZbpEeH+xF
WcmA01Hn8Ox/aMGojJWkL2Q+2SIL3BsimETor0oMLnkT9c1C7LzzBYLwVJUpB/93ttPoMrYVA8wy
ZiAEjuqf9dSrjGeYkPq5ZCYMcbEwj/7ukgrZsXDVeCBsYKx1KYLhBCPyO7s8p4FQDzYOcXIX+MGu
JS3MFd+n5gJdvnRc9SU9VyCvn0Yk3Q6mGBKefJgpH5vsyPgIwzax3T/m1dSwlW3U9X18kPO/27/T
3N5Ds0pPQkowyv/v6H0h7OfxNVgFltcUH7lw0aH9Dh1eXzxrvH0yNceVYB8LpEMiAcB/zkRXqGOA
bXQKNlgW6L3W6jDwJGJViHy8jgQLdpLOrCw8r7xxoJraxKJr74ilv4AKSkkmh9MTe9hlH7vZa+W9
C0jUnGLTequFAKGKcItKRVqfLaq0szZbeq7VaaXNQ4wA18TxZKmf9afCxzIpdWFapEUpHVnJKGKc
dL0vKP+V9Rx2k1rgVgaigHbUulOVr9xHuF2/lGzHdXxmO1DNL8R7D4XKF/5zVKJQwX87muF+BY0/
9MBm7I45Jl/BK6+zi8+hDxBOQ4Uthr1v7lNNfyWFYQkfvbBI0nQ2uHRrht3L6ZdV1ICnY6qmk2d3
DJ1GBQ/0w9pazaAJOg1qzev4VN7/fd20eGLbIIxu6bht5iEqEuFudHFJoVcFqQvY5yE9KsArSTxq
S7iRd3NiVeuyfH9YdaOjiAvHfewxeDMS4rs7v/BLKqrJ5+jL6uLvN3uG/7uCYsPWtgvTtZ2TWIb0
p5JYQW9HbgjHvc1NS3hljAN8X9Hw2kOVT+7zJP1JK5uZTrlngtdqrvBA2v2hIDu9WOQCSA3qRfZb
cPrOrXX2tlSzvRPKoDL5eCkieQzqSd5NOlS35Bn6/qCDkMqlA5q0SHIn5XZ9Ie91kLK9nAKp8J/W
dRXqKoL5xt4iNES2SqScDf76Tju0zDf/HlyleS3HIyZy0RO03Bw3aVX5Tis0py69bbtvIe/8HlFU
sr/i169qDZTKA5s0zHPUnB9t84r9ysVsOhAVTS5R0p5xJoIvRWmccIPzCOg0utuq7GZLxzFR//f1
bG3XA+07cKR/oXGwvgle+ALYbAUAbish6KUjj315k2FK3AvgryoqNDQ0JNRonCHK5FJyWdqhsdzs
nDQ/oUnIM4Cikz6cB46jhUP2pyoCNLDP2P97bfPYaHp3lSX2T8tvnkJSICJ/TD0Y/RZpwInD1Aq7
CRVRCoAw81VubyrLEIWielZJRw0Dl/SOQybjKggAbaX3x7A5F/OraJGqYghu+3v1j0Y26wiYRS/s
YzvvT6rlZgR8r8aM0QJAoymeLtMUyopy1/LBEvtOmtRlT5TyU7UpsmR22Ryc1MFDKSJN0O784UTh
sGzurwYZQd8CXqTiHKEGWRHMOxPI0N1QWAT7PF4C7VWqfFg+vjP5AzPug6CoK4fFzC0kqfGwnl6s
8UAhhILus/6xoRVL3X0Ocp2Rk6qM2iX32ro2IdkL6qFMDROAM3dbPIHxPSHWn9Exrz/SNxQlmP6T
UOhdJPOgr3zqNr0A7tB9XwutckYrTMZhqUh0XvQfivxK4Nl3gQpXXX5QcwXhQ06b+t01G2nRi9C9
qovLT8Ux3SaP4lMs1d5GUl/m9sjHgCnGBpW6oA9xgmRrALeAYDYahG8VtzCq2b8w+zSs2vXPJeal
AscOTxhU/ZLk5arKgDe5TM1ani3S0ebAeRAHvljDtLHCq599dXZhwZofI6ODePIs4ovw8LgPycqK
IpJpy6FbwjbWmrFAlCTksrxlNXWmO8X53dxwmDDBCn7PSl8sD4xq5VLDaUVfkl5gBvpfFk9AW7YT
lUX3HIY4grTN3tixJpfFcLVGmtVqZS3ckAsPEqBP9Aj6Q17lUQCoOiIg2feJHqQN0yC98IV7yhhi
FA6WWZ8xKcFHTGrQ0g78Vt0mdNJSd8aOZGZaHBlpwB/6o516CAmWfoFC39GbRQvLmGajK+k8FZWg
24fJ9/PKMiekkJD9g6icTqQawXAyeUSGhUeW93pPq8P8+jLcknKf996HFeTs/J7uPD3cIX6rKCS+
ApmClE4cRT2U21G6XEXNMdRmmxc3LBMLTZgmeNybe0NUw6NXEPxYmb/Xooyyf2dTNxIDAbza6+u3
2QB+1MkXCs7aqZmUx0j5dUnufYwaW3hUFdt0xGEJySTViyowfXLf8BcrXfbZGLuGKTKv7W/jjPqu
jvN6cACCgzZIyRGD1+Hrj3VGfpJ60WUaYselNLuPEVxmPoyNpEYet2wxMVsgXcURGOLYfG9UVlNH
Hmq9g0+kblWxpW5DVo47HgJD/1Wh085dWczUeLVbJoUTrDJ2VFhQos6hceIf8xZYf6hOuQgCyC0P
7pA2fMCsmQktoiMZDNR/GCtVVexSxC3lmNcJYfT+UPmUMJo+lBeJXBwlFv81uSZ4PnV8ZHziKilu
PctdUrGU8LGTjgYY+l1a5qrIH6+P1LYn3FGNXnlZ6yINm3R9UR2rUthq1C13REzPKnh1ujjVxWcb
+IVEc97+gkL9k10x4OpAad12TpE234VdtEya5QTGRe6qOgt9+xO52KgcQ0tdC72wKvsIMGjn5kOZ
+i2ZFVhdATY/vZkgyUjPUe1iZ0xh3gZ/UTWvBe67O4D99z/ogyzFAjAMl1CeA4AjxNUB9RRQBNa1
rAy276rWu0FvO7iX4MjUhNfE1rncrxRAMNE86so+xRrMs8h+Ed72TejpU9l/EpyLSPwYxlcij1hE
AfVRReM3LIY3oxzW0haSroVpoI6RXRCZPsUecX8SC58W52WXWgaIaDkipO/QAHln988CXJDEIRzv
u1O5nyIEv62h/cELcyoRCODoyGoW4EMatk/ojyRHrETlDbwM67u2mbAI5oW8ZXhZhe2pSqFr3MQ2
xiMYcAHD8CXID3iQswUcKILohSxuYmFj8GwXVVRY1OwJHpcpSdSg000hmGNX9a4eTjONzVbaWoRc
jR2iet905V9aaHzCmM2AJGKBXHEzK3UfVqmTto8w/Rl0R4LGzdDCPBGPdzJKpV8hU1LvhLsIIbOv
jFpM5E212Bnod5BXH4LFIetr+oZPCbIi0N7++a2Q6EYd9q0uxVe5lUUpWeZKDUO8Hku4W9/3nWtt
IL/c4MIed3ogan95NR7VHWYkgDuDprXfnnLy1PiMUAMO0cFOQyJv3fdODnCSSW3PPem3kNP9KF+W
ZKQQ4encMfRQQ69jjo+7TNwnaZY+D0E/iW+S9nuLel9k2r3gBDQeoDSOUzwjSRzgM+A/xcy6L7cJ
IYm32B+r6kTAacI6Lp6WN/vI1UrsKHcgUQeR1m3GDT/gACzQDYqk/ofCyrt5KRSHD6pYSJ1og/ef
7i78O6cJWaRW5xD7IHMEmsA33l45PNO/ddjYVX6R6aalTKvwltTrR+2Lz1V12/K2SX5zNlYk4IkT
PaqMMlGZViqe1baAhQnwCabR7yaOe6MuyaMOmGw+vRbOu1eMwWhsx8iheWCCUIsg3g96wkRCuD+f
wXNfiW+QP2V5fT3/xzGUt9TLCQEmysN4C8TBeq7pvoSPYarGjjj+mbkOT/xlzUjLH2R+JYQlFpQU
AyxYVu3JP/XHLHVwjIOPJmHk91MIkE2jBOYFSWHNFVMMVLzGT4lXu77pG7kwFhiM6Kya4dcFCvI+
mQDfbd0CrdJu0STIkfn1gT/7esM08dBPqQGoEuGOjroniOg2WMWgwEkhjliQH1scGcX23zaNxD1w
FQwWcKQQcx1GHaMTgA3JuilZlQIf3dCOw0uovu9nqTveNqlRYm4Rzhf3qLVgzBBm5f0KxWi14OKQ
I7xXloIw7a8RxVBH3MC5KewXlXq0WGtwJoutYVYjMcJMHxoHIWYoRWLDfD0WMdRrHHj9wrJ8svxu
zMGNn36Rpy0P8SnNbz10RFs6idiNthUn7sUhw0I2q1hBANolDWW9XLPD1tySQGobxbr2+woch2fb
aKRf4f8D1O7g19yWCSTLCoNqtKS5yfpxYweV8V6jfB+7WDlPLXM5sLvxGk3gB19aN0J3Qe7vHY5v
39lpDU9xW7sEL85SGVCrsov0UmrrcVPh0roaMvX8bvF9HMWGHtfZSbbG0CB3o25Gg2fbU6b8136e
xus8A1k5KE5Ea/j/gdlKKFiQsHihH7xg+a1rtekA1iPuXx/pW3wHVpR+MtkDrQU6D3EpZ1uCfIA2
bmbUmYn29XbTUO6Qgo4IQI5trLo1gLZFYJQiuNbmaFKCAHDJJ4eQKV+rkQDjLS4njvkl5rboLA5/
Q6KVnf9OiPjSNXHv0fJanPQcL/ige2hQfRFQqgOE1E42E8EwiiObWapCJEct2Dpp+NTT3dVFQ3RQ
jjG6UtryDkBHO71Tmw6UVpdYn9wbYdTsxZCQDqtAUnHtlVxEr+kGWo9ZWr41iamTwrlcD5fFhYpC
XeI6jD3LmsV/mFptOFqkuKomlcb7sXXP+f34JackCOiEwGIIeEAbXxTeSlYz6MhZSjrYG+jf/B6c
NgJotQSHG5RRvVqDUJfCe1mSe2s/UcuyZfURPuSK1bSCKhTK8xLp+0SU03BolxGYSKXj5jldDyaf
37wloIA73HUnwnkxcmQhizeqGrTvej0w0kwz+Mi7bVsiCZg4j/zlxMUvjG4jEsJaTpg6doPPESD9
IlvettawU9tKwOXbJS3cVNkaepnqxUU8I+bfKooPudn5ATvkOvhhHSivHBWj0DzJh/3eOcBMLG9P
vPbnIUIYs8vzA5I6NE9Hrd5NC0RW2frCaZw6b+1lcNuJoLHm6nA8d0x/13hFunm2Mtq/phA8g+Gn
IBSMJrPybKCmMdFRCFQNWz+YH8jZeQi+q5LFtN4c4AZ41XGNwysWpoTP1T/rTj8SHxi0yA91WrU6
S9+HTw2zEgNa6NzrFSXwX1pkjgcVarM+S9cfsv8mrS/6N/jo/yfXCRnnkH16brmrqR21JrF+YxB5
FN0tWVkVdh5qbdjJUA633oH8W70Oub01N0ZygNnZQtRnB1iURy2V0qWAuZJlV1vv+1RLWMNwVKiI
n6kjtNyH7+PpLn7r0GvvL0Us23lDqO14Vf4kMZkmeEXwY0jgXE7BCMIglYcUibIoknSUnGLsxXnT
O6h2ch+EPDtAbMrlLBFVvYrH66CdgaAP7WUo2ydvaIPH8/viqIWQ0ZO1+JLAyMEtJc1UmydeoYDt
nYG/gE+pFxjEcu6g/4A8Eal5GES2l7Nld11p17odXIs/bxyfeejw7v681BkRjo3nytujwaZqGazy
Cr9g0TnvUuLb6GY8N5OYI573D2ZNhft0aeDoIqHpYa/q2lW/LHs7GLnTRZbpGJQwWsupaHrJxVsx
No3Joar6dSKmi8Y4gqeiu5Oghw0D5w5B7SKcv3Dhiy90dRUPLDwjUWABpLAMRy34kBH4kS1evrsy
y4L0R/i1DZkic+oLIcNDfJcsfppyPH3BPpYEWNmhVHJ3NkRonFbuEUgZuYszc54BfxaLNNhcJsQk
T/oWjmjeMP52OIR6hGy39ebJ1IykAPnMHtDY1rrnXB0+rGwvc39xeUJ1eZRoTe5mTtRpWxVzngk6
YT6tJ+2T4tJlext0mbqHFQ3mUP4mL7lfEekoBuAvFWoar6KLYk1MzkU+prrbT+G3gIqY8kEyge6m
z7qgEIXSfGINbYoXiLYMICioUt4TjnWRCMxD7U46B76pNuOP+WQfERFbM/p8HEtu5Q7H/9AtEWB3
pIHtxYb4xI/DuMeY74fRzMIKI6ew6W/24R4YgC+fmRJMalq45i+cJPwKqgXz2SnEyeKWG0AfPzrS
pg+Z44ezAWeMiEvB5OXumFvv4qZmDQv+U66loDTy9Vd7i6wE+gUE8I8ozlqgExcNNN0hFo7prXsW
ukibyIkSqnN2QWUlDuvJs1kjOLanl4+Kv/+0Y2mvEUwmSUA4A1YtMHJVxgYsE7zF6y9G3u2OmxnX
6eo6ntv0NwIrR0T3WLWpb5R/Qf1fpTd2BHoDgILuEWCrFq+QGEKfBnGSmrroSQzDX1A/4DxZPkYX
ln2v+wtOnYFi6pd3GQWnw+OqzG290SodeBJ4ow9vYC0TnB5+71QBTT2U6hPFvga3UpeYTBtier7Q
voGxJIBAs7GkGQUBQRq/UGZvZAKbpT+GTPeygHj5WgBY0g2xAYLGNh5fYynMxoYKZB/2qe2Uyvba
wxGZUT6XMEUSSe0UYbAjmOdrQ9TujPm5ZhLTReo+rPciW3rC8zP3k0y7lVt0yvTQb+CohH0lBpQJ
6AHi6U62WpuqExnChKBwtkb2w2BWI8UiHHHVSAWchNzXpUBf20tP5ZMRdwBueTpfr6xzNuCzgJzN
GUvb3X1Us9SdCbhfy+1wHFI2kvdtTeOjCvdYBZ7faP6w04PDmpvPcS4J8ZboxVLWhA4LFSndYBpz
kAhMIswSBRZmxYE003ZnWF4UCvPgsXb2gIYr5TW/yQesUKaZVljl5UnMUlUBpJ4bCBvzg4XOtDbZ
u4glxe4m855udYdK+U+HeUnLl6nXvjiN9zk7JajPpqcYlLILHLUmsWeoYr4JD6/a6Vn7TDO/YFov
4iFdCXy73J0Y9fCZ6suMbPvSq14v/mLUgfY/zkJEFYcsnWNmC5YH15IWDC8bszkQCd5tEwiTSGpA
TiaMIW89jREyExvBKBrwOmhBwZrh3vB0M9q9/8wgXFVPFFjBhTa9FFXLiC/34zAwG8Q8ZTDIoh6U
irqurNl0cXKs1zM2E5H+Vy07z/twtbXfGebZhgzPR0KcDmyuRhpXismzdZCkklw7uOgcylsmzWGO
Df9Ho2ovUtjvSZwzFG2goDUeZtoY7mF0mp2P/ti582kY854rca/O+3Fie4s42mdkz+7Qjd5teMG/
EjBvYjwv4/7Im1RGhxYSysYMTatm2W29HBXXJxcMBFrry/yqCtNmc3B/AYfTp8x0LLP08sUqqG09
bhrmOnJ8EPMBCzXrz22jIrxM+fPT1yy6Uh6vrvogNfJDIzM8Lbn4XXkGK7n7etM1Q0hDNj3Zo9+t
DK4aVdJfgo6JVQgMBFCV/RFN5PUixdiMQCF/EQ1p3Rnki0Hm2dbP5o8aS44k/2LQhz+a4Q3ccjO1
lDTvYDdQ3CD0m6/Akn5bXzz1DSeAQJlbfk8mGwhmmhZj6r7Vw9z9Q4RsY5QuFpB1R555MHZGHrGv
+NRaAtzbGMEY1XRqevHe+vKRFAIvcSFk/1nUiBT82y9a4o3iOENBWARAf6MHSsWqmYM6U9DOSlt+
DCg7vIjDAmDOTtH0Z7QKXchQAvo2D7godv+7d+5OhZKhvxgt+36K2G6Rr2quhapPd2u2CHEN4rfr
eEMCQpDRHsigyKtOIhB6pvI1xPdffC1ZACxN8jDrM6RK4/NdKdp2OKiRfa15NcubgSHOqPsef5mD
0RD/NbDEY7+SsbhCgEpOxgkx3GMzOehTE7XObu1pfqCHHzAD7j+R+16Pno5GF5rjz4U7+9kIGUsD
IWh3RcjZBbzCa2vQmB367Yl6xIRRDbNxByacQr537ZelixM7vDWe/Sw/GL2HK7q0nGTwH8e3WihV
gi6Q2m+wAYG0kKkgGmrq2V4Imj6CCu6qAPwhtt7D6qmQ50Uzpq8iPVvatuQW7Mw4T63HSi75riza
OMoxEbHAVH8T1IkTVRChn/rktPJDgptwlZEVAu4lICvaoj1z9ybMRtSYylBY2l2TK0QWLPaq+dfV
E8MoPI1riaUKaequhoEeECQmT0BeGy8jtaqhv8kr9cETn5GtzCWXD1HmIrvLBshghL5dklrgJoZs
ZnF9CM1sr2wjVsre2YKNFlVH+/ag8QDig2WK69YI5yo+nR2otfGG7++1UQmf/NRwSCyfTMPXuAPs
NUHGUpa2pbGmqUvS8IL97A8soWuTru4Z7iW7GYY+1eN3fRGwVrhAmyl5sQykfHPX3Kb1T63y0cC+
HE7s5Sl4yG3U3YBtlOeUQyokhJpVyZeVeVl0xjLlbGum2faRG9eq7xA/fDlRBX0Q0E63URdVCwdz
4dUSa8SRThCXsBY9hGfb1rfCCDqhJghxLbFc3XSG+x9BEZi+XT3pTJ7+UBzbGPMkDIN9EtZJ7O5Z
j7fG9aUV0fUccMy1SAtKiPkd/cukS0j/L7jPuqbr5mDmP/aHofZhmapxE+XsYNYv3+Hgtdjbsca+
2RHgY/nN/CGYSuN9b/zZnzvjl/kMjc9lR0hpkVQQcz/VtS6nJpsB8OpZZFaDYkExqovw5OlUiTJ0
Vz2pBHjjSG/ANidYsgaUN1CSVu0h7zgVeVJM1oHAHRwBb/Tz7GoqloyImHKUiU9BD0j8MGhT6yk3
okbSORfV6k0BlmgbsNTpx0tbrxXSsflOvuCz7i8Iz5WO+CZpJoWvH2+arPlKzjKjfVIzwSual99h
3HNYUlUBFFmG2JqDr1ekdmS6d7rKNBZXM8MewRQmup8PbGi4/t6hU3hONiA4Hiqn6o4i53tn1f20
UK8IAqfl2yFTIE+JmBFk8sEp4bp5oKivcsR700mPR6uKBkaeDDA7mzcPbfJDeUo523xKvNngUGyu
nV1EXRrkJ3PXuTBOczHbwdGLW5F9pVhOFaIeGNRTine6xnfN+Sw4ABF/0Nwn3qLuZy0QFsdaUAE/
Vl5tFvcbRuZpsB9i6RmTi6dsGUimDnIA1XfmPNhMDKAjG+yYb4TCTFgWK7aLdD5+nw2Ht4sGlVvg
xY1guurdrRL9/EDoGRjfZQM/8IZpPGu2pRW6ffrt70oV34xO11IZS/X4MqKi1G6fprwK/AAv2sya
JSnh8hmrE/XXDLQEohXNbBILx7wFHJnm4/Idv16tTwzgRRdw4ge9EC9p/+MpXPm1wms1Axag6oSG
/r4iGCS7tRsp+OGRslv8DcsHu47mlll3GMdcNTs3CFl3WgbjDqtucIfnSKK69iLHkP2h+eVEzr8Z
Vw8PVYth3/KQz87s68uX1qLRfFdurxSTk6oOxZJfptGBCNS04ko0HDw3n9iL5LDtkeJh+Ze18WG1
5Rpc8howzQgErNNPTxi+/JsJdBMGrEpNRAoDcTzHNDAhZ/AVV4ghjtDhPLFbxCX5h1kPVBic6kZo
phVliOBX0IOUVkapyHYlN+psnv62D0pwUagBHFA1mJf1jVOOwKkM2WwsxgC8xpS2Cktkq4ZhSs8k
ih0BqDXK3CQ2mXT/MN6pmjBTOgu8io880Flf/lTxSN8DPnxg8M5As/p3vVAPpiF+XVmzcPLANLNL
v0+1ixh+hIz4RZPN8XHgU+wp98HMQRAGPGFqqTxswQ0mzffZ60NptNbl/7rvpR2DMwGnFnwwrMyJ
CLj5CZB+Y911MNCXE4/fQYWCJwMl3FXR/3GczVsaCeTRE7IntWP68CksxHQHe9LrKuXgFzaCvZ+J
wS0M0sT13Lgums60GXULBGsWUFcFDlZIIak0vWUR0h7oBTrVSXaLCszc4UUJLduL4Nzl5WYhdJ6R
fwCqjneTIyVs1ZT34zuZ9s86O0sr+RaicDF61Z85zirlLObSJeyMiHh3aGTasRGVas1vgcu262vv
zmc7BPXztziOr5TmgMfku2QnPUX31bHpDBUQItv4hWz/X58kh52H7KyRrPDnn2YMBVudrGc2XTR/
dhTFEVEM0AgkbM7KE5qa6q5khMVsyI6tujfczDy9mHhaqgWa+pfr+9aCwuUmIguckeoebMuAcb//
vYIB6RJgfIE4y2j5DJ4uqoFbfH1OROm9L5L2JP9nqdsF74qSirHsdFC1DiqIMAK4vQPS4SjW7/ft
Xh07ArG+BfrswmQUEqhRbDncJzFg7Va7L2MkXzb11B43HWifO4UW2xYwqj8pAXDf/46Gjda+qSv2
YUp3yU/69QoJnGrxZ7/1vz5VdMBEp6/ig2vhmAngDFP7NQ+Vg7ys6+W2Dyf500aPxaRnvV0XT4TL
HlV4ZM2J3GCLO/LTyNAkdPoaXEl34523QW2jcbeK5EMMtSf+rw1c/kr7p9xbdMYuqVu3QIwwSDhw
wPLYhWicwZNAAQ5tZIpa5bjauQkMBK1C8mg1g510OrBTs8/qRbrdQbqaU7MTZtPzZQVfYTL5lkSq
Xh19z75YotFx42MTs4ILZfcVfl18kotCs+W5wjoC6SK/L+A3tntO80YnKIPEKPNS0mjwmOjlgUF7
pFPiFrXzuActkfJZyaPrXDhzK+kFC/2bBxxF0N14WiTLBf5/GUJ9qKeZJk0dJUNL6c+/Hf9T3CLZ
LzmwMHlKaF225y+5u1KAdPQPXy15+5vFqbYsaMQ76nPqBSpxoLmcWoHetQX1lZLNQ3swPhbbo0Wz
hubpcLuq1nwCM5n972P/mYATZgAKgmohNBT2PEE7mnz8Hv+FWoVFjAc9JeA1R35SqLZHZmPXMnOv
Mvp1+cxb9VYKeZSJ77PgAuXU02YShyelwq50ytvtenajTHopkI7MCUic1jPXesTlLeLesREkNma/
R5eF5ENXg3GmVusSVSsiR719imJtLUjaID1RaEKKlBakFCbB46BTVCTr/IxD3hodUTs0smdZ2cD+
gDHt5P2VhJnyltOYdV+D33MtmC4woD0c+v0pQ1tIrp6KGt0poA1FmfCz7w8FPWbtdZBh/oL2ag7g
AWvqpMBXp3iB5aOEs4eUpeDEFj9dkLDri3LHY3GPIRqbK5Ni03xWqRbWvwlwap1b9aeNGCnhtiXi
AWnRBDOzr0VG2mOJSbUsBKqo9idoZBctFmJKYNmHUFYo5X/2K/Ba+i5xtepOrG0lfs1APnsu35bI
0Q3nGfDVfjOPM6YDkPGN/U4m6LmRdMkzFg+2wGheec3lKTcRShqXL8kbA4yfJ7dw0E4Y1xAn7CQm
F3bJHk7fuGnkFe4CoonIS9SRkT5UEumqNkHn2AMDaRDkLVoe1Ix6Kowav7ltWOnEfS5xEB+/SjmT
hK/Lkuyoj5OaiLyZhI84KqQzwp22D6GDKN3+t8AedWUbio4NV7ON5FqU+dJ0e8W8cL62QZNyw6rU
FI5/64yENRQ7EAB3qDZGGZl2vb1nagJA5uiNZpczt6qiVgUz5OqpFmYV1+jjugp0hIbE8NTlsi0c
dMQ4dZK1Y9Q+MxMwmaNVNdxNzxwPjSVa/JawxmBp13tTc02DW+xSAVpGGiqDv6bYk1F+Y6OBxrfG
Jsy7NAkMoa3WACTT97ds0jKCWT9kX7b4Yy+mN2q9nOmvhkLDKtKe2E6W0auH9CjGqqMVNwho8CVW
XH5S/npWaVifA3qflZDJFrysGf8ATiYUCf8hY2jBPWAHQLKZun+ZC1z8D/QGitllUszr+CjPC2fd
OP1XqXN7JCDBTKiVarpfMrZ+nTahBFzpScNq+sIV6X5B3Cb345zZ9VflAojBlt8APcjy9U7eOU7O
ov5ZsQU2vdlIeOTCiN34IfKimgXW6oEARcRuO23N8YdIL3Nv993gSoO+l7E29KdBCvlBD48rA6qy
vDD8WrRR5dpRA9QQUF+0bx7HxPfUszl6+HxH3PryMbLPkUliTKxC4IcAFuyS4xmAj1TITqDkWJjc
1jOH+CNS1KfEgrX8nRrwrKwliltV6KAnyry7FiOrxd79YGI/YOEV4wMxq2vjnCidJ5aJbvaRIZxI
IbiYH+VK7b4y0CJvn95DBqM+PxV25es44lZ9Wk9N3plEVHB38oSMXQhB0X34aP8u6mhlO+PrfSy1
qPx+vC+EuzDzXoHfLyMIv+r1/dDTkOv5W4HT5Q7Fu7D+eFocl7eXBZ4KQpsDkJBk9wUmwHse5lCp
VnzZlaAugAVoz+c+5ajonYyJFCTG0EW9mui02h0fe81TjheyAZx1XIUvF+Ys/QswaDRl9bGPwmip
RZsDFqVXAn2u+gxsmLyxNLSog9PU8nCKB0YKCRWbOiCxBbR+8EGxN7oalLd5C19cmMw4SgUGnUlQ
HzLKpzBNd8BKibUes5MmvjsK8w1VQLXDriljr7hYqNeZKQ02EMDwBqIoZ7L3r4ru5xeUSksaOc9K
mefCi5FAbHfYrL+m6a19ZG2ijptkp2qaKcLivt48U0UWLPXnp4eI9js3NAJSk11VezMFP510O1wm
X3YvtfYzimVYRKjCggi4aSdW+Gv1oWcBhAIaivYe1B/RXM5/B16iKr1J1UwXczDUxsnJbJw6Z4oV
4lRgQMf9gUjMlBCXJLIgb46d3/tkAC55KTheuRMLkavzWZPkYPPW9YYst7DZlYe0XaZpelkga5qu
gxnUJ/YEIMK88st12RtM+JWdXdLPGf8cIStDUxr7nvN3mteHCxKvwnuOJLvAzGmaxmuzF2UQi+gG
/OyDjayMCBgmjz1Xy2XaqB335HqHMoBaQ2wWs3G1ZAnYiIsbQsV94SpRfn38S4V/OKH54wYOIPmO
Ob3iV6S+h63T7JTD4fY9qmRC7goo+eYDq1KvHflDejVnQadt83786fgsvghYKpWy+e72fFs1uGvL
dOu0EXNE4NENX1khdNzCtq9g7tq9CymxlhW/M0w+g9zOfb12SLpW098vkr7gFYhpBkhWsaqQRY5l
jVFAqpbENp2yBxjkHkscCzypANuSJCx2r0Nkrch5RlZ3N3kgQrN34HeLIy6sE/dSXP2pnpgT9v6G
xzkSxC1imgJ+4muASXgu3n4UObcjBtwOcKDIQgKFH0i8UE68tb1dGDahbQUz7w77lJK/Zeda1kOQ
3wgVN6ZUnZ0RBBUJlqVoUHq4DvTRzVWoQzw3YK2K4cY7rX2nTxYYR7+r6WDGz51bsHiSOkyPgqkE
+jjzBAN7bp81y2RODOZYZs78wtGyqO+LHHiphAwLeADnccugl7vj871flWxMIkQbMRESaDkT0hRZ
Veko0VB7cR54epaaaaPxw1nxYaT7YU+hrjS/TzbPr9PmF+v4nw37gg6K8IYwI3plUhf2YACcJIbF
BilKDAN3GgISp29oQjTqOYyubbj5NeyQpDbxMCxhI1I9WmhoBh7WuXsWi3/lmUqm6UQjAK4qAWZX
AlpvBh0sGhDlr9IoNrwrOb0Ni6DwxkD2AGqQzrI1FU0CUZ4KZ+/XgPObPAPq+Yvkr/B7wrHMsJH5
CtZ0ZCiz+Cqk1GmD0g+ilhXlVNc9O6+/yV2/EeOuHZivC5tfpc1XMxfXIN8X7h4vQ9pMpCNCQ6Qo
Vyh+O1D9NEjHQi9WxgzTF1VhMqz4Ad2ynqSV34+aFqVAp4JrsCIxBd2ISq06xistAfpBbUtRU2yV
p5DEn1y6b4ojDOm2fDDXaHtzVqLSrwGbWtV83PIzK+ip0r0/LA14v92JTVUa144mAdBmDL/zzqtK
yoJvLXLQJUwF0eRppKoEvtuqTNwUEKg5wkfX61ofHX2s/oaOCid87Ps2pchA0cqyHaNv3bnFRiZ4
LVQWwdwFNSQTnbGL/NP2DoGqkij5aSPQHC0rMk7/TNjQN6KHcnM8Tk0bjprMJKuQlXwQ/d72lVce
QQ44V5+E4Krg8E/v+E6w4pYC5EPdi5kDkVKlwvgLgmhIi1GCCEa+GIIdmD776VHuoxSOPF8lwpkc
ErLWWbDKH7Tf/M1hulwHDjSffmTFpw6Tvk3I9x85b03GMxnY6j/pPBSMsfFCiaXfMqoY1hiOGdc9
MTpDane39+g+P5RmTI2+/yLj/BamSIlV7avfAVo1310xe/QXu80rTnlonRPVethFLzhFQKH14/vb
jaU/0mCQ2xQnJ7/M4JRWF/NLs332AEax4n1gyGxQlgZ27Syg4k+NEcoAlLGSXTcIt8777imlvpSb
+GME/iijM2xto0WMHUokiAs3PLeitmE5lbhQASXu9+PoFqHEIE0qiFjTc3Vc/73RPcIlFoqv0Ui+
cOUAEh+cHzfcxFr9ORVcND28KvnAn3oybfDjdLpQXWixEp2U3TGTMkOh0DoWlFIS83G6IVFbExCR
EB9i4M1vi7bYAy8ZQwrN0uO6THqssnlUimm+VvwiQKPHw4VSGdB/0Vf+MOEEsTACZ4naZPOc7JbL
IFQuYUGJJ6bSYRUzPjwALaGY2GZC8B6o/EUIrPzC9hbryeZ5p6qjrLV1Gx54vJUdZIs94SEDVtRX
ZwyNFy4zfH0E+fJf3U1A/0safS3NK4V47TLebAJWPdI8ZTAQH4L4VDgGNuHHD6ydN+KicLGOuSzP
m3yyVpNmrK5zpM8B6TlCV1De77GUVX8RlL74i3h19et5vG5jL4DsXqcOy3Uh2u/2utDuj+3nRXbr
fQIunk3PPBZutJZzViV3OYw8H4E/SWOqaa3Pj85emVKAvjLIDb1olXtDnIEbxEDRbAwosUNWGfgv
+BRLOG4TrWs41XLonq2nFW3kHO1zMaFmwk9sNbmgC2nPYGR5QQUjNllcNcvMRcjxgbwSY0WXG4vY
f3E2FtPCsc+RjZuelb3/tLlGBY7gq5pFZ8SRtm307scrjHmyoa5IZkpwsc+jXOxUU2VEp3Z9EJLm
6818TLr+yVuZcEwdGfd+/rijRJZ45tm1cRAnVWckZr+wM6yJJm+LV2DdCD0dj/YU+9yi13mS015Y
2M/PXB7nu2CcObP5C0VyGZu3mBFUv6M4yIuOXgPxIr9ew34GPZ8vK7v5XKkvwWQYaFFvYkBB7e7B
9lptrkiKFlHwiXT7sM+fml0zIRDb2BBuEVMhbWqwz1LaJBQp/HHWbjBN9TYXG6LRVMn0NcScH7Ha
ajOTjPuv6cVZCcZmh+vY7wy4fiP+e1tMmVYXw/XSTfAZOSI1mNO/SnNgPgPGnhFZi+rqbqJ0jj9Q
hHtxrJ4EHYZx+gEKBZpbzlzmMFXh9t+Nn32/aXmYiOE7HBYsNf3/8c1J4JC//38dnhvdOiMLC8nk
lnIY5NMSEp+7QiG1YfypJRM+QuYvuJB+DYxfiaohG74MDUg3MT0BuVF1RamWHBAjbL4ETzxAQ6rb
XFnxCmy3tAWTA9DRx+6VmiBdvOa8ta6rkdKISoYTZ+5bV4yVucq2jBSn16MtDh+coA+vdr6xj5Oi
iIvSeNZlskpZTla5nutAQmqTjkDwXh1ztRvaKLJK9HyQMYashRL3W0TYS5O+6Ym9b2hGhzHCgtgY
l2/tEyCvvZY1Y9a8u3xHpdy0RBQuCv5K997ey9c6zNRBvygwjT3VDw/5wXlvcPryYOUs3558vWQK
JxmjZRnICc/rIPh3yQwBSInsdI56136gdgBlK4SoZBfaPgg9LKQSam3YpajW4jQuYuBKuBMm7OHm
pWOmxuDklPxhzwBj3sqdE6iDgt0eMOHcj0iPbYyQmxIaaKlLMQAux02Q0nd+P/Jy95pqNecFwTQK
Htzsnw8RH/eNwqQxnfxlx8ajc/k+AtPyQ62dU4DN52QGbTu9UP2NAVFD0gvJnGY8n7xZw/jGXInq
EYDWJY+Hx9QCXyX4EiASvQXjL8RlHGFbG0ws+Avti4mHzYH/vonlprwhxxzFs+tgI9J5DcavB4ot
sOzkr+TsB0L/1qEBcnojYpOLpb7/grHrQR7m8s5wtKp1cjjEyOIfr0cDGsjos0JtFfxPTwXmzeDv
EI/oOgNPwKLT2F06s7SZKtyxsnpFdxLVJQ9cpiIcYDJkKiUWFcmm0CrJTa+ushcQr2W+CtAmxU4c
0+Dh7Xly+cy+kzgWfc+Uov6WSN+6SAZIh7a43leMqv7UGDt6nKkWb5UYLMv3Wqixx65AOk882KU+
+x34PrNeKaHrqJOwg/Crw1mBq7woX5tNajfMGe5wM8opEb5UG1BnLd9b6X8vfOJcclpl5xfG5WmM
EVEdfsH8m4xkr2oz5uSVZGS6ZW0gGL17Dkva5Ea3GIKUp0MCyNIDWu0Ypjaiq3g/OOfMTV/IBZyv
Jkofb2L/YVsm8cJx4AXSxkEGZTBHL+E4VCxcVL0v7W/Xrkw15kRNUTAeb7+5e1vP2In5GkpRuwv4
iQFe8JJ5fpMrBpXvH0WHMYxNAjWIEQfCWSKLxzH4oFcPuvNqrHlG/3NuF+et12nquBLWE0ZwRoLd
s0tF/YD2bukIDexknsvHpstq9nITZXa5ZVLGJAtCIb2GSWxs3IGs8VyCu0RXuTiz9+gaM2Apy8g1
grTuugIDLtkFNi04v5b4oI6zWJZQGPdQoV3Q1dIGaERHosNp9w7rCOih6agfIq401QAlHxKMxyYK
mla7BGrLixoI/nrflDUeaQqp75LV5R5pXoodDFWPEeZ3mNm6TYjPLLSOeGeqK5KLvvQ6BcL8fdd2
uuTKrnAnaWn0gknT/Lzfekeul+m7S3olE9FZ55K8cB91QDg+9efrjIMjrzSjkayGt4ANuzOXLLck
8kp77G2EZWLHYN/MrRREAnUa9ysr7ZZOgJSQvmEVbMRVC1kHikk932gV9NqFkquXv3RwAj+iRRT6
3n3NSwsuwBHPiUKZVgsECTKELY6qgHofIJlkbaNem0DjLZAcZVA09nLvl6/kiJeq2EMBaX+ZPpIZ
Uuj2MR5IdlX1MFvZ5cbKiO/GfnruPDKecOAGR38kVD5dCRgIKaEUPzYWV3+jkJU/R2weidVGn3/X
Zsmv0W4W1xFWj/48LeIfA0HOnt19p4xEIWBVUfd/64WLw3gE8IX6DdMsIxa3uCYw/jBELNpvsm1K
yf1e3ZxOxKU5QqhtYKC6hivMrx0CplUegxpCNrarZDb0BJ7ld5YvU8tAseeZdKClAL5xkgQ+SBZ9
dyvlsliMpqmkzgTF5hXGvszjbESBpHRJNFYxPBLmi3l8gp4BM+Ub1eKWm8yrGQRqCGEiC3sayghV
sB8SgeeKwpIygKQkF8sTnWn97gl2BJJd+zW2wyrHZybUlgWkAOLYjuUpJerqlRlcwY0gGtcQZHMo
/6wb7Dp57LO9aVd5n7cpxrcWOFQ0PmakF0s3IhJWzG0pPTk2S76RE91LHfahB0yz1AJvOgwdkcS7
QFEyj9d8JVwXJrWgpEWsCbG109RJZ54pXlUakI7FvY/JDkodRwqbilgJyqnrXqcHl7/eB049SwCT
qOZ9iLJYFbTmeBZMKBnEJFT+T5FCwxQAeILYZQDgV2PlhxULVNZdejOVsXgoSwtsI5LNLhjWH6Er
XNLm7P6gNUeYgtr8bHE46uvGp3tBA8AqrkAbn1aAEnZzHWQa68ccxlPHMeQ/PRuDURrHnZuBnAfg
mG3r67F5rllaittEW5nGGcgEch8gD/yC2Qhx3UZh7UaZc8ytetwR5dWH9TAuFBR9sLCgcqqlXjiA
G4vEr/RedlNZyKWXGvXudzdbkgXp4XeBtJO+0gXznH5Xg1KgNTiOg70HlQfktz1oxtu+i60Epxt+
mcFwk8PWR/P2M0iPyqOkl8CyXlWN1ia4UkuuR4weHfigWcy6xi1B/ElxTFrUPscRxjQ2mpwKC2sW
5wxGnG/UB8NZUZBsHE3S1Q9rdpat2OUk17eWC3eWA6nTTZ63sZK6q5t3MHAtXJOoaSSEt62FeIIh
7LJ5nB10K5RP7W0rA7oC5qhsP7zUV2rqLG9gAljPhG20ePkY2z+i4Bb4uqFNxe/NMInaNW9yjBdp
xByKllbmtDXSqVDKdTjp2wGYzA5zjBH42ytJ9lUBm62VEm/Xi5cdQu30uOImw4fSPmll5KwFzy7y
iy5dDiRZseU6mzJwj8ezvDL/IHsNjuRGgdAliiwCt3Yi5fZ99vi3GCxCkrWcw56sXhCnqHbfKra8
iJg1QklPDZnZzQXbU8sGbXFTisglTysL4vKQiHGqhjoH3AheOj+KKOuwmVlFacNi+ght1Iwnzcji
oqTdV5PEZ1nAyLXjEKpyDIbytqtY2xUYfkcaZUIbe9o7dxQs7ldKpDAtYZyfTEe79QYb33VmdBAw
xWvg4Q3h28bjzhyGCAtc6kGhm6MRGcvbTp1rvT3mJfMd4fGI9fmmyi7TjiEeoPBVYdrP1fQcClxO
O6eyJq90n6MGG1M80SKyu6+Qwu6jOt3J8PZ0V1jTIrTgrckWDjTOQOzlYCDozLkpOoVmsW3cib3X
9FcXvE+CgHM+dBa4M5RkeQuob56oRfwjqJZMUAt0X6bJXWoLo/54Ckh9k5jDSsCKrWaa0pZrU6Xl
qh+831Gw+cRm3NgYulC5ZfRIEPG3YdjzzL6XdqdcTX3xFfvml06Ppxey5j8ct1DwbqgKq3LgENAk
6qJMY2e4u4qviT6hppf8DOxhW5RIazP0gmQmT3t9MlM8bdIBjtxz7btUzOR6wdRZY9VCA2nm6imD
9ayAWQUEhTCoq1chekVAdn3juqhI9QJ0eqvWDxWyfXScjloGMPn8autTMvHzfuBOZHPhXuVjSzUP
loVMLZYpe5nxHHOE8rNmMJ7mnmMx7TIfBlrU2W1m0a1zvS37wUg59g0dfZ0rBXJM4LLxUZsMZybU
Gbmf5XUXeN+6Xe6+ioVS9l1ev1FiAYQ2NM0K0V0iTGN5MSSy0hb8IQIijbbMoGvDNHuG8t0ZQJcg
qLvMWKReQp0tkwUggf2DrbMOMHIbMNNd0Vhx6siMaIaFUqYWs5Jc9++3Eg3QGjKipDLzFXNfE6rr
oz27KvsIGM4ClbK0xrpWX+yYl9IqbYrIfTt+3g9GdaqQ9sgH9dhYzg8Un4S9GBluu8Sm/ZMye6Cw
3Lwo3R/Ko+PalCg5OzT03nNjecajEHcew9HRYFZGDtX/k3Uw2IRmWKuZ0olDTvg9wM0Hhgz+jFKV
I0s1OF9PoDWahgOCZb3IPdPbbXKDzMQr7dBKHanaxutIz8uQanrXaIsU+YktlZ8NM9qDuVGANhU0
Cqj9MlSnnnOnGCbKtLJMXLape+esu6gG1Zf/UsFaxZRb3XZlHj7fREEpBRxweSXPDtcXLo3qi/z6
CRO2b76BgG4gqvpv8cNJ6ly9v4ezduTyoSaj7gyu/hleVXuhKRwMBxlWtbqURzmHKaNSL+hoLJP1
UOquGtVYogQb+SisL1Nmb7bnHN1Nw7Geahk/WvIzkG6WI34UCk93Vart8dYL5RoqM//46lgD762u
Wsw1D3SrvMPTHyQckXL2RcmpvS2NzcNNyrXnkk9X8nK1V3hJZisl6GQv1wcfL+VHwZ3wNjZoswBN
c0ytJ9DTnrNXL3Xly1OIC4SHuG5OEE4UTJerNdHTpJamldAuyjSidZE5KYzMD02wKan8pqvLReQA
k2Iq9G52WYvLcFkMor+k/YyMHYzJ04KLCxoG0gW+atTUF2EcPXPBPaSBoR5FauXxG0ydU+AdSEQQ
JoKkMAyNbHImFPoRCh46oOZqfPrrjt+R0Z2suZr+zNzO31RR7Uxs/oG9bLVMrqRculjijrPHmjWw
ieMuSJlLhuIvX0ILKk3PAHjCKx7S+YJmGa49pF1Xu2wDMLDf45epfwHE2Hkv7ThhFqacToqxgZRA
Hv2sxEnapIlYTEaGQHKV1fY6n982fY+Y4U2Z0HqohRPTRarcml8dTs9UB8Rye73O2BmEn7Z7mYLA
EZXPn5Wlo/cOGSkeh68svqZgj2xXdpbRwPly1HRzOFnP9RqqiK2utUvbWOR+OfHvNrI0DdPec4Pz
vY/Pt+EvGWi5ko+Yf2uHMoZ4ycoBR4cN/PFgvaRKaemBZqmUWqCkU9Ykx4b1uFnkll57TPYVCRL0
q9mSSggYWIDM3fXK8bwe0KUPSqLMLyrPZnlNbmMced4Bo7mSArMRD2zeXCr6X3M4IbWYY4drl1o8
jtoBnDwvb34NL98e+9zKmXAn97HPxC+UUHMzlhOdpuCZcfvaUfGJ5aFQDbrUcWWxp129gEwDs7b4
KWmWzNMImPnkLpiVZmFu9gD7JnsPoG1e7W0EHEwXAz0VtrsHkjHMGE2FAeFJsxgElNfPyY4aeAb2
JrOtIAEh4nVBw/pxbh8HaqdbIn030z9mEM9tkHJwtvhu5u8Yv+5HTrlvTuvzlGuodT54Vyx6dqed
7p+Brn8juUvhnef4K3by8lLe/URaO6hshIx661kvwBvwhGDjI6FhihmWX83PHaBQwKoK5ko0NFKc
j70J4XCzke2CMFHj7OGKARYoro78G+kfJ8W7ALZCNzt/uX7aO/RF6l8bMpLB1sBhqruatl50+BoI
YFbkWHZcCPGqkEHGT6vtWUKiW7ZDdStxWwTgYNrPJqmfx5wv/BUiJGAHb8Rn6tKJijGJmCDtAYG0
MvEEIMstwnOjm0lb1iJsI0GlgqFK2XS5BnIJuK/E8g0QFPH+06JAZ/gvcRGeCtFl98oTkOTp5e2m
EXbCBAjHaNKSTyF/i8vTEpV8js8FKsxvj0JJ0OMaOzkjUBysSfdSXGRsoj+uJHWG7maBYxdYaWfv
13XT5PV18oAU4XORqjGcM+Adz31N1S+S9xzwJsX0TDOyOS0/di5r7gZ4Tb44pyXnB3bqLYaryHsq
9GQcCuR1F8OICenjzpuu+hB4iE7TM/lBcOhSKa99v1aUtKIsUks3carBUuc11XFP/i4FdxtrrrV4
h4k6V728WxDR81/M76qFeji8D91BbWKuIql1IPiOhK4+t0N1YWRekP00eHPwSFLsA7rubYvk9cQI
7ixV5l3CXayJb2xa7pxxGU88f1+MAN2SjVbBsurv/LP/Sfbf7IeILD7L/HX4VdzS7wu2ZvYOPSpB
Lzjy2I1r+Bbh/wN8R47XGtXSwMtRKEBzznGn+Q5sGs75jAIr1ybH4vMzB0Jn2HRASFrduQZTa5AY
J/cVtapeazCgVd7EKhCGJaZSKIhqfg9x/mpD6fYVq899HnX3ODxZ/udsok2U8CnOJ7DafuAVj2o5
0wWAJ9Lj2rbtH/d+bO1fKuZiAZe7cQOUx+n6GY/yBL4f5tLzhKd5FLjeqPhrRnbg91m7EB8sGCko
8GZY3U3qy4AZzK7bAgM40xYyoQIpDdnqxnbRJFU0QZNqi3tK+31CPUfThppdsSrcOqlc1FFy4mrh
T8qiBvKvhVKWc1tF82a1/tKnY920wloCx4Yy6hZsvsKRqtV1tkxcLmLeFn9y+Vjb+jMGaRt/bD0A
ITofuGJrcoQMjq9qSJ4M9OgJ9U/siHlnCqhala7j3Qe8bDGM8D/FjbFxGAP8kDV09tVlHGHW2Tyb
a5ZbE7vSZ2PHW73yCA+o3pCi8+mTHD8JSb1blcoqpmv1QR1JTDcFjvf1bomFb0HTPCiTwfWnK77n
EkTpVIVgQTkDmmnCTxh7qqDGM5SlB0fHS95BUBoRSoCNSIZYoN+IAayVzIU0G4YOCVnebFTtm67A
3E6F9uT/P4LrwkKZBBUtO22wJDakwpkuJ3WwW441zRQrTymz5z3vad7CQTnhWZvHNPtY4y47Q1nC
Z4L8xxQsABHezIre/ZB/D3Po9li1Co/HiK5taFaYMfFhROkuHCggqy65hq39QgXMhUL2QqJCjyG+
jt9B3xJhyGRz7vGHxw1YV+P372vnf+pnlPesPbBNtmwCLVRzCE4rFcHyeXgqIpJxTBscT+ahn7zj
rObk8YAwlHExI3gB0pqL8kq4n+iFImYpbQWvXKgDjVUHBExD+fpgkUbMIM7Q+OMVlFlKmuAlmME9
xPgfiu72xAb8QUoyMSodRDhcZJC+RNfDD7djY5wdxxrvKdebQNOAfNC6JyYBeUb7xQUZA8vYfi5b
kzH2J63hScfP1omCFpkvauGID6PmO6mfUA9Q3C10VcjBSZL+2R01tGa0MmxgEI1dxg8ueLf2UgSt
Piol27FphhVfin1Aa1vXZGZEZMARHNvCqJFUNtjiNheUk/8wd60coUKku3d2I4tSvb/6Tb1kok/j
eTyxJNuIXutxtOClkL8hDJNUKVHaJGTRfZv42pIWnWlBMnGVxeFPAsyAQmocnq48uZGa09Z5NO5N
A6gV2YJ7N6F0F9MApXclJUieWGpJ8AqNL/3JbChyGDI63yYaAn6yPy/vgCqojqYcpthAmDIz2hKy
fkCdwZ86n4hn8WnKx7Ks0Y2HXPmH8IjOSk8D3jpL0nWktITs9QwXCEUckzznGwB9IJ4EnEqKtdhz
c6eQCwtGQA5uISPEFxqGAHC78ty3HtoDhR2uBD0E1gVI5pN6Yss6I7iFLT3/xUf8WI/7zeyQE0ng
qvYAEGvzgJ/2T9j7YuhqyiBg78RI5RXPDrf0T4UFt73z7JFD95fFUoeGNgoMqPdkFvFBodlMyAZB
zILLetfVeLz3uKS5IdVRGrOBBEKNzTf3ieEtTBpuvFpgtwxV6vp+s+GfIpgMpR8qkIpOB6NaSEpm
YbCxu/4Os6UoJsoQK64G7+2ntWsXEX7ETnbUvylaGAgz0uEhzI8rtlLnzTuwKw4NSb6P6Ogl84Hr
0+aAwtcmM88d8eE1akbHYgCt2jdHmLdZIEOc0xiAe2A29y12injzB6LL4S3Ix12Xs4Ka0BArpmWQ
i2L1ZCCA+N8Azv614PGNNUGKbf9OygLCUNkrls8jg59botVy5OHToqz0bM9wPEIQ8dpt2Tw/YmIa
aYGt381HIPUWbyLNc3zPpR0k4GIkR5txjgG8V5G3/ZpPYo8cSao1TBFYFu1oK/4AyGR9P10y1Zfr
qJrfUhvJoVS3+gMf5GyEoVffT9NzVcBo9dQJZcuqTe3HLZGblIB3SentDr5OTxZc2twzln6tI9/i
pqnnu0EEiGN7IREdYKiSMzZtbx9OzX7xnYN8Uu2C0+RKRCxr6xPxYlxpe8cw6DOF74aCa+2ClowP
VhesoMZrJh6qpJ80WTzL0dPQCBN4CIPPDgiz2/00yyxKRmthQgxdBiCwsXwRxzzoHLniIbsF3jEu
qco8WRpXWc+4wyZVuwtwsH6+0GE78a0Zyjh3tSEqffPekhMQjtdAxCdKBDpjRGqU8QsJCm1z89Ua
5/QXdeWtfLiDIIWxeB/DYo8ZsdPzOKVeLBgqhodl8kNMO7U2zqqZPL5daToJpe32ZGhlmrGJemmS
9c8NkU5FpzEKsgM3uEALMJ4oB1Wa9KJGx5IpRA8BIni/LgWCpPIZisrkeMB6WsC0Zr9l2MeIYSmK
liPXdja3nsoMCyBw2N79hJar0NwNN+S+jqWTbzFLLD8FSj6OY7MNJon6U8uM3tzaAcpSHpzqz3ew
mH3Q9hjE0hGzrcp0ZDRES7JOa0tLEJ2ExIouICpN5FSrYpx9iOnIu1mHXVAq0VUh2XCWkaACswpX
UruGbONP0pqZFKTxs8sgBqtyA+m0N44khaWfrbZJyGmM0IXOLJmOyySSaueNQ3OIDDQuAKR5mFV3
mXIB6L+jCKafuIMGFyQTHv4T28feGDVbhw32Qygj0giMEun8/djxH8lGkavwMTTlzOfWAkN/D1Qi
4rKARPbIv79Ajr373fqz507JxmX7KxBqzPJR1wrY+xg4l7s1NN5kUPs0L77T5dF9PQt0h1gsTO7/
Wqf8PeGrsfaaig3/tPxCU6VL4Q0m1XRkjo2R1GNhNPlMxmsxzdVviL91uGgfQkFkwus7xKuHfJZf
boZi7WNCembyQuURgna1+eoyJOD1SSzXirhJ3/kiQHKhRok9tQ3I2tLZ+y/Zi0neqz7l5lY7vxNL
XxMc+KgOofo5Cs/3IpQKQYB8OR/5oprYRdq3nZnpw0KxQd3LIMaEXylMLVD2g7kyqUxVPo0jOUlJ
mXP4ZP9tAVsx0tZqwdnbVCBJUCdsZtxjOAhCYNIyR9NRsCScVpSZH9dLILHzTrHTPcxeARAH+WVO
SYJQy1my5i9jgmW3dt6Qz7yXTFMM9COLHgkSCESrePo70cwi7Ri6UsTymVlINtf8Y57qHU3xuJ8x
imLogBO7z2KMM7vZJt8/O5bHHd+0uQa8SyGUQoHsb7Fyi3TNur83MSlvrnpLG0cakTapU+fgZMj8
0qq8OehBAbFav3cbUWv3TIoidgV86nqyAHVutafsXAmPSqku0O/Dj4emt2pKV2X6RxLQQFi1ZMEr
aLDYok4AwdQQmKCZ/Kxv1erVmmHnX+Aox3dFM2Dyht3R7y8zaazpJf9kceVMRJW45QseVCh5LbO2
Kivc2xuBEZaF68f5byN/oQICVGXgSmEHR6Aso3hhY49+G/S8lIlnNoKjLqdcg5vV3N4gVlkCqBdJ
w59bh1h+o2CHEnMfLreoTY+SjfIC9igjKiCsHjwy8GgUzMW1qWXm4Xwf1yCu1pjR2jAAI001jUAH
A1pty5zo3ulg8mCBHv884EFZRv1EZQ/OyBOdK4HDv78YG8MgRlVQovaXtpiPwkAKVwFXhpstAtpL
yVL++46X4ZOZks95CYyboVG8WdFcZmklu+Ar2VBPdC70W7RN0HGx82+EuaZVWxAFA9Jx9DTrNMNC
GNefm4Dorz6UwtTZdQF5w05b188S9nFsqFHlyitH58nNVQifffS/V4rPUHW37+4+uwoUXK1jyLdO
a7bNQpjFEbpjpM9f02KOr7NDB2YImk17DVIna454urxWtQSdcWUJeqaqw6dX8dpN+XBupXxqcfFP
havmJM3o+pD0wN7cfKf0v7zFtgyaWPcgtyn1Lnq2MKteqEITKvyT8uX+H+ZJXoJVD5gSaUFluZgB
/bvIO5ANORcc43RYP0TsKfsXSoEpFOMFXqdBgx7jWizmLEckwh9EWMPKCUP/CjjkzUCc0fOE1WYh
AI8fs82UCrCi14TlLtavpmdXN/ZA1kmQcyV/yAlVN4ABGy8XQuwZ3npIUpF+2RaGNejOQzoI+poM
q3xWu0ZXWSj9/KNdv0AjnrIjxmp0KyTttHYWJGoqmYdxm6mQWO2M6Kgx0T0UiC/1r2IYehjHcQdZ
gO2OQyQ++3lscAPO4kYP/6FXPSqjRzp5G0VdjQDZ0v2kEpoCjbM4D7B9sXVh7n3RCV4CvlgOZa+D
totwv3q8KumQQzjiMaswgwruqcAtcIy/mPlBzPbJyuSE0zkxsl/dgzgKzv0lF8tfMttSB23eQj+t
jwLjTTTQefwOkCLeJ0In+jabZJtF2X+zEMdbhPuzuOKxofBkEZjFd+wRM9VsQRafDgJFYUho1trO
u9rsWtkY6q2NVN7seHYcCCTZSg4YQF5j/Akh/lcF3vkiRc4Zzs4ztjxZMK86G9pMp+HrPIcvlTWj
H0XvPiEVy+0LQFI4IWAn5x52MmbicCZqZBuheYdungCjnqBQ49v0KYqAYpPzGOwLcIKk2PYJbfOR
UJoNddE6AhVT+DKeb8ZBVQiyXMj3zj1jH+I3ntB6kZh0y1+k4Iz5oJ3GNBfwXL8bQlj2IEbI8+Bb
1PyCpKHEh1MjqwmE9eYFJevrLxbERKI2VqxIVM+mzskZdg8Cup8kheKOI00TFc59UxC3GhAVdtxf
uhYP6r3fdG2kdaNtl6X8pIf1xSBnRthQ+bfGaGoUNjLM+TOLabwVvXkAXq1TliaCToa8os5gyFJ5
5z2KojHzCcdq5YkPc65OJFOEXkE1nnzmQIwuzFkjpCATIm89aWAl75b9wROm/jzZoZccRUtGQ+r0
eVkH3o+K5enoWH1E//VtDSNCHG219jx0cT+yMrexI0kqz7qsMpVmzZX5OboWmzFHD/xojEhrHLAe
uiemNyFdfgJqbkL7siCuFPQGda9fzIaZokgC8xWT5B2oelm6EkEWFS4TaNpyvFywv4zL97jVwQsF
q1LLLZYpyPdiGOhSIeEhz7zckIx4daZf0gPVw8s2QuKyWsrZJsMcXzjprSnnzaBWBhbU3hm+pV6D
u7aW0jdNWoyAsgcLCS22Q26MQzjqp/xtbDquEVT4w4WB3oo+H1YwVDqbcZgzbkZ2T0OZVvaSgDKe
jFmQaTB69yeUTCMIMC8PbTfzpvbyzyKcxBuekY7x990Gm1y5lx8qd3NfdlxCOF23sJ0gM6Rj5LE0
7aBiLCulvn8REpWc/0FUY+XZq+StmYtoYLyqLh4vFePBu3KDW2KOMIvQY2dqNe08jxNnqPDC1/Ph
+iRfHzJhItZSXOy/79FGw95AW098RMbRNtEZzwbKocyJrJY5I2iogm1tvD2UQMD8Bwsr30tAUnHg
nU18SjHOJ2dxmUEmhLV+0iPgw1s1ItKsbublfqbY0vwY3tDofJCl31MgtUI7AlDTEueHsA6lm3X2
bVIYN68P9x4gcTbBu9zmA+Ekw6kH5Uvt/cS5xrc7qP1gfoJtBJN4gqmkLyXXfjOYIA8Ws/86bDAX
e7yZWX5tSjuyrMomOkUE1orC5tsweBA6jsYsKMcgDb7OG3jY3VunfNAo9Ra6c8tijTszJkX2nG/k
fjDl3K87TgjyT3lnerHDrwt/BtHmmJW98xgQWkfli4dnVTyzAKYmtk0Kt8VUagA7hWGfzeTkq5OI
6jjncwPftFtn2fkgjIbCJd+c6f8+lgM445KBcJcy9oKhoSHhjNLFivza9eaacNjd04LtvHKis9dq
xXXMndpkLbbXa8QfDFqns0cMZWIFI+ebm1+5HAd99yah9/LCyOqLxZXu8wyN9HPAfoxYklWkbnDA
n/VdcUr4MEUBLvnrU2r2ieJ/ta0e2KkRTggljf55sJepN85z5LUN/nPeNi48pcrMjyr+FSW95EmF
Tb5NZ09xRPQOak6p/7OCR3O0Nv2OSAg71qHZxBv5um1gWvJ0+EzbbOwG6NzpOQzK/2n7JCdQrrAi
ocjRosUsxFD51GL8o6UWDlFzPrMvzCzrfZn+O5L8vrWmdtX8cE6BwIXldDIKx/jqIX53ludh2OeA
rv+4RVPccAjRYuqjf0dBB8y91wU8Dt2dSMcLtlZsbPYAgTmryEvI2eg31YFfYz6OXWzVy2BhAvHt
4izdG1Ocwlts9u6CzUX2H62ZWkyQWmPmvURO7BQfhDf+2hOFd+pLFZoCpnC5y80k5ZTJbU16rIdP
YF94JtkjCBfzAB4bBYCgBsDv/OllZ1ImlOkJKzf8j85VpuO/LiY204BUDtlGmWxaR53vOeO6Ct+j
j7e/CtwOutgaq8r/bVPvicNwJn8Vc2r5FpqQj5ZALf2gfyp+U/1O5ZuL+4dUSFZQV29WhFf9fCP/
9fyRYGIvNJKW9UnK7gb5KvkCzF1XLsCnNltZ8Pvz47viE19yudfySeqQp16MD6I3YQZLCzU93D0n
Fw9W5VyyuaqF8jtUyuegkXmfR2HWjCPi1BCUPBYpUx7HZqfQQ39jS2CpOGk9w4ZYiu/mXDMcSaXc
bllRvOURZV/aP8JkWMhMCfDP2+Lbzu+2SOHjr48SQoFn0Jwhvwdjz306VXpCZPPhBtwMDSxs2ooQ
+6IMZo28vb/Xceyu5GJ4eO4hFoRCtZ+hClt4k2fF/b12ARL8y8SxCB32A9CxK++qIXPnBrFhjjqO
R+jUWgYZAyD5a1+gDcc5z/Rc2Tca6E0qNKPDGY9KKhYfiQbnjaqfl7SM/EognCHx1JNuFdm4vpx2
hnbfrXkBdqMzIIXlTuv5vWVMm3L4T8fSg42Ky/r+lCQyECsDBS2ZfdJEqMyatWcDfunTRYt6nfgK
r4NoeFFH3UZzPdgiRUvAt7kXeJM4CvoxEIROVyN5hc4xin9fvYi1ElukX2zA+s/mdXC/fpzVeUXe
tKO8Exmypx4zLDi0iL861xSJmFlHFaJje/DYq7KNXXjrArFZ3tL22SyC03dVp79fqWS2Dt7z0iVP
yZTD8Cb/hqPiadjacRhozVsQepAxGl/krC6Dm/yPAoOwTqsNMvybPIsRoGJJFoq/6JPHqpvZvclZ
J8JAzbDFAOcz4QmekTY+tbpKrtU0H0eI7pxy+P0KtukDU1h5Mw4IPe0CiRmB1PeeH9imLOGsFRr3
jrDeV4/m2TqO3jKd/DEHh9J7eoEX7W2BCqMsmFVD6hbZJg0vdcZgmjOnKthfSBZHIWZfqj7D1SIr
Hsg1z/ESJCm2AuB3XB7mahMbDXp2qzIc0dC193a0KF4/EVn/1fTJxIuGRwzccNOFhs3ZLTDLUQ6l
6UlRaEUYEiNBCK9dznUdpjKDRhMK+TmQv0JPTJz2kkzJmYHBWXeFy8cAGpJ3Qf2N5d1QwyNvwMmO
KCsyPKPOk1Uu81WvQBLuL4cvXyGRBfQ0+L46tjBF6Nkah9wLwUkm0clHo7ved5Mm3KJJIOCAza86
WNMXeCciOkm/xXm9IjYr63gYyx+T3QRQkFAlLRW0EEF536exEqJScX9KsltWKiAAJ6nTpV9HqrkM
ldGzb3PIVWw86hNXVohpmvp1w+EtlAwqlYUQHOOp9ocEt7OObHp5MNHZ5t1lVEqvwF5A2aldqTGi
dtDVYgJWWwt7aI7SV6n2f6+kQGYEvi1YFHOo2+4KyGHzmYbPahKDmafICoz3RJppgMaw2wC05QQG
60pSpMb3P2bzQ2p30a5v2FPTAUIYkdNTWyu3lTX2isiokTDm5ZzqU0cS3tsaXmTjD/vRgh9s2tLZ
zB5+uFKC7VAOiYBuLzu7F7wdT9c5zoBdf85l6BM8h8BBm6jf9AajMCQJ7XCx4p6oso7nghYBlGId
IaBHWC2WkBVgDiP1LR1nrTI2RC+axuPCEOcdRb6r+vTQtq+XFMFh3p/Ar72HwNeCoYhBMH6k4xMV
1WbYu9Q9xBtq1/FPwEpCyw27RSWlI6lbk1Ha6kcUncqqrEwo+EXVsuc7Z3QSXNl0ty0S1K5L4YgH
pKois291Zg48QnrVGy4Z2B4DTpAI/08zVYaJboD+XeqT+jwRxkdd5YIwnFGmqjXACjgRyktm5hyw
bkvNKtghz+AzGFLTKraocC4l6ybZ0Xc5u+41j8wc3UO80fKvrtG0jeG6nIf9jHnQhD7IJzAsb0QJ
Dssp0EyT14OtZ0mvzth8/O/Uo95z4OJzCiiRn5YbD3sSjJ6wftmWwv2rweR3msmoQB3PlK2jEy2V
ONAv6JrMzcs26TCbJ6G+diBF4wdG1/FxLHPMzNTjUC63s7IoggS13gmU1BGeR0jAJ3ZDb4T79bKt
oAkKcAEe12RWEQT72fzKbEeDQatbyBXCa+2ILYm92r8uifMzrM7Yk1pkR2kPuLhT1CMuo108P6Yc
SWQzrbMWZeonyjWHcTE+Y8jp9k1EqDQpv40ty5yXGK42H4gD7TNyeVYLPdTn3kBLzw/bEfO1uI+s
fh1O4GCsdGgM8B7Si5bo0YQQLzDeSExLQOHvANigobv/fnnQlkvtaMjHwjNFWTRZdbb/gPLZ8Vva
P/CR4Bk9GgWApvstL6rs+GSzGbW75v+P6MhR6jkdIC/5M1SWV8WAXUtYddsL2IUU/AEE/jmUhxso
AshnnpF/Z4RNTBuPt8ghyzz8xyGCijL70Xfo5D1zf9468VmZDQGP18FxQ6R7OQloTUHDHCfdnzsK
3B8z+h+kUl5PmddNNLyyC587zR+vpsJajPUUVtglTCzGnwp+hcKIczYiJ+vIxvX5dkSV+JjolFVk
eHzjg9dn5XwpHqOaYGl/J/hPlNIA3ziMjOC4QUsIg6aJnXOZg6HSvAYzVPB4P5rL1ZS30yFzYO9e
ALrk8jwvtSH1HhGbwABqM2mdG1KQVY4hP4NvIZm9vXHxZ5vTIxKdDMQOY6AFu3PQD4bPcY+VKSk5
+6DRK6OmeQ6hLCkGguzAjtWo0ehmnigut7c8VUE6CVg+tQoY3RnbFEd3DYSGXnFR2oCHFSabTaQ5
z9sQmN3VFMzgr78SRBHNDajlh/ijkszGGfppOKx02AgNwvKex/Eo/4uW4gUFZrSgWXQ8rJRNoHWr
aP+FLr3xhQ4oAweyr3d1u/hrgPTmp9qSDyNNveszCwbLtk6Dn9BhCzvsx9wYcbA4nvQnvRLL6Ojq
rhX1tMJ9ewHTPBFKouVXvhm2+j83gK8NNRio9v1li2rncPVpsYkvCByYyEBGOlST1IRq04OrS7XH
B5LWkak0N9MKljHbMe/TtdmE8EwzOL7fkHT9coCQTw9t53btSsjkjNgkLtu3jMspcEJ6D40oLnkB
8WUWes55ACcppFuU9AJ6tsdH2rEucWsso88A7CMSn9duzBr3pYFVGxOGKyx7ElcmRi555fcIcRZT
hFflyAJvuIKgXjsYo4ml71vUmBEMFAPH67cnE4oylt6dNdXinKkt9LF4nkmK/8x5j3Cqp1qmstbj
KwTCUybFLxVI4u/XnzF6be8J4R+TEz+ZTA9NP4joDIpxcnnYmYPMb0gnwXomEKO8mN0pspJ6YRRa
I86bgMjaIdassQ3/G/WEuyQie8zjgLqX1ZhAdWlY0R3k+x+0Xs/wNIBnyhs/r94TxkwzlKSlj+F2
rrsmLXxzyhka5xwZIT9LSDD1vP4wkfNIJGMAXAMXHEr5SmsSQME4pE9RfjwfNgxzZA6nzNM35VRt
G3M5zWu2TO5Q0l+VG/lcObbqQPRecDPsvvJYT3Kx112RSI8bHlagraf32dM5UBXyVvEg0YFvEfhB
f1Vz2BGXJI5Qmw/WOM5Rn7Z/HLPK/FS5FOJ8iGOSylidsoNPWo9DGCMOYU2Yyg+XLDpgV9PU7lEk
H7tp5fm5pasW1c1XkTFtCGWfiyvy/YuRz+XejoqYmKpfmYYPirWmJSkUsO5ipYj157LBeJtYumLm
FdoFiaKNuakgTXH02YsqsgGZwcRyFnQ88shZjSLB0AqUrLMRJHNcNHkUWfwcZpmXmk86s0Zi1eVa
bUSPtwPrKyxxJrJ0HOaabd95lDPXTiSuZkxgZVCXWTpqo5c4HMcez3B5VAcswieuM1TVh/FUOzab
E4cmggdVybkbPIZ8QHM9PQ4NnkmrQu+y+vvQ6FQgdJzKMkfJFY/QpOrIn9a4vOlsCuGUAw5W/Nxt
Rl2DSFeo92ORoo+OH6sYrZyKquA//msExbgt4tjUh1teEa1+uaKlwdZWF15FgN3WZfERmjqIbxs2
m367cLewbAqPloUXMnMdKobfvmmTXd9VaOB6tuAeTpcRWVfzXqINXfpUYVxe3A93zhvkXyYZjAI9
GrKtqVN0rstMw+BUFhIxmPd7aFjqJrlF7a/ObHWon3TE+BAAwGYLVbOhpex3LJx3lv5l/SD55dWy
wWTFxDJrdYpiNyfeyeyGTnqeCrnw1dlVLob1z3L2m4iTILypbuBtJMb5raIpAjE1yw2LneNgKVeO
I0Xb7Gc5QTXwbmSRZ7o6rjEd//w4LyNwlrHmMCeFHFHZCDItixM9rBO3z8L8GAjdHZalQTFM09db
iQwEHTjHZp5xiDS20YiK5PxF/F6IqAvrwZ2EqbpEzuoTPof1Kb9Md+EqirMXIu1soSZEaFhxVnPG
3QXB6uKucm4UFMM0SHMjHT6OhRZws/ExydOrzaKV4JBzOMR+tqkZGpo3lcYx/pAOgNxTzQs5looq
9kyLDii/pFW9u87FxycqCXyTquaw+mar2IZrEUofXVHd61Sth0g52qtnhXg6m7ILKbl9gGT0QAZV
nB8rZG1hvu3LVnIBR0R/IcejZ55P8+a33e8vVjqb8g6aLulQJyzpHonmHfgIus84QOf/Lg1N4/Vj
LoMEhkNgs2TaOlB1dHJe1XAfVJ8MO5PT+ClrCNSFJH6JK6tnDEdVpObexYxPToc7vJ1EGRhYXta8
0Ht02EQWtatRoo1B9Azxz9Wvf9P45x41/xEuDUTkw2EcnYTfB7lNjoM8nW1hSfUd7jaEjVVCmsL6
gCiUizGx4AhmtwMKNc8c4qaNGZt3ykkM5ho9fTRZr+0oybMdGyCoSE4Uqvm5LugQDP641xOdUq6T
vztnJDvGG2stqMzHmuu231F3nGnOSGXJmJWY2dceT5KF8/wjR4Qa0xFCWr1NDUtyaOvMVa0Kc6mf
DSkjzphyyPT5QQzTfKXN1Mb8H/6Se4PPItKG8RDLvRGToSlg5LX7yim8V5ix/oWT24j6tAaiE1ER
w/l9XA7qXBbWbs+zLVAuOj8mFlf+ZyWm/3+qT+hHKg4JuzZRcCnr5Uz28hpxhoVUT5UNkPUBl1qM
+ULf/X7h+JACnI+bIE81cfgIq78wNMn89nlaLVE7ZOreekZDFTyhZc6EVCnfjiJF+/Lbbw4u0nXV
GwOmisJYVew2E6nWv9dx1drpanGzyLJ8HYSLJhQt+1jL3G3bniBipzXbZBbett5fGi8QA7lXc3l1
MRDQSgketcw/mn9ryG93GRu9sIUzWG0Yb8QzcIZWfdQBTubhPs6gJ750K4/hHH338T0bsAB4UX/j
hnZ331wHmu+M3LRtIl7ukGrB+GWRGVKqsnAuaeUG/f7GtPVZrYrdm8CMEIk7YLULQ3qAwNWlrBEV
dDNTCo1RIbG1WAhPyoK4vV7NARWhLHbrA0KgXLunxMRSqoUDNkfe6aE3AC4OrTmIsk/Vwj3i+/WG
fhgqnT3y3uEEgaybb6mvmcVFPyXRyuAMF76NZhNygkVzz/9kIdUdSOEl8w7ueH5vGS3GiueyBJFk
f/jZmS6B3RorcazMxo/FMez2rV6xQdhpDcSjs/AqPEklb61soc+q7nB3Vz7lW2W46ZUclbWtUo2K
d6vdFfleVhT/2VDT661jplkD1qEeC6LungOUCL5pDJOSZW/2Uov49zDiJL+6G6o8nZCZjZxh3tDu
yPJ6rbDbCq9KTZceGD5neB86ZPNty7dbvai+hQ8UJfQTdbpUOz5gHERtYc+zc8sRU1vf/cAjzpQX
CF7oyqcD/v++V8fGA+92nVZi/OPNiDFRqiTmt7UJNFQuf3Kn0JDFyFoooss5xb76D7sp10EWjli7
BY1wEPLhXNuAQiH7onLPwtAUf/hpuPtU4glzsGkuKCucIiB9d7q+rW1wUAhNug6mPszyEyWDEAhU
Ug8h93Bw63u1HvhpPtH1svDpWf6XrmaGMq4sqyrUkxEmBFpyAhi7kIUfTMCVyKT4Xa3d9+PIOE+S
UIENazF1FJyao1iNiX5fG+CW62JgXyvGGpArKWQELlotfKczJ/PwzXtfIyNidQO29dqDPAq1X9e3
KqvrHjKrtGnryBzBTSDHkj65RIKJ3QeX/F0vN2+FvrtR6fiw21LbA+/mOaaHjmp5I2Ud20pZYe7H
B70IFLnFTPD3IVdouU3Di5kOSa44BGaIoHc764co75382p9jnQilkw/Ufotc5wowqpEN/CrFeU7M
59GJp5ni2yYcQ/ZSlLxN7auKAQ1x14+A8O15NETR+ATDiGG9FNfl+R/QOR4ymfb3XbzW/bM7/cv4
WhaXwnF03PHtZtoqsWbpQ0EIq1YT+MHKl2qjdbc99cIjSLyjzWeYtlKHNcAr6hcHisJDiLQa+lKl
LA8JdSRKMdtjDxqzpri/onU/chn3OzU6JB/7yjrVF9qBQIp2+LuATcE85PM0gK3n/4yofJwkvixH
oG5vGj4Ovpkjl5klLp4G5mssA72UCzqQH98yQfos60tGxPfWR0Qye1dk0/XVJD7gs2ifPOff3VLJ
NVUzFJ6FQl2ZG6VLf9cG219nMFSVFrSfCQYmiCgMV5HDqRcnOdY8duI4Bcnz7HdNVCYGu3/8PD/B
GkUHt/OkOFr3/fPV1opvF97oYdpsEtm19K23/MYVCf0PwRrCye21EjD8Drsr2tUjDO0jXSrXfYad
EMuxuPSHO6Mv8eCTNMu+1qXunhqTnWC2lOSmBfYF0QMcm58UDdjixIkgsCwRGmstV5ea31119ldh
sWj4isRfhjVxNc0G7zGVx/fpIUmbykoDLEY+uYIHZLR2vQ9Hs4yjZIPs/2M2pJamNu30l95SWqg6
7Dv5gmWyTw4UhwPnVEEr7wZi31q0pk8NhTuGrYtQZpADemFEINkHGov0WhaTwFHWnR6G3xLs8DZZ
ZMKQO3LHInb+nFp7zkKRldFGzDxosICml3BGkFRcTAL9Y+4amFR45KtkoarUFqdthU5qFxf0tb3m
dpNjCOII7cdSiqBGH5Q6bc6QquRc94wR2Enmps/5s4Ch48Ld7nat1WiaO+QlPEORS/nuf7ygnvvh
Lxu0M7vmhwFWJlMr87HCIvscsQwREARpR+zm708i7ux+5fumhJvZw8CB5a1oOnvPw5Z4ZejjnjUS
JU+oWA0wBZW4Z77hlPzy3PwyAge2xML/oZgsMY5NTVqN1HUicHfQRPVdgsbkJi5NTcx+R8MmXD35
hYd5ManR8zOwG/Gol0RSOQj51FUVCgQBrmp3cqMy12lSPVYHuTmCUsE3BJqyQCHgstoSXA+FQdSw
srkVMFXXv7gMotrgsV5rQPFcO10GIIkS+4XnmreSPZgTw5SvJlUJF7Xq1lMfuHCf6dhB410xNhkd
/IWzc9DVb3/6kEnJWnMlWqG8HnED69n9hCxodbkjcAti27Ylh4g8umiqWfRCFXkXPfoXa/gExwwy
sZb/OdEfoQXCoYY7IW6STNEHM1FC3q1xi0xZb9wlsILcYmborijeIDOagixOa1VAV2ZdFoDiBvC7
KIXmJ4IjeFfg9AWyZ6Bi9nLslG3ItyoVlOQYQd2jN09qURV4rD6XSxxDXgKCQKq07cjW5feo5ylY
Gn447eT9toM7BLKhm1S2zdTgKTYlRxqt3H3gImCeJgFJjOsZerl0k8Pk5DhpajvEIbmeb/VxeWNB
ZA/ztLbr8h3RPyKddORbv5/W7DPAEEKuu/Gnld+9A6VPTiSKxLsjhLL3uBvZVeLiSUNKTCl1dOTk
AZQs7VAMxVPsbgNNK40O/y+c+i9fidfZyEVJiPecGIrYKfm3hUQQ+qTSLlceeudGr029FKK/eOoU
RpeEoXzwEfu4zHruv1nISu3g8oIKud1RZVsu3wrN0LyeyJx3psVRBuUZ1E46EtV254bFbc8uEGzD
czOGBiYp0NTuhkdkveeN3uqRBQ10Q6zVB6wH0Gz8tiSseo7tXVn6Noh/Iv9OyiSErn6VuojD2aJE
MEXFIzqN6VJ460zcBOaUbwazXLMWYUpn5XZSOALaaLUHf+vVjwF85n4wrLxx+J31t0G0U3LddR+7
imYwzcPRYYuFDfFyyJ/32McWTLcRndrlSOVvgEqzJV69wnyaKsDKPV3VJqExu8+QLGbAzfgrAmis
9ri3B0nw1BWhtG1N9jy3M1M+KL9uPD9EFlOE8sZytXdlvWxewNePImfBqdoViyNpSJ+zHiLs5yL9
qKXCGUEdP6hh/DM09aOMlwXpe736XYHrZVFJsFI+SwBdKC4Im4oRsiG0JTQYJez4FexqgjmVMwRw
tlWZiQ2qhJyDSU/KX0YbrybnJD1DiB7/u5AO0fKBLUFNcsrefnQCnNbO/KmRaaeZigZvWY/K6RPD
wMkcsVD1lf7OMVmG3PbiFy5e14kpEjad8tFyWcl4GtSC3zN6pWkthWtcR30I4aZy59QiQTnyR+bb
XKWu6zSq96abxXHBlGz0g2fb5cFEL2BW3dDBH+dInxq6hKLrMUtEmVIyyFhosy1mJhkzQb8/f7xq
79oW+w14TgyJrx5/stKAVmL2ncZIpk1hhevOh6L08EZVcBTGkvI2pCoqHt04him15yoHzZydy755
eTJD0UhTSkPpv9CBYbmXBI0D3X23gbsx0MW+eCTM286iOa4TdLI0X0DDJEAluIqPLeXTg+gsy4V3
Ou3UWHStlE600u/R9wfoN2lwNy0mrZdr1bxMmbMyTE2g23hcdycGrKvSEpEWM+2JRHF/1JlhKiis
DCA39PL80s91Px6tc7I8cUmUKdKjG8NApPOhxlZIFg5O9OKYxt4zg2uj1nmUjI7KHKl2FkGjHH3U
qVgfqJcS2EQ2+eE9Vu0+4lOQbHcXIUtZXoRBKu1CHjMJVcSi9pWfmQC2Et9Er6cSm4FVdI0/6J38
x1RmbdcTXBnjjyWQQDw+Wy8Zj/gyo2VqOWOcRMglfAPzRI4BmvFM+7bAILmlu7IOBV6UiNOCqKzU
3Rn+PgtrWvQZeEmJWJHiYrIFBmoK3p9hq/G6UFpA5EJmTvKy23hBPMgIm+ZvmQc5z5sGLp2q7WzV
6VJA+QUT852QWoJ9ieq42adtob+fmYYvGSOcLQRI/6Xuktiu/r4yqQoxmckBCvtvIqBHti/hZKM5
zbzFrPFud3BF4La+kgMTx+UwmV553Gtiyc8g5a31GvsK7wrhCPf3Cz0886Qy7TRk1R4hsCiNY57s
V+40spvYAfHQMR6h4Y52ls/N+XCkq58Wu5kS+e9+Xx3sPsQXHC93yTGnHJCymY9fD3rw7X22kgCm
+bpFvDW9p0IS9Vqma/e8GuVeYHbwqVnDFl+V0JkCtnPhqEDfcbPjOzGZDnsLh/qEd8tvtQbZbXuo
nSPbfMAH4JV7Rb91j6CrFrulxIlnR4DFJXjrDqoUtw/+kECKwUm5J7COJV3F+oirvHmMOMxqJsjc
7B6H3w/Bd0JaT5ZtwgwCYEygVbtBBW5KkvOYxzhQqWmNw/Fd4/9Ve05PODfebjSpH84DWwokO7Cs
QQIq3GaiC5Vqw6cNCuzX1Yij9i6s61nkGtuz5QzONIcgm7Ioon2F6rgVWdYi92lOaJteWz561C5A
rXDC4sVfPBxow9IN/X9FlgV1DQk2QBezMCAEphZ/z26ROQKnO85/bfaQ958DjvObEKXdQiyyVRBG
6OwRdpiKBcbC5r/uqNF2KQyphGMFMXw5Yf/yrp4isx9Hc9g9HkYQspSjfiQca/GREyHDI5FuFLJe
dI4Ue/VzmbzKh8GB6ZEmwmBXkz2SCfJsqiUvWs6peyOu08LkUWPd/AjnVygMjDYyJvQVgBdjdr0m
WvXbphjiGL9dvKDFRv/4Xn3i5RiBNdH0ZfrZ2v6A6CbW1oy9nTtyltabKIKH6Mj84WkHzXJ0VUjj
CMxysbWb8UJ1Ue+9C/jzkN+BgN/sPJvLQpTOR/uoBU+dEOcmoTRr55ZCucrYvY4ZMN8prJ1h3De+
/4zBKwK+XnVyCoiFTbplFf2NM+JZdejNZfeSV3cvhsGGxfDSZYlC7pRTCbSVkV91assh2SZznaFN
Oy9loGookqzNn1SCqbvKyy37cIh46VYzh8sptvAzUgKI7HEHTt85nblID1KGqv0CmuWo7XPZpUB6
CMXGY2UDcfFTSs1Rs2a0Imh1ZBq4yXz89cqKUp5lA3pQb9kwsT1uIWiqAUIt2huXr6q4DF220sAX
jJjgX/Dc9Ye2gEOWe2DqJD3zSA6A64+2w0k5Nbxf6P7yrsHwhUh/WQHyPoHqLd1cKB+TsYJabR9n
gRTyVDHJZd53R3uryMz6pHR8YfimOt5lYf7kulyQzJFNL3Vn7DblFdSQAymD+jkYT5DwXquLzQlI
7H1BiQcARybd4iZ2LMxhkep2EMv/QBTeb9IjvSDJWX1c27SeVTrsxSkjRxy5JIqBnD3fjjy0klD5
2kjPPXjB4u9PtEyLxri0nHkl+jVwbZF13+9m+WAeRo4j6RMt4kWQS5MkjKsFoVDezfwf/A4x+PGY
SqXPC9Xak1VGXrdFBmWnj90QlDtjr2QTptCJSO3O52ZZXePFg0LlRak0NqCf9hAhlXrW77hJx4oe
Agt9cATQcBhxgsfKNi8VhHcSzRno18G9bfeviipT67jiRFCVD9mehbBZGTp4eKfNxYNEaq22p8k8
IEcISP6dAIKpU1f4H9ZpqrGa7pAm10LMAqTxCgdZ8l1IRKEahgUBuAEhMxWcE/ZOc7UDSIR2P3F3
NGuyUJtTXYs78e9+efFXebOcLL81OeUBJAwlVzd2QVIwNz2gkNOLiIaw5pbWOAxU1mECVDiuVaGR
/S3I3HlK956ssQidUr/SRK3OY6nvD3ODDKrP/lkkrYhIavXX73RyTxncA7wpyPQxOJwxLJ4hWMld
oIKxQMPIbrZI9YP8aL1KcOergolqgw5RcH3f/4HSQ0kL8VazS9xhT+F/wCSh5QGU8QlS/FVFkGR9
WFOMkwTdnQjE0W0wRNYL4M20F+toab7aCR/kGlqSXwj3GfmC2ydqTGsB7y072CyntyPVf6SymZKl
Hxyg+oN9xmLycy79JqsfWyP5LbMglEPsvj+KXkiiAnDiCaAPJBSvklTkPWbcXBk7TaZcEx2lDvhP
vWgUQzewxb5jZlqGJxls5ePAYfNemnvhuI5crr/rqBzyo+TtMZHFUSCacAAKA4WCBtuM7cg/BEsX
2k++YYZ4Utjm1mt6DiqQEwjLWIFApbaXOc6nR7Qh/5ldzMMpUYx4K4WpeQS3MqvvySaRlC8LI792
zBMknNj/Kj9gP5WIKjIF5GGuscKm/oINdbUzw02CzOS2Zielyd6ak6SiV7xgsQkJL6EdoaGkGDJK
lW/gPIhDfXjk4vWHnVHV6BnVdLuv+PWuh7PsiMHbsc+vK6Qq2OjZfeOnO1pzlz4xUQjRtV4Hvouv
TqUTm31va60btDTGsJzAzL6ZGUZKyHwr7RWyHvVw0v4gFz1WEMSn03V8JbPWjy7BCRoeKyR+WjxR
Qyr+AHtwR86U7ryOZhPTrlVo49YG2q15RWKHxY1mV43HQgikNV3EmIU/bNV/RnS6Qr5D6ohoZwGo
avKvdRzyqtykjFqI1QFxs7BM1JzwF82qNqX3bIWkS7la0vZrYj6vzjQNSx6c1HTYfhck3nuL2Ftx
Udvx3eugajuLMLRTn29fT7bDV54veqbSnp/dHpIoCqCPY17/QYEGGVWijo4hxGUCgj8Tp+lsCgLq
KZyLfA/R4mYQug5XWmoYNXN9uyfxKLPKIAvf9wP4vBI2kNc+muiqN4OxWnjUUNxzY5x/DTZIc07m
F1eEBPBem219B0t0gxa6fa1kfEyxf7dYkCuNfduvgGCRewh3vdissSMc7uuQghnOlSgR+j7tXzpa
0EhzCMbNHg1jee075lJzzxgI4mRlIuJdGWPCF6xkr7vygiPu+EjeBBdEUCLVKXBsYkIxchxS5eQJ
UqHXNvd3cZHPxwTQQM1NXAEFoRc3+7CPc1epnSwqmj3ocbmwFB2OBoPhDdXp/c64okpnh/9/7qTO
5PSt1WuubVA2ld4rlnSybuLSXprTKuAXJQKGhGbfUIFaP8QjktZLtdGQbYCYyx7TdO+tCJ1rP5BN
5FgcpPTmuYrUdwws0yx6ql1SMpgUWRqF6X87lCfhk223P7p4DXcXCQaqHQx4ihAIDgjsLPG4SuI6
ZXOirTHUkf8XqCRceVGJxn1wWitHTJ0vW7F2nS3zGsY8kYqEBOiJPTd8jZjONHRlp2LOgxwI7660
ZtFBMcj1GHydrx5QpfJMuTvUB+iEe9tQWvFQu2pn3ZgsjLh1aIYShvASIHDHzU72Ed4+sJX/osvk
kiIL5Iax/38WjurPByESVCYhT/vA7NQGx6ztppPbO42UO03mL4MojHCZT6XKTJCLE0vRrd8cqO7R
IVkPnsBXWRFjjiPWH8ljSFWhayuQNw4FmM8dLh5vJ6fljByMEeWSVxVIfcxxPEONR96VJOUz7xnp
5/6O7w/hHJccsABH606sEw3EO3TZlo4skO/8aB9599GhFNbqvqNUzAc41b1rOopBDdt9ac+Akyfe
8CvomqRMuo6Yv+eTYP3ab7O3Emsai8/MurCfxVE0SUyxLso5sSF1oVYT4P+3j3xZ0yYP6tyqVAlV
ikT+/aI5FNsew6/hLAvqDwmrNdY3W75Bwrzkenw83nlDHDeOI5yb2uKyyk/KPuHopCVXChoVFTk5
oGO0J5OAYjuSqm4p/6BX6gTw9EtuEKQPwpNf1iQdGdHm6QqHgl396ZSM7JqLI7fTz6IHyXnbRVmS
LgxfXQ+rWatoGRu7zLMcIBN3DVbSmFkbnXHY7mkgGaX75eQoNgXNxWhZG5ROud0XSEwfLP1fixQd
hpZCFj4NJToMaFzM5a/cjgw/xgT+QVhf+KvD6BCYVzaBZb9z2/pWo+fLXPGrVpTe/GLimRYHnLjM
e9/aLvFS4b7fr5neDXxPtZuE3zcL3QPMN+f1ukha/F/yu4kvZ15lnppVDHnkd2qQYqS55CFVxpyA
2+V/m7rogaIgaV9XgcyHmziLD40hGHcJTMYhO93KY9eG7kPa0UC5Ujf8Wa9J4TriUWAbeQ8NZLJf
cn/i9ivwLUp8mcWYs19PFV6RQr5dGcOHH5fXAhr/m8L492iu4tKubjTcQSOko8Q6R+cZPm/VVYY1
lvyZ98ruukb+V/Pmn1eibNG49s7uvmWhzadQy0PqLZXUqOSwZYz4EpNRXZEvymb+XWgZCzJA6Vel
gBF2t9ssoB4aoYOJ0Skg0eJnL5ZtRbEUM/oXIAwyx2s3LMfOVzjPowuAWBSu+Vo9Lg3VkOp+il78
7JHU2D3L+N7ZLtj46RJm5eTrTfipSYNCPrZN4ylULHMyK5TGWLwNJ9ZWjmMSBOYYjrpZOK7OmXzh
ekRNPtcGh3opgpGP8VKkPk097OVMN8uze8w+iRcQzxTElBHZlArImDq3OScwhgW/PhlnNh4iG3gu
zW3Lf595nJzBUI09buyd0khGTL08i85T5JQG2dAFL+hbxmqrj84+BfxOyBHlWrh7Ra3xWkCRufLg
qZJj97L0GG0OJ5LKlDPH5LnMMsr0t/VGMR5onc0SShtDLQGpRBRLgfyfcRvq+9JGtRMEv7P9YcHX
rh6VElpiHq81uWAzXY7VJusBBWzeRZ+VoQMVhK4mUTL5foU3yCt/VkGpi4Lgw7CDodau+yuoJZZx
BkseK7pkc9m27w9Z6Yv4PqBF5kMa7A+PzwrvTEQvQvRshDcVjFmopE1VuFtUdD/R/+29lers0g61
gs5xTXdxIaqGlVT0Rc+w2gEdYp1vpADS6Hoo9FSFDNqRpL1GokTgS87D1XRMzul2pJjNCAczVZP0
yeEKF1TdAsheS072zCS4Az3zbHVDubDeFytwHJqttMDbq9FiWqPn9qyVb3VEajFP3mCOktIJ5V+F
f/EUuLA5LTRqxjyXgUJtYhExVurRLEPLL53QIpGMhm+CPlZlL5EfYOEVRoZktc2sAdv1DncWz+Fa
RrNwPeXM/P0eNlW+C4GBotShzNbHMByRZZnmxP7oe80t8ZOWqHv3aAR5Rb/Xha/qwhUckSfRQmD3
128MpXuiExPccLNTHVopY4kAMl4GXQxv2FOo1RJJ04prKe7k7evjFyhawKN4gqkgVTpIgRfenmti
Ib5FRf2CisGu/xS7jmAdKD2o98yGnV211feXcbAIf++HUIFvF2NdKUmVvleOiEzXpRRjEv5GlD8K
VPuRDCVL7wdKY+U6KxabhogMTn4La1jLv6BwlpoNS060MC432Pmw+v1N5F8HvEQqC7qNkKcblpNx
PqX5GDxzokZ2r6vYIByPFJfl/VGt9Ko5bYYktf+XZO7gVmxUcfEUWm6V889W1sBqVkpCwEHQqD25
sPuTTqktYmwjtuxmLWrgoSBbHQzRCUhFn8Vq8yz/Nj7AFavY4uXa+yAJKyiKJyB/Vp4d0ZKTlZOS
h+TWCE23c2LVcZGP4n9IgZTB9OgU6StH/1zMVSFw2SPXXCcUbVg0itIjmbtVhP2qPdVoifwiI7DJ
4wnq5lvLJ4XDEXf0BBrFJnoxFPSvss+mgHSuKf4oAbF0iqacBV0h7wkUKGOo4JWPHku5WqJBvw9B
T3xNwAIJH8T7/zYD0dbYNUag3nlGzrj5zb3F7+hdy/Lvv3NQnQUgTGCacXcza5y40NTsJkK0OzqG
uPd6I+kg4WacvIGjWVRkiO23DEpetvpdpWyd07Oxu19U2mjEoKYLJfyvdKyQo3f6VlhgrKyKoVWM
6tiSCM6S6h3sjQAc3g4IUO1uIZdbD8NHa7fH9uYUjd3QFjvk9ehZ1i1DQDx5JuGExH+m3ROWZqOD
Ny6ZgVc/D0sgRLaJWW9GFKGm05hhBWZsfs+NbV+WM6xZX7dlC9NDMnWAOL8T3azkovZ3Iw6sIzFQ
YP+S2h6F/1sLe6tXS6pAC5PX3zDkOKnR9lRqLMFd9LoJKeXVe1NC2osHh0IgkrVi7CegoWJq/3eM
1hcxrRq5EwiEVvwzxidP3sppeOt1mhJGIV8OJF3QSpeHwNDY+Lw1Gt1UbWrwHAQy3khP8RzZ+ZtY
GQ1sbMhVAMTb4E0KtpySrVUwsMTeq/fagb3qMGvBaQzsvYfW3P1p2JrvAfeTFdx+vGh0YcizEWWZ
yLyzuTHO2J/VQNVA/ZqWZ5oknQrlHqF3cr2HqEvR1dJbfuGEc8T/6Ywhg+vMsXUMQ3onaLYA00Iv
iQerkMkvit3NM3AEIZtboJ0kfJj+8hHE3W8QIOQVNKh2pBhfP9W6pd8j+CbZ4OSrdvx1yNqoZc+Q
/4fK71zI9mXCES7BIhJII8tR7AkbDcZCN+f651Q0hIe2k8mmVJYw0rwCD4T5mmc+1kraQfL2r7/+
KeNLUR+PlnwzKa7l4KItacef/u59s3O8FATCifDvMMkjmW8dICXR7o88EgTvdTmF7g4DmzYS8feB
eQHOqM2QdMZ0xp+BmVwDkPIMVDuy7J9q6/ed5jpEsKGT/JSNcmVbXIlmlSWhJ93rIYlN5gwrNRjo
aDKPd4KWacmhzm75HD7NARNquxSVUjQ1MPNoPlTDyLCKz3c4W3h5RCfK7aY0IBDnyN5AeLM2j9vO
A4CD61tE24xWeMKeB497p7dfvIgf3FNb38NhXT54jv4Mpeky8RmWeWa3ayOLkj2dIwbKeOwxlymb
RUV4a6FII+vBXL+xUGmbFOcRdlBWfHhqqA9UFb0bqiUtKcomyxjWFVN66fq2uDwheothiFF4l8Gn
n7izAajlNIjn9/Mn9+G3yAoGy3ycHglDadql7uzcJIvoEaPMDJ7IhQByEddOnTRS/4549yGqG1XA
NdepFYzUJsHGJEfnmJNQSlqDau+iaGNE2biAYfKy0vT9SR/6fLMP+iOlp4TgHO0RE9nRFtKAh7ww
NQiSu5QSaLBegblr7ZA+xOma8ThYjeE9GxLmlsQiRnAahSRNV2iPBS8cWPJt07gqOSw/1kHX+0tT
OtuhVIjy0xMLOT0lQWxay1DS1qeZWxjK5S9zeHvjfTNJT8I6KqlEKvNuKTJ7YonXpjGox6ogG4RS
vubCyxtejIQNJXUFdj6iAj5qEaoRDMYCHwgx++WmsP2Ldh0JvSgJ3IwjVEtf9k35zTmetsv8kWXn
JLxxgb8cFkaW9QNAbNushMN6dRZpbn1o61hYVCD4bPp5btMjNDlFDbgfRZq6WB8eJYof50/0mbft
Qp10SjbHRDoWNAlG03pwq0tYw4nR6mPNF710BYK414NKG7L5HevnWMUqXMeSGWnW5NMRWT/AUJPQ
UkRQPRyU5Y4MovAb6Du2ICTdY/47EgG0xXMSz05vl8fgL2ZSqK46OXUW6rlDfspGiCRFUblTs/QI
Hp0/B9VGoEYX8aOcb8p0qpH1NbP8FKD42NCNDtD9OTX3XtiHPo/n2wnGQmX/NvIQuYrur3XE7KML
IFbNao/sRNXRFsPu4gI11hPh79C/q+kGktkWr9VMiFti+BCgnAJ93923fR3Ghw1bm2+k3MIzjtZp
o/43tirhFFfcVKOVRaTfrzEcIB4aHmNF4AB6u+4KmRxN/s4dILqWIlXJVYSLFV49mNQQFbTVxwhN
DokTdAtnPZfzLFfm0rAkuJjeDkDVr5Y/XgAsfMonchQd5I7B8UUXJsaPt8KbEF+KS6NNZRKZ7+q2
J92DvWibJwmVxroiCVib6qBw/l0cDHNBn5hL0dtUAVGFyk2jqd860SMZLp/YsieNLEkno8vdTTvq
HUHn8e5ybxoQ5zYWq/3ss2QmPzFqFMgRyeYJLiUGWa/FZNfAzLYnQXNQ8sIrqq3y6F5KoiqHF1aL
4ldp7ic5XkNfpYKkfmDLZX8LmN1RDSnInwKJHQTRq5uUCFRQVx/WeZncWqzcW57rzD4hu4DvPSG9
z6E/TISS5kPrkvx2yYFZtx7fuG//yt2kFVEIXL4wq/65SmkQtmJ490FQGYhUkgRv4kjRRBiSnS5I
rEOv7KhLVRdpfhm5J8QZwEr0XHjt65cAWSTK/L1rFmFt7ViyQs4O45GeV8pPWhdaI2F2+mjBkd03
iPzlpoxdk95r0D6YgVzqcyK5YMnh300ky8PdnDuYho5VrKkTPWoEjt1GloOpXl0KWq38f6xDfZ/t
89S8Cse2XY+pdUAT4cqeqWjBc6KTC+icW5OqaaPB30IqejeCTyY1ksWG4g4K8mADn1E+G4nWLbp/
blfSMvx3aU/CuVAtP3IxC1x1yQkfh87VoYSfSOXBV49UiPmcx+X995A0Znksxd3STIeT3dtg6C/h
tKp5V1zXobqSAapmF1Ee+Q1v0Dfhbd/cMpc2+p6fuebSRYUxC0wvKZHPA5G9rX9gGprFnfMZU0Er
ACQTaAQIhRtlfmB+7n0t5s9bamI7sjT4IGyeDdo+jdDlvqDD95pY0sNMHpZrH0t7G7iGV+zC+K0T
RX0SLdgsP4bvX5brPHBK25F0BIJCq05pONckYTGZDLp/3XlJRoYov6tHhBcZN8X8cySUxn1x1THV
dq7NPxCdgS98IxT8FXkNo7W+bdD45oaA12PnEMZn7VcI3dNuhIdBoCUbm+0mHCM6ilwo/mSPgL4r
0fZZ0nvAULMErsPImWQSrGZVZoYn7HaDNKJbB3CcIbCNdjZpG5NzouhmH5UBlmR7tTy0OJ37vq6X
1SpQQPqxSYYfleEIhjgO0uOFriaZYHkCopzFyWS/Jx3UoDByNm3lyBDV05XSTz2PNcGSHiSUF3r1
HeiNmXZa0vZKnRDGg6/DgjMWQxvVxgbiRaeFWaPlu6TxlOaPAaG+bE1aX7qIMF3KgUVUoyg5iG93
uHSLWQT2xXI93tCdWGGJV9EG0J3njE+JF3TMKG4I6ZNZ4wW66skLexA62fNvnj22XmkEA6raJN+7
Q95yuqJ0ckwOmHiSC8DBsrMbidBH6v8ysgBrj4V063Ve870B+BfSaZc1aPj1e4KCUW4YFzBRxQZQ
IWWyRtMBrNP/e0MjAjAM0tavxSXwobwXfiQbCCUFif9Eba10MtkrCRUXSShBdAyQ+LxtTIOVCOaD
gLZVbsauPCvyBRGN7mb+221txu3u17er1XN2Vd7q+g3kSd3Jy7YgJbrw9nZ+fT8rFn4DEsPtBytB
zz+Z7DfjQu+jvCcCsQma/as8P33o+SzXlf3bmP1vLVe6ygL4/W+uCrTsNIBvzjMkl4B7w2RdbDmK
MkFoQFB5c0+dKvQ3i04s2gUMkfcUsmlYpf429qti1540Cz7JDVrlw/j/L3cghjtvHj3tvfs4NST1
Mkz0TqL+BUg2UZ9BNrsFituufe9petP2fYKQ4vTCO1xs6nJq4CgsAj5g0VrD/ZKk0jkKBBUuSnsg
j29sfehs+mFunPwty5eDI6dxwQizsGYj7AWTGjyhBnVWLMxd6wgQnNnNH8fGvwZc8DGLu75M/jDx
wNhSl9//jGdVL1aPD2SHgOdAiE8ndjfJZ059w4wpplOh1Q5w2i+64XvnxAVXpSYoghsPkmC9ZUhF
o9qEvWDEZKmZuZ4R0qTESVarUA1nIXW6UpV2ZbPYe8MUJH3VI3oi6vIAut2D2Wy+QvVhOSVZlewt
WHPw37cvoidMEZ5pekR2Rim3NFNsVHBw0QtGoBWtg/LPhptYj8Xt7KiRC1zPiYXK4IR/AP53UtyB
m8N8PxN/nVlbnhfZvrBZgYInXgjObBvSogroh3zD8xCHgnT+SWzV4YmK5sMtn+2sdC2UjYdjGEN6
w1omCVfsRN/++UHpjNT7JpLDZBg3M/f85c7rkepJ8j7A+uD+Z8AzH2pZz9Qwnj46jTdN4c2fJOVg
KvjYWLFKtLKlDfyKgDSwCj+x2laiCQc1XPxHTQ9pf9xUXDR1Tb4d3yRHFz20RADaAwct+aGMErW4
yFW5PF7CoFKpjTb+VRuEVkA0K0gwctKuAkmQRzUhQ16P7ybna8yZSx3EsX/gXQXITmw3cgupKJ4D
avDwNj4AatQ625AwaQYy7B8nSbJM3i9WTju7jfax61wmRQhtCrx2qrID23pEZGwDBROU6wLykikQ
0dE7FpP/eGkMA75GpIaswGH8ZbOl7SCOQ2nkP7I83527eXeMrF5OQgbVkp75siugQ+QFMInkguS8
qdu6RVkN8Qj5C3Ss8L1WjgmubZzmrDMcspFhWQ8xPc6fKGKnS6TUv7m9l/sXaQ9m//pQankdAUnv
UibgzjbhdTsnLxX4BRcSj1iMQgM9VhFw+xarmHgb9GAThD4z9o55ThT9K+Xc4MmLo0cgr+WFDfiT
2cQZQ78WQ+IJVdrFa+BxvDMXG5RrCcoHbhNvH5JFlWbMMhDNLbgswSTdZ3ihgG6FumKPaYvFKjeJ
Ryd0opMp5J0e3rNYW2U4MsbT5O939SP2RAf6e09r5OaS7XaZ9Tu7wMPoU5i/FPKFf6FoD1aRSs/9
1IQFpXkTYX9R6JvTdze8modJo4Ypx6xjMS6SHgf4U1+d/vurIWsFetfVY1dbRz+tt/cUsakVrNZ+
eStj1IAbEY9kApIbIPyE5+twG9RY7sP/lh7QZdLiW+ZJ6cA9/hR0z2vAU95aFiYs+XFSZ/Rem0Z7
/TH+omJZRfTUdqGMFw5Lo7GLmuWfh674rR5P9Y6LJSLhxqZ75UI6xJc7AfAG4+O5jATsP0InwDSe
DnbZ0nU+iw+8h46ZRQBvWmi/VXQCrNjkWlJaizihJoE4AYeiSn8rDqdh/BWNl3wvnlxU77QNjjf5
HGEnsOLNzxqDhexxzrZBTuHCjRaiQY09krKdfLpEm66QNQ3YyLc621aqeDnqHDqT+l94o7piEykZ
kLKbiLaWAb7JaXc74TIwN2QWduBtV8Kqsh43yZyxbnNbkzrlH04QaJRcBE3skF0xvlNew4fD+PYn
OrlHPONpbqEKtF45R+HEye849Lwj4ZIAn1hfUGku/6HmShpiLlA/siwip1clKAPBPkyCY8qcwPe2
dvf2O+pB3YhrfLG80aRidajydzQ8jZO9yOnwFeqDQ8F8sPpG2vQGdDOD2fEOM7FiladE6EqztC6i
vmUYDqzj8sBXCrqvSch49QOrHEdnxE4HctUb2Z+qI8YRYfZSJ2EA6yAd4QP2rFmJTYyXvdpaDgxO
64/NR++BFu1ZoOyZMLiHgHqqT62j8iPkkqzZgoCX/VGQqJUAfph9rWLPtOBYoiSX/LyJo0YamGvX
PUcVaOH2pIplE9PFJagquNZcsUYG3cv4905ruuHUMZSEKGV70sq4nVRY5PYnIMJQFUFebl0zrdA5
T+xvQB4IVzZP9W1uqobwKqEg03Z6rtSNVRKCoZfLNGqCgiZU00iGl/8mx0Shy9lsmtPn5C1wZuZ/
GillicDILp/GA2GFiKy1EMUEyBqlmDvL69LwwAwyuPT8Gd5Pt/yesY6xzlt138UwZfL0OltGKGSr
e9F+i7MiyLOhHxZW3NPhJmA60K36EZ7jIZprWo+IFDjTchqhmIrE4cO6iy13McJ8UswGV2UCRE+T
dMP5faUeo4Q2XdO90jX+Db6i96iUieIjkZUTY331vkM0BnrVIbzEve052T3ucmUuanyGlNyqHE4Z
6SvxIg9SBtVhxGhCw54Zzi4S5HPN6Kd7ch3M1ny17bDJVNHkY4IfVKALtXGi53Wd9joLl6i9Sr8m
ESw368G9y9EdGqNcQayNWTVXAMb8bgEt9Ownbfp2P7mSDitJIRmtp4zBBoItSpmVHUUlatl+e9v2
oY974ooPhizSFSTs2WhPWRnYGpIP+8hpfDrUZ/+8Je7g5NU6VpZss6hlwPLjmxbHTaaOvROR0boE
Xu5DkNhSIa7SkV8aASvF4/xtS7L/E8TpJbXMvMDnDGLNPDeD9mC/TulLqKcZbXMk718alesTTq3V
eOAWoOCtILPfq2l1u3OIeDHty/L4rB4GQtCF7R8TjNfDThn483h0mcNlNKDq5jODCBHGv1tQISlf
py2/IRqhZW1nKzzZzDWJGIV1Gc+AbyZx7iz6MxpuxJPMMBULx6JApCHASLFmwRZB3c+BM0pvFC5D
7i8mPu0JDQj391v4FuVmwKAGDtiMRN0Alj/zkeEI3zzHQwyVjVTbusp5vYTlDkDstATsX1+bc61m
CH7egoAKxyzQxIbTL6gWrsAiygqgEyAZ/BYVldzamDmfWDiXYo8KPWddhAK1m5hqlmGNVV+YjMeh
ZjAuEdy631zq8Lb5hOuctpMxsnNAhwb1I65jrPvJneiLHvOS/JJZVQUCBZmQ2P8shZ+iEYtTURg9
eOVDf6utSQJM7+HhZSEO3ABcbIi/PsEuYHq6XK9O4VEJhRQ81sXlGhYYUZMncbM7LmgLLhGbORWZ
OkRQG+2rIaGAf+qsQ6f3Y6YwW12JD/nSJqISHZ+/mgmzuDjSXuwLCc8EF4fF3jKTgqmdDmTp+l23
SwTw7NKNwvCYPpouJa+XHjJ3m8dyWPUHv5AyIH187kHt8zgjAp0NHnmoqCXLTttkgTmPUOMf2Roc
Hn1QoBs19JlAltkT3Sb3zMOhHa6f+oqDa+xl/NAP9CceLAnGDN4Q7WeImVvgbIoobMa3mm2nNwdo
UgOE3fCO2KCmRFP5m5rMtyNtUXz2hj8R8cNCLbQLMnoHTnZ+K/izLuew88gEGoDSKJqjdYAIVsxk
FnZLsjbC3aOKjF+ICtYv3+SkzHc4eXPcKJgVElLq16O40VLVqOUtax/HUfKDO2qkDBUF9n2sdfIl
+GW4mAHcNTdqgDGdmOtGCTclTlfr9wEjbqWV3bdwjl15xIQ+8+RoNapog6O8tnvai4c/JS0Yhykv
Cj5RzuvNaBFd3YO5lV3nhH249YSlPnDZP+2Z7z00J7Tt6D2dFCeCOF/TeOKWRlTooqG6SgL8n5R3
H64AroQ9MuonOIDPVujr2ofiH2iuJjqSWDocWNXzMzL95G9RTm9aogD4ywcY2LpdQbaGbFpGzN15
DgBzAp1OT0ZYSX1Phtj/R3FnyX4BdFiWtTWtg1HyupMSeV5+T4ieFMcZvWiQ8nfFJ81Pu9SMhWP4
sdWnfap2Jp+D1Fi3hzHnlpcu0kBTAHuefjbcBPLoWRDH/raD42H9cFB14U+C9WhGqn2LK9FmPzII
7OiylVPnvnSm3W0lVAadv3kVgPRdcENVTkM6KnyFxZ1d0fbCRpSz5VYWEHxRJBfkYXLENK9JMyJO
yHxPLPGJF3b50G5a6UY+6cRJa3zDBlGTja9Wt9hOn6skg9VDDMmupZYguPRPPQF94ThL4TArhpHh
sHSL+i9d9GYKUtr+N1w/V8rBdCsMTpY7dd+js+uC2TSyOjVN1k2OGJJ6vF+jwB+9J51a/p4ga43u
im7TdDdG0k2nakK60/i46IY3NsW+A0ya3HgnURA63i5I3EN7CNe9k8ukwEim46WaAPDgxemLKGb/
tN9qqx0+2+6cnpHwgx2SPixhZPeo7+igp8cHh1oC/I8LD4GP6I9XojLsU4de4FYyTO9nrz2JPf7M
kyvqmoBgZHBI08Ip2xK6od14NSODLtE24idAPTaqZwdRCddemWTzkxM+Iqm+8cKbx2thP4+EH/au
Aq/KR7pgkKofFf4tCqJR78z6ZcZ/jDFu2StY1jzDXI1BKgOZ/aK6SAt63M7DZbg3pN1wpwq5Ldfq
9qnEMAAczLvUNqQsvPMRw63Zywk1e+zUn7OrvHoJpEicnryxyGQLx4dhUZmpcFs+d5Rcj6IxblzB
mcH9CGmkJ7Y/WLVsQrv5z4C2TDOLSG881jLTY59Vhq4zBy9V0OLxeHORjn2sD7pVTqKc6lTGn45W
80jBDcgU5BaPFwhgWfs+OUBePXKAQW6KbIbtMzlmBST3BDBQlFgCVypI3mtndbI8dSMD9kvEMlwO
HoE0l/EA0ukHCVwtJ62NCWHStnzefw8MmgyTVV4bOk6uBN/zTQN0mxSsW5E+bC88KHvYzgc2PzQR
kTBRG7Nr7YuEp4U2HmPBNm+PlLWazL4vQlYo5dGL4f1lzODystPoxnZmXpG3+Iq9Xf8b/BflAMiH
TmUzdh25sQGAZa9mntpiQ2E+364LvCsPAgEcSKNwGQ16l2PxBjTsexxeSe9EXSjzikgWUWus6tSq
jfEEY+AVqcpipUMD2lYkrXdtri+mCgo/zA5XFRvW23O1GotDo7u5qWZmWtpY9UDm2vvSnhEUfz4s
WRbKl+BZlo511pIL6jWbl5WSvM8NbYM9PniIAjhOVwjbI2GsX+M/2sQ2ul7J7gy7nNy4UHozHjlb
l1W2zaxvj/YOyTyXID8DcVw0s4YDTjKevb59jZCRKpCaQzVVQdFaWoapGIoE+If9reELHzhnI4QV
l3lQEOOxJtqaVdd9tTF7kW7y6cvaAUpEvoV5BNHUt6HimzzIB4Ll2kvod1rRTGmgu7RdJu/S9Deb
c6fldeNI0T/W5C7OQv7BnZOvmJX7qetWFXRiW0GoBT3atLItexPK8MqDkxyMdP6+ml7shpcDQrEA
IutCFgvHtWXZV6gbfOdnElz/LYlS3mgr1iS2uQe3VM7crfidFvuHUaVD8rXwQs/NBkxrqnvgF6po
pIizvsAB63ZilcE9Aooix018fbQ20fW1fAnQl7A38HBOwygqz2KyYCs9SN6gPakKPbmiAbriYTqa
15PIEyLgsAyjIyufauCMOUXxRaCUidJQc1pTSigj8k+EsH3d9xn3XdjVRH835ms+wVPEOZpumNrG
YeP3EtcLw/xP9ymwwmb39rxl4RUQSiQSteDZV42m000lry6KX+J9HX1WbL532JuF3z2iib4aGLKw
+Jer/m9oHJFJBKLRJtYApLazqQAUWMwIJf4HORS2hicoiCSKtF2JQH2OxwKZ+PO4iWXmBNle/kNl
vlmui80JkmAKyTQdQofdh0HQKE5QYP2D+u8r0AIpF67f1PZYVFuz/o44qr6n+ulYX8o4idYHIPma
jwPFC1lHvuEtDrFKC+7c8u1XHPJftOJLUhRdxaG7DWbUHFtuqxhgtUXEhmRQUAxKQFE1EvwkLetg
BpkSMkMqUwyTTMVcHTANaHUCVaOUBKb5d33zMlOIBnCk7TWjHBixi/M/SCcrQ87e4U4OiWPG/EbJ
PbIcYdy8iwfSKeic0pCCYXs8PFGsSFfHt8Y4MfiBjGv/sQIuLXbAeoMuOpiBvz6lEvQaMIJxo0Uf
3EQd/IyoQ340XB4V26MI18e/7PjE2OF0BcQoyuecfqdzstDmbKGfqnfHjwIMYP1lRIu9zJjj3S/2
aVQA6Vlxo6qGL711pfBl5t8VENiU+RomIt/pgwO//eQ95TTesyzW0NR7FnUOEWLHVm7CXWtGq0lu
1UDP1GM9E2BRzLmZ2YGCqQm+KxYyf/0xP5i3zoUOBAo6JF0HXA45eN/kHz/x7xWnyqI8XwtJVHGX
SSm5ecb9vEKn5sAQHi953EkForlHMzU9kvIev3OJuSESmWthQ2GRfkrCgiwVjCzNu5syCkWXyOjr
2Qt8KCvz5FfgJtJ0y/p0ykbujxp5akqA0UCo2+loxzLPahqtt3y+Z1GNC83o+xg7jpjBMMtdH/BX
1D0D0mQHqv455FZJniZ/imyL2/rNlH3J0Ys4JMwZ0LSPNaoA9fdTcRpJRQf1OZbUU/q/hL/LroYX
RLR+O+qboeGDYaQeKKOaDZx1BCZ2nEdVL2H/llOuwwi2O7djLy2mzB3cdjKzwGEW3vejk+BP43Bj
xrE+laLO/lBZ7RHjo+bUp0VFEjHBHNdTynDP5Er7U1tCMwCharhhNcW3exu9IBwFLn+WtTh+Oy8e
0t0RjOmJzO3/NE8Sy7ecuEPHPX5SiEn7No2OxArg8OLjhvyUNk1zsXpULky9NOM8m5LRqBb6Eamy
txKMObbyRTQq9vUAT4nWWn85x7q4q3esoPsTU9l+S0HzQEnG017fo1q6o2POALGQY4fFVYkB8AEJ
BQnZZBKhkia4/pEVjfuag33H5IY1a7ReyAifJLWQqx0iDBiIgzqCClC/DWpgAbanX7vUGoLBG4Le
iF4EHEOFuin/a9xor9rFUUJfD4vBWAo4JRky9V6J++5d90Cv77rOkTQnlzfqsIjeY4LDYjZFhvsW
j3XMsbpdR68sX0X3a49ljxto7Otu1hPyQF9aCgBHUzz38LZ5HaeUqIm0U+ScpO5SQz/XJFRWioq/
HET6ZmQ44CXstMpDhVXiK8ioiG9TPg330yJ74+GCfOEgm7tKopmCqNuR01VKJY6nQqeVFi/72//X
OuBOYRXop1yb5iGDxuRxqNagg8AyTyglPrTNPEwpWq2qmAAiGufElKbnC+d6uZ3gR2N9NY4+mvPy
cgepp83jozyX8sg71ysorW/1Ms9sTyQgq+KuezgX5vux6gRXQQGbpUc19VREvbPA+CW2yIiIv23Z
mpjjJkk8BFed8qyMJRuQqLJUyN+FYVEvJbejgEHqgP+M/dqzK7rWcFReSR8J5SWk1L5FHl7v/m6K
B4dGK/nmmic+41ZPGjH6Ia3oS5C9VaIUh8bLAnWEwwLR+s/p7aczSYhSrcEMLNMHxg+khkR1bN2I
cWSl+4LRbMODzbA8SMGwXnKMpZboHXN72Ejd6lGKChSSpDLD6KE1hXH91xy2Zhz8H0Liao18Y0Ak
xXBAvCUIZSG3y0CL7mPYm3u/RWg7YtJ7zO+RDHypS0DnKxjAmkkcBvnnXwmXQzE5t8Ws99hVKTLD
npPE8QPeZeDkrQv7laYunucy2djNHgki9CtLsp71uTBF2E+ufuBz7OktDg4CQ79ROp9e/Vfih2HC
bUUjBng7StnE7/y/pv0eUI0sSB0pscAs5W03KHOFJMz7IbZze0drd54JW/TfOpDa62kHw3RKKzoK
A+59b9Unog3Jay+Ma/RepUekp/mu5VGqN84pxU9dWAY+9xLKd1O0NuYZooibxez+LPc/YWyzsODr
y7fbEnK95Jlxc0PRlt9Bl7WpF64L0ZS3ALLqsgAu6mDX28XYLr4WwXaIBq0aRltjeORsHgoCn3mP
dfP2uutgSHYjx1z3gsXCLc/28wusBIyK2/r+yDci7YMSNG4MhSztIEIMOqY/xokfZjxVsXO3V9R/
v3Pe1Phq9tCfxvzbtw2nUsnbgxHtIEgUWAL0zUs+iCyvYm31lGPC0NbhMCXG6qQbPWOmTz/F/Rb6
O6M9KtjRYBgXl2MLDA4MUScHKx4EVk/l5ZgvpryotXODDpBkViPl2L5DnxJDBjX0xvHRZ1XIn/jL
0gOrAN9PS0WYOJuue9rGjXCjfGNMdprUOgaZMMItF1islYF9itMxhbcMZwtxCIsqelFLsZx708wW
XyLY99g9g3x+vkSxmYtQDCyPKbkcCR/Gtge5PQWb1ucovsbJYD/7J/+h0kEGfX7Fg/aZ24PbRQcE
g4zTDWywy/mE0TUhQBsyAdY6AgcjvaXjDz0AkIKMgk279AmxVww+D70wJf6Ikp/E1Jw/z6YeJLMz
J+jOCFH8G9GdmcADXPpYyFnbJbpn8oB4Dw414hwKHHi1DRcgjadkXSN1fyVkq6QwzweK+gJSzuMm
E5PRIeaoG58mNRV++rQSQ25IfTGqBj+fgd/P1iVOdMWa/EYLbbmys5r88THxWrXCPgcgGIeu2ZGA
SrRhQ6/T46nnvViZGB8gnUYWsh3aI8onG3PRndkdugDQdiramf4VpOD+uYNcHNsspP1v9quwc4Du
cflV2gd9Sb2+GkRkFWLAR+I6JLl3U2H+AGzrzBv2jBUfg5mAzRxZWGkEQHBw+sPyxgD6uJ8UchRu
xtGqbh4aQfNC/wFWm99HimYYij21Em2TLDPHqQQOC5w+SnzNOHTJC/YFBxlXpnJCC1xnEprkUezs
klreFWxOu1Nr5VPUxLjtS9leQOAEBeh7uENJbgG9UiKysRxQZfvwtHy7m9OEnyd35nXlMy1IkTGk
HmaUEZqByVyzmSx2tau8iZ7+U59YZVhrxuQWhlUlKm000NMT57gsKCrE9Chj0+wjrL6K6XcRy69k
TMyJO7vwgtGIrmMuylibpf4vFjDh2qifK9437YS5IvF7cs9VpAlRl4Ui+lD3tCehVE8ttZnN6rZY
wKN+9axNkVwoEgk4PpCn89wsKYPWcAoF7yMAL+sZTTYmFP2D0tpdn1jLrx+aQNluDEOH+5qBkzJo
fgpoK/0fJzKDGqW7gPx4vEbIdgIUXTIR56Be7aNTwugzCxnzfsQVDQXr5TrW1tGI6y+b7JAOtJmH
2NvQlsvjIkoS1/fXUOCF8HKAPOu7p5E6MvlXplZBmI/ac87pE30x5FbzV6ssjJelCP/5R8bt/cxN
MEuuODFdVmnILktIrO5gxxLtFcAgK8D9svxctywcD9OpubonIv1zo4p0xF5Lpmf9y2Mylf/dk9Ub
1XVgHBN+QHL4aPqoFnWMf+zk14ir7VPoBaiHM/m5Oeyc3/YLB++T1Zg7murdJfvs+36VFaLsFSEz
e+/K9DjnhX7Qjb8ryirlX5ORbgTUz86jMdV4IOhqHMM+AhqhGd25jL4tZCxB5buKoT5AkYdRdsga
HHd1rmCRU8f2P34pmq2N4GhyvbD8DML8lhLL5/TDlAO7Mg14Ylmr9DPzdC2Ux90bCHTxAZzxmqf5
863dN4AV6cI8wjmHISPT/KtHhydRZr7ypMG1hj/0Pa3vOAq66lT2P+hgsi5Mq8PQ8BcYVc/wcV2t
t6/yjaytCC171yh3PWXwjSXg32CV2Rv9jIqB1a3yqncuKiAstNiADpTQYy8Lm/UpU5pj0GxcUzEk
XxixaiuVyXCKtfkDBDqvPoXncbw23zPTHjoZUBmA5yhX7jGMNhF+NuL+Kiyz78qQvV0L23UEsxt+
DsGFmi0wh0Cfolv1H35wpI3p1ch5P40VQZOL0aCFG66VNPN2cJZqruv8ym3FBNlvjpVQ//a/Hvir
h/w9heOYHs8EvwB9JLmFI8q7kILeuAQalnN08OgEff7l4yRj2qEOwWsgYgA/4Gkzs5/dqqk/OwJl
B7jYGbpsfTZUrkGb2/wE9lPqTj76vjetGp155yNbUh/9ufEA80ZE9HafurdPecvawTORDJbNlqTi
yN3Uu1b7NTW2DcqbQHt5LqfVwNC1Ax3S//We/cWpBNvvQwnvQqVO8tX3QP45ZIPN7IVOdMQxGRZx
Yv64mKuLdcwpom8h0V3i6blwb62OnadbJYlDr33K9rOjZ8Qvsa+udCGvJZ3zG8NW3YqvdP+j1mrj
5u723dnbT6ZsLZxNY+xzs5qLV9o9tBJAsepJtBF2SMTV46v+/il0Q4fLod2cWbWZ6ClB2vEaKVKo
7CaBqL+lxzt0hVESqDdLlOPowmVI4Z1HHyK4FBoI7fJF4VsN4PKJUR848QViWsYzOoCdMo115Ekg
ECRzbVj02efDHprMoY7MVQCdI2gDr+s+/l+XYrAv+E7Y+LwmYs6iLQT5ae9odNOtGc78fZnD9Juh
1L+sVYhBlkNsvaOT0mLdiiXfaNpygz9xx8xf28pHPPPgNXysEsktQvf9n+2fSp39N4ReGjcCpEFy
5rS9OTqVWzprqiErdAzQ/cHcmBbXptWyFYhLu9VDIqWY1ZZzsih2pzzCa569OxALxl9U1HXjT9QQ
ku/RTquCCkgOn9EjWB6673KENiF04WwedMUGKMqcTafr2uFgMIxP6GJndiKkr0MzgyuQpP2jkeMi
MxxbSahEoQN9rDJK6Wx5Vkx6qBbUM53RSAyTXd9245wUW9w6HB5iDu/kbvMmB5+GXpTiWoRmmfPE
gqn7dusN3PQjFnr97KGkyHrC3upkgTm8Tt0g7fXEwBGD3wCf4eXtpJwKwaOnrOAh6aKY8GOzHYcb
eEAqgj5cmbWyOIOTIR8dIfo5/qJfzAXvglaAonPuCaD5cqZmxutus3EEl2chnc4rMawaAqZbyLA1
+Ga5dzCKSbV4RAiZDK1nzI3S26CYwSpEMGchg7jqE1TcAzy6WKuecwHrQ1KEj541RF3lnvWI4y9T
uFEBULFZWrmeWTSt7k3RZRZRL1LFJtwkIKwf1r4YnbgCqFQZK5rVd4wIoRRNVQhrzp4Jtd9OM1bW
UdR3f7JwxR2HfpbGD73kP6l1CD7pTzBJzw6q5P7iqcze9u/pRNsiL6GYf4ghcW2wma8CugdR4adw
ZJQMxwH+G4C5c8fPzK/iLTcUmqdPFPJH64MyN7zW+/B4lFNVevT8k5G/C5TBySE/AGLp9McydBRM
FXkB7bFs/FgFIfn+6E3IJ7F/IYnQsGXtiXlATOhjNU0LNWM7KJApor340RNL62YjU01Ik0LbWNRM
MDpPQBAhg5Ves1NI3EKWRqGk2P9S5fkYsGIKhV/ZRLqLwJcc5m3s7d1EKFnL2Bv2aXjit7wH2MUL
BffoCKn5S8D8zw/y4YVpDaQf/v1Hkj0du0Ko0qevGTyWZbT5YnNxf03EpPSzEc5WUSp1K/DuVLu4
2MRZ1tc8e+cAK67v/MEgtikxtnslHI0ouxcAdV1TV45+V+JXXmLMPL+9E4avEFl8t+PhAooC+84f
+fz+9q+9EnnKaNmqfQ1nV0ox5CQUzeyw6a/E8exI7cQoo+yz9JWu8WT0JmCXrWGqCL4SCyviMMbi
TVydioig2671FYJm7jjbDohttHytzBI/SeQFBitZ79ena6yGDZjqag3pPIKshCLE9yQ2dugf9fLu
g9M2+xbmeW+4Ny3rgd7Gr+mCfAZZDVxHE4NC2NpwzNTRrddLOXFe7LpnLUgQIgHD4Ge4W7/OQXcg
l+RoofVHq3sqXM2RDWetKEGjc4WMvr+F3/fwYzYsRFwoeU+G15886nuTFKJpM0zPlrLioWJvF50m
pcfl/C0IhfJ1PYqzSv/GFUTwMD9n39lyfRWyb+VpqlwahgRKcO+BzpRrGV6nZwPhnMYtQrusc2X1
7QEBn16d2zfL2W7KtGgJxXleamSakCI3tGC4gbO+ogjyi865Pjuy3tEpyeEG85rK22UjIMaksa6q
Pi9kMTxrHrwjBuV9FjY2oT8eaetubo5ICRR2NWob2IqUx4P3SPs4AIHcWCXP7syGCNjPcSSNTADv
sT/VT6ngSC50VuaCK28EFdnXwJ+wDs1kJLxLLx7ztgSZQmVCU+fDreBWK7x4BqFOVynrdii31Xyu
odgSarwqDphryYi60lptynDeRPkKmqg+qb7NKFXtMbxb56HohO64fRFCs6o18y7jocqKlzP7v6xL
khlP55WhSXbwHRbAVx8Khhc+oZ6AsKDV5lePhk6Sr7S6guoGAmlOI9EMYvbocgcJmbJras+g/Slz
tTilyVYA+FN0LNDH9RPvTEsb0X82aDTkGVRgxDn71HDayJ8rERz1NB8lYRkiXQkC6XQSS2DJMJC4
Gp+CIUlYdYzoTy1lai8sEVTpewpmZzPMzKLIJwwpow2nojYbXVuPD2rc7Z6CogXdti3MzSFFIWad
qS8lJ7qtPDC9jhJptgQVLLA3pHx+3BqhjRDj8upDOqI6rI9wIruJH+ueDeUOjryizfv2tsJXNFqu
/srimXlK4U66dD1bN/zbKW6FmIxWg9v/FEsMOfrFWv9qIvZPsr2DLnEFXFsVwnyNlhpNO3nAN2Qr
AuZA/stklLWBePcqBQ5XX5N5I68iLYcRMUoeHsKRVIpwf1HLLKwVuJGgvYyvw6r39MrWVqYjfb87
XPIq8gkLOalfdRVCG59R62CKlsECOrYWd38/qzCpAnaWk4pNwbuVHcbXmnjqhowT/J1MBlfv/2Py
a1PBROEkrN183n7HtqVYmIcJeACt28nMkOxNxMzgyb4bAhkPQ+Dh4RLE6dnaRGdeLeXJ/CAzn1Z5
MCznDQQClwadgqbRIIT8lmz7YuWl0ws2fF00WwaLBgSY6ZZKxiCBVEQ4hyUajqU4OCbLv/FZSQBg
xGrvK7QJ4NXnb/UJG2nQHNfv0IEWbcSQbp201NYQHYEinJHsilO/ojc4XSu8fTuUx2a29aB7hgf9
Q8JhxFDuN1Emntb0fYF15lSuKY6Ek7xfY2g5sRIrDSrueGvQSBJfM3ul6dvpLtCURxOCNes65nNB
8pf56NNvkJ8itLck5mZZIr4Z1fuPdwVpgZpVoKXoynMybroM+o8MsUOVqJBWlCPYGk5f5sg2rCCJ
1aX72wsxmvMR2IHI7nO1I03mha87y0aGJunimfnaLhotui2rALkodM0pqMvXUJtLz7sNX+gNM9oX
rxTmfiZZf28wLy8qr2qyAOCXJ/eaC5c+rqHKFg2U37fN25BLBgsbLvIFywFa4Nf2CfRQjg3UHxFN
f77Mdk2tOTqZxRGD7qvNdQElOYbsuwrawmV6tUpgDaoBuZ/gM4em1we7rEmnPSB7GN4XP7u57YxF
Fs0S4ybXkGk7FajSyoVeQ5iBciXiaYPX2CfkTNW4ODh46UloZCUILdpPd+E8qYneZSrjjnxbPYHI
Tvch/ELD0DAe+XEyNRmD6JglFQa4fNOSdO2XaKgp6/D7RBPsvXOrJUptdGriYcw+T2aaMXrm0Qx/
AgKEDZApQ8XiVfEcUpwK1CuRpkxO/gbmm77J/BbYVvdNIyMKuuI47a/qK8rMMs7rcF3BIE/CNW1L
Cl15RbKMtWGJgnpSyu2fy6VUFTmhCHjKvZHPf7oRYyxjOIxctOVPYs6DsAs7Tr4ZPMLe6K2ouyjd
sU1gaYv7CD6JpeyJFzcX0gUvAKG0U3RmmHdvR+oqPEV7C3ci8Of1TjIXJKMl5x0VW5L80iAmHH7i
JepmhxYXeI66PHHQsHIMNDrd5Ogydy2THrF9q75IWJyiqcr+AArmAaESPssNkMIHvtmhV1Y2wzYx
KacW4goUeMkxHbU6E8vnrr9fSGKoNTsiSfK5yLp3p4gkSSFgsKohzURqFEbslIU8r2SXYZBjAk7M
MOVXGGhGOS0KJBahhY3KAtI263yiofXAiJjIOvKHjpL6QzpA0gcMKQ99QMMrCiVUL5jKdPv/Ci6T
QJ5tm8JTVz+XavKU0d8isBrKS8zzgPBMr7Rd6/7ScfuFgKTkcDOlsWjR4QmuLIDw/h1+gz8Jc3fe
UXhO5zAwrxXaxfqaor6pTg3VXb7eYwW6/zSKeoEy3NmuEHXSV/8fI0DNZOQtd1LYywWjMgh+NYzb
nwwZDJXbUF6pQn7tY0RgjYPUkdRlzvqwN8PA3HLSd4kBSPHMFTJ3faSM0lbhWqci3EEhJU7Wnwgv
gCFX0F7x3qiT7T2+4HShFlkA7GHGoC7Z4BoLawzcW/vK5PEvCk11oWvTIrgWDLUdntRDTSHSuAhw
rmrtg578+Dwmjomy99sQDxe83/vIMKPbx2Cu7GKghwT5OJ1kwAGbqonuy7pFkjug72a+8QRwFFyb
UDs9XmXENF7EF+Pr3NFkB81qW+s3X8Il83pH4rNvBf6hyWFf811kySFTLVjEv95E3A7msS/B4LBN
1n5hfb6gY2Q3jofKmNsOUYq+02wg8B+9P2uuO5zAWcI07FFutGGiXz8OIIXLcDEjdyb5myFL1hll
RT+NKmUOrjktPPDAwyhfvpH1pGcWUOVXppjg+prVHkG/yI8eWZKQLKsCFCIe5BpLvPziv7Om/x3l
AXuMHqPJHRztu8nI0Gnek30Qc6KqeqJrOzImbpuwvWG+20RqMce2RlgVilCcOaKsrSYNg8E+tFme
QhJvXOEbv70Aztvj3NdKESSgEwfbsMFa80Jdhi7/LhyF1GOLNXOi6xG1zTNMpsNGw32KJ9hugrLV
HuWzB9sEiScj0VL2wKNfEKm+rmaTqtm6aWKTL5kR0H+PZGOLmL4ajqrUBs/CAJ1NKPju7fnG67jh
bv2w6dRWlX/2sKDza6iVPMnhqBbOf2zzTV76n7AjXtp6GM+2mSi5HPcroHiGoo08zIZ1E+lIK5n0
H3g11Ql6H6nHdkpsl9XJZnoH2OsIQ2v0ShJFy/79g5fvhnCTs9cmHms/3aLjNDAnYJy1uk2IfKFi
EjxRihRco5BrhVoq+xwdl/0FLZk61QPR1pZ/YUXiAAcydmdiS61RSK24xONjTbCqp6oaJNfTTAMR
Wldwlr0lRWjlJsErNeSrhQGgLk9qqaBBfeumC10lNfIIriO1fvUzass7lvBe2KaaMlhwnNFvdkeA
CcziPn9847F+ONj3hXfi/EsEOTvZ+wTsTo5qLEemAQaGfV/xI4uSA9zv2Dy0qSdUVu7jEZFZMNJl
8RiQWtWW5zn+ck4x3LYOj5QsVxOehEN/l19+yOJa+w36r/lP0pnDW0HYHwEmPRhFYJYOz3tGXnct
e0dwH8F+rZGpjCEWr4bA/zaOmNtjHLclq3oY1GQSNw/lYOC5vzgUCnc3S7uCSGubuHOO0pxVipZV
b/ucBXA2SBRb47BUitOltCOnHS87Q4lKPTv5YIJ+BSgLr3qhjY05VB88BtVUCuCJhccS4QmKygvs
7Plar4EfQVYDNVto0E73ZjMput4bmwq2rYFDfuKEA4BJ864cXn3UgrYdSpTafgQzpaU8d0r5lS1e
CzgiZ6ikgMI/UYX91Y0BddE77MzRHsXkluJ0ud7A8mTNSbMbfdf/WEJ5W2kf8GcEeNB1Mp2JE2tg
WgD8n/1Xab4Umi0ughOpFeMTdD7SVTK/eWCHIQJ0yLStaYyxLGXFaBHTHolcV1e3PXgSNDxuTPYa
jJM6ZccjCFpVlqdMJslARC1wyiMJPAqD3agJPLKMFF1pf/AzNdIC0Oub2+3BvHwrcUOBxFhQqmjf
kGo5/Kh+56mE+XLA7BkwoNf4Hf+doFZb/UF9nufp5UtEzow5ukCpiW3h0AXmwqAJ8igDYevXLBML
zAzuw3jypWQTH7uLkSmqzwfX/XcsbPEfifbe5AMCqx5keL5h8QBG5vARVVWLYLpAbJI31xxl+YEr
rdK7k5T+CgXj79I5GqN65Fu+xZ3qRT09NOG1PXXqnGy3qejOuYbFDibPDWEN2b6mz8jop4H8fuvL
txkjeHHIKlu4amf0i9sxmruHdhgPlwdQJXkazhDMPJjNZGLnH4+CqSwOG1tCZTHHkTgcsa/8LDHX
7Y2lMycDjwar3Q/M91fegGwcbQ/buf5L/iqov0KLU9S15wd7Iik4yLgF8AYwhA5zzWOEfN5YeYlj
lleiPxJOZnlNj45NPOIcrGYDGGPpRjMOBWqa/MBvCxf88GfRKNSvGIw4X3FQmKjMblcKpaG+JBuJ
AQ2b2dLU0CDJQ8dz3KbfBByDIco+8CPZefflmX1+xmtTVD1nL78SUqPlbm+tmZyQgJJWlxCNnJ55
AiBumPA4vWYQ87tqTxjvjHsv1Ho8LogoncUw1bwy3FeckPhCL/xDm3LI6YWIBLwLCtLvap+f6i6B
+hAz7ZZo6WPsesVTBJrH1SOkqT8gBxHzRYDvNfHsSoIP9rYmlKp/boOLHSBsCB67xle+gDBh2UDQ
bvwYhUZDlXkwjKQN70zuMDusFSLGPfIqjErx5MhAUAtD7LDWE6RZU6KEZuI/M2icCtdlhFDBVwVg
izg+f2RXugSkvVVMyyYr1gb8tjlyZEhAlkbRQDtSukxgIi58fWE0NHIzbPX/52jUSaHRzfqtEAwQ
un/u6iRRh+o1qkouzlMLEDh+Ks3GWziLbsMn0zz8BLSA4FpHjSbKC+3f/6LSMTYtjtwXFZyzpMs6
P7TqcPDSIB2sawbGkwTGsOiI3kqJ8sszgwo9FedX/r531d5WPajVhpgDhMZbPjqm0sLfxKG6lsce
PyP9BXdF4gdwerAwNzsOfxM4vRF5W51aj4QWlZHPLfDC8DeN+S3xi0dm6fGN/ZF9lxFQiDXY0C8B
4s0HHtiShA+y6mqxaOfso0numym3dK6p/Ukkl9mHmlCoccajq/BBdAlJ8/0cEq8PStmqvIe1lh/c
adACgZZB2MzDXAzwGatOvLQmlAoLDjRQWXJPEggrlyhlOfYVoIyjfhFcodoNjvam6SmWZplSUskS
/ULqrEAMMb5jYc0FBUT6KPy1PEIf2ECMLIIiJ3Rcu1Z44zLAXEQFLnlRvGtHZI/4vvFeYnE8VQt4
F01K9Js/Iw6/Ll2vswnxOaA+RJaNcBnpwaC5pBOHrCdGoQirMGPFeQHB4QcXOUw5AAiXMXi0eWV9
um2G5T66/Qm1zKqsA1OhFUoCGw5/jt3E7hewtWzRSQva3/XgRfO/FMTalZI8yawsFQSy8FnFaOSm
qdviCtJCjog4aFe2kEpQ6lTBOovjXGYxVjKMilGUftsVafV1YEo20HqaZQInir6nlY6yKawPTiR5
Qje7dh5mHW26zKYzbj3asNAgX/SjZKkbf5TXRb8+v08KqNDwAn2pr17KePsYOAX288dXtQ7WfdQO
jlMdLXAHVLsZkcEsvHwjwi/KF3fGJ4ssaVfYVTya5KyMHV+K+2RBg5TNv3PjpShS4jymjqp/lQre
kuuuYaMFTKq22eYy2Nyx/Eb7ieYoytgEQvx140uAYbyC6BOByC16RNXlENasQ8FnIU/5wlWwym/1
JB0pig04xdcshg3j9bmkNcyy/hERqEmjlCUWw1q7Qw74CDIYO+WUVsdJSjuW30Zg8hNfxaQl1eR5
SuRCgxF3tQThgAHMnjS4pICewGuE6MuDcI+9edKv5p/vMWL4dxUZdBn4TiwhjVFtV0jUwQkYt+aw
bwvX6xAy3V1Ln4EhXfntmXjHmBSak6FRM6HsEL5SaY7lMAxbJSOqIB4EPufOZ01Ce9l4a40+rNbf
2xKOCbFnXc7kK0oKm1/4p4Cp9IK7BjB13WdF1/QtKqqP8sU6KaxImZJYg4ZDU4LF/yaom9oPDoXh
aTaZcDk0u/3ReQoJ+Uzww90Y32z60R4QdZr4W4QJZx2wLBoxQAhKKQh7hscYHr2SrKN3ymm8xGoZ
Vsg3JmpqRn7uBBBJws+uNTbiITTOq9+HOfT4fnqrMcw8DP4sw+nd2lTG32PZapBbpcVixDsbGXjG
lipEIFqpCkWvLACq6xq02PmnNGnfPP2WiLacTCNqwfeh6AOnE0MrfXARZpzOHV4qjNo76L0z7/Hh
BtbE1pvDXllWGv1Q8SQVVrGjoyvMNO35OXh97VJLQ0g8CDM8aRNOFWLaTAvxeEIFPzPEFaDoWNIf
Hx73LdUt7LarAI4Fn71uJxIdVbcwCQ+vSLPOVnoNHNqb18xskWvhtZid+V2MtqilI8ENGZ0474c0
MH+WObMz4qsaaN3isk3SQ64RUiqbby81Pc5w37UML+0MLfVZZLmOIU8zFe3ijW0RnZt5s2h2ZLAn
pUbprkJ269JKZLLzA+a1kDP10B85A/iaBuA3EybBGO0n2+k5pn0/8eLAHijrHtpswcM8ptMMLYuR
dHYOc71oE9KwFuhz1Z4TCUdsi/XQPiMs6/g1p00TI5CWO83o94+5GwXKPRFdly21FsgzAJEtcFsn
YrhTiv8W5RmqAAks1yZJAK+ZRMgTuQlLMgmYl5NJ3OS5sbOBCimzPL2aBC8HKUo1BD8wMvjlzw6b
FVKvzLbhNrTme6kY837kHNanS+Gw8EBTdorXYpum9BvnlRSedfX885JZotLs8CzResDxcQxtfUYv
PwESQwwDrtNPjJEYpBuDrBg6OXglZDcOybs50Xbe2VVNfsnwA1MLW+tOv21idnw268MFeujCEEVv
r7/yGk1lKTH+3KuocJE3JuwA3XR4uliAG0IhLx16/2JKq6esL+msQIOGrMvRj3bHB7KT3njNHUDc
M4YVCi6QTOBVoG9WrPOlKFys4IwUOnoa6uOOwEThUnu1jOnHFC2Xwqj8rQrQbtJ00Y/DvspaIH/l
xtb9NpBbzHRwPa9pGh4wFbVTHU1C/JaTQ9T6Q1Qq5e/7RwKgnTjwSRKHgKNpP+vSLjWdw3lXKmtg
khrsp/AnjM1gFsslkiTLCtWP1BAh+le+YsdRipDpzOVtvDYX/s8Z3kzAC9KL8fjD9hUl6U53CE0v
wO/cTcgHGjZOLFpEdS2VfnFJ1s6Eyddp3kryJbFZs8q/MSPHy4FVjLGdMB6ZuAg5f8SdXNon4PHw
qVNI0zxbwgcpasT11suOuwTqr3TJaYN+iUFMeelvz+aZBaq3+ITfDBusY3P3kUzf778soV1F1FQS
dPuTRe+0iT+qDoX5f6Xiljt1cEX+Z4GKBylXQ0/maImM+stw9Cr86+sOT5pAy2bQh82VHCsa8Azj
Y/oFfmuW65MLa0tnlXrSsrjXk62IREIl43lOobo4/5pGE/QWWxx1xBT9A0PHDFDh7N/oKk71jVWX
32kQmKwDHuszW0duw8ufVm/Pn8/VIcWMowGEjP5BxXw7fTwaa65TqEe9PDCf8roIoDPKCjIDPI3M
0rskY4Ghkpmb/F8Q3/4pk4pUer+Om+eIjpWxaNUY164HS1UnOPk5TTELJZ0Kwau3zumuQub1lWgJ
IkkrJPvH9adt1FhPPQKsNNtu6wremQPJBpov92NDWk5VOrBbGXL4aiXGJAR6I5Upbt6U3YXelckK
R+Cwyhi6OuTlT0U13IP66YWvKZAxeEbtums74JU7bmV00MUcmNeXBzUqVgY65H1EShR75NxOdYPn
GyrN5zwfV/k7ANTu1T7tgYIJ+W5GwHcIXtF8KWhGBNvlfTUN+zBGBoIFaLf/ITAU9uRr7GvDdt5P
KD3sPPCdWq0cH2Mo5z4wyq3VmsHQkrOf2x0IxW2S4UKbYaRDU4f0YRGvM5/zd0CuOlwcGm4VG80u
oF/DN8i2p0tAbmzbABJ4EonLweWKV0ocGb1CysDQ0wthZJ5Fhts9ub9E5y8NAdCf5ZEN3/8HLIgP
DsIY86lfs8UpR3DdEkJI+aJIJ1Rw2H1MHqfNV3zthmwz0b2LbqITPb0HHneanC5+4BIEx0fN60cf
fU+CZcQVZ123DL4kJXeLN1l6+NMeJgNvNMcngmLz3kL3hUA7vvF4g1L55CHrF3E+lAudrzQy/ESJ
//pl1ZOuMx8kgC2c7bcJhLg2VCFEdQqmSlBdxGb89VjIjgOQOA/ca/iEMFfla2ruHymQHNhk7xEx
li1SRexsAINFw60JOzVUQKbSjxQX1qR4DlYDdtEUWM/WOk2VVhBYIuqBwVUEe/H+5lKAxQR5B54n
Y2rwebB6EeNpoxF7BHw/k9Zkh7ZG3TOOmz7GRpF706K8zBuZCcWFlEMxYxrrHVAHieMBeCAQJCg9
iuJODuW2x6m+y14RhGBeiFgnndX1Kr6fkKxnLpX/A28PjZilbGbJNhFTwtsOdfbNFDhKwiXeWJ/f
Cb3fNgzZd24TuxaQdpbqZEgszmHQwgXc7LZG1D3/aTlprLCgxqI40hdCvEe6EaxPG9ruaa7qpK8H
2woIZlLAoekBpQdmBBeid647PfjPvjvQeP6zhc5ojqgxN4uHsP9GuKJ3bZ1kbMSE4AfAwSkCssqp
DyLx9qdbZNqVI19wNQzJ+CZQWZUf3fNza3jco+QCr8EG5RwMin54fxxrfpksZele0PBvQ84mxwbR
ua1Wd8u7+4TNlvAKq+q0zuz9v0Z6hwDB+YIgEEc/noK3fbvMQDd7DsOTtIWmHg3XNpTRtampciqi
VwZOEFBgjD1g7tpJMpv+gqSPCdiw7ye4L8zuw0CkvdaJd82rUbzNAIGhreKG0r7z+Dmruwp/EeGZ
5BMHY4vsPiP+vHrL8qjl3AT0C4+WbEuEWVU63O0rk6GVSEdep6LlMscTbpYuv4mnz7DEPZvOXaD6
ktmlPEYxz9qW8rsmcJtVbBXnN9y7nN1bLMSMKdk5k7DtH4Auir5dQ1QYLjsvfRGir5XLdr+8SanX
9z9bd/0ufsTpeoNvfuQG53zh9EvVGtQCLjBm2R560HF1knsBwywMZ/2S0tMvpGuYdg2Vt0/Ei8c+
CytDOObmU0uJdWLFcfPeYhk0+n/th/EgqxMRv6HUCLJ250nP8PVsRlWcESNRFOh87KWdpRH/j7qa
8ekOWBeaHiBvXBNNO2fs3p81SjJN8wYiFbHGlOyrkRVJVJsS4+vOGC3lpBnAqcs88rXNEbJwDiS4
e7A4n3yn3LNmp0ryxxaAVc+sgpcvkC7t4pD8M6zfB91QkGG1zhotQuKrCStqgGIhs9UvNDVCvmaM
DTPe3yr03U2QFn2ge/UzBTmFkw11teS4Osjpi4WdfcreCe8pvUfMZShkXplh0KVPZyjubrgWTN92
QgKY274CRwFt+tT4SRzGvt1DJVSl4J+3xTMhF5kKV89NwMmEQ7xvZHEaBi8mjE4Ya7zmMv/dWdT6
tFsQqKOaaFRX0rlY9YuV35iFtbaFKvmXLQ9qTvA48MBD2/36oVWRGGXIs4+SM5apzM0bm7g4ZMtA
JwMFnTpIrGq4P8pgQ/rmbVVHyqSCPrz/zra2Z5ROaJjWt7fIF9ZXob1kE7+taCDMwIzDRN7s9I0c
tzLJbpZTUbJ9oB5pDmgF0fN0Q36kBVnvCZY8oi5Ip6DEEj3Khsf4EjXn26cr9jjoLThQL5VwlNXf
WEgEMPjjZtLA45gN0gqdCv2jsW0ERtpgvdD59FCDFOYMXWY9a1GvPw/Qa2YCdeug4U0PDXWaP8fX
VrzNkMdu6ltU76RmS6FBf1haUlIOdkC9VszQjIu3eOndVrnJGJqxkedK4xSWSelIq5oiT+oemHK8
PO3KVQ5Yg5E5uSTVU6eZ3HIQL5i9ndqBIAr1bGvJoLSxvQhaedA1WbBaIygI7h8u+RkEl6c+CpST
NsHLl7S/B2g1BhPcsE1EToi4UsxroHkQ1Ui+EK3Dr6F5GajheXuJhSgtUojAZ6YWZMIRanKk2o8i
GwwWDrzhLbalfJydDY5h4yFTRwW5+YS+BqwFGV+pF/xZgy/YX631C4+kGqZsCEDJ0Hu3gOkpouwC
nf1AuG1QMDVspr+zyjZprTlGk+RhOTcIAtTj33AkiBdwDrdw7pN7p4sqNDGro1RMRy0wiXEjuShF
kZD5Mh694vNded9xcUBpQVTbNGSpv4bwzHczPENdGwRWEB/j9jX8OZ1Tb9dFHVELGAB5rummwFKD
RwIoXP/xUE1ff3vNzz4aYQxDh8mXKPxJadZdhGO8LzpmYDjiKAyOmgQH3/eYqW8AWr0PYo59JeAi
j6NQXZVIFcr52O49qCoW2mTTZHOyIYJBlBcQkb1qD5v1kqp3kE7fAqbEbiMqRzd9sl30Z5ZkMlvq
u6168iOcBidK+B9b8mlLe464e28wWDGwl/4V1m/dkebhijXheIX/oHimnHW37iVhN6cAtp0PSzrq
xXIzR5T4K6JykAo4YJkcyMLUHMcjYsc27rz2+ccKr8esB4Ey4B3esorFWuVvRvPrM5ApSbWzh8Qv
+CMe2nmi1Y7aE9+/hQUm50XEiAxgXvNbzpJahopaKDaDkxA/esuC7H4TOEPdjI0tNlO07WAuhqn9
nBAJSPhwzc6mAq8sDXjBSXtbQnafK5sD0a/SjSYKAGi+KUzMMvG/6W9Xwmt6SvmjimEpxMxhBLyg
VZNwr83tdkYxEGZAPGHAbn5P+mGBhTguE/vPpKyhfL2bdTlvbewYgjzvfjqC79ZoLh4p1NCoz4DR
SPjZ5bsgYCu3E3jPiH/BotQ/UNkPa2aGueHU7J8YD1GWtZBmLnKtxoPeR7xOwgHsu3ykJOJMByba
Ys4n9RSaKlVaeE1cVJFoOXFDGmpd60DlCEx1y8AMtixFuKBHpmtLKkjL0jHi6QN7j7rn4yGokIgo
AJwPALgVpBoINZzAU+MFm9oODb6zZnlMokC7ACDEtOm95SWJOoyaZuGAHh0V9BoO6BEEWCg7tXmt
ecDjjLbys3Yv7jvkFY/LJNi6h+L25ZvUv+uCaicVvTzU/q91lLYphh3RqXJ139SMYRUmS+c7+c7C
IziqNcUJhstslYMpvnIWnYv0fDalHLGjFKGAd74QBNK9QwIPI1G1G46ouGk1w6nPW0nL2ce2h94v
CqsWZRgFBVBTmY9mxBYMI7iboolcOZm469WQFfr6XJR0Fw4C2sdUrxeGJZVTjNRgJSaj3GDGmhGq
LhOPyAfNaIjMsIBx/g8OHpRWce600ed3bWZc33iXA12Tuk7ZACXMKK53hJ3S3wiGNohhp08Dqz5I
su97Ltj8DrD076VVPW+A8VKiTDNneJ1q1IuhtATg/CqMBSlnb1APtZsHROy1QuMSWm3ujJjEHUfD
uk0Ag2NTq7BnPOZIWAfaSthd8Lxpse5VHXv/8n2VG4wEdB93w2sSJ9cG9JWYKCD3GoOpn7PdXQ03
jY/86si2gv0q1JssIzJxPEklGXivVsHYEWgdVxYMH3vRnP6FcyOW2X4SYFQ1TS565+vMQG9hqD3M
/KUMgKD03x2nTlYF8oL4M8eFCDKWAr2uBd5T7VbTXuCHagmYVtAzLMlHDyD+EDbQszacBIPlx4jV
1Fp1Qm8mKfuhDBU/d/OlOCH2dG323RDK4SYsWSsx7d994JbF78Gj80qqZgdiFMmAaxyvHpcd9CyB
jcFuKC2qTvRGDI4plXKyVvrwilOV7TUTuE1BvBvZBanQM3BiLNykSiWOSRb+E0ZgPxjnkgY275Pg
0Twure/KgngYWGHk1H5SrbPblmwn85BvQzW4pIS683y4DVKH8zcif4sGFgBAIDvGA/Agft/hmRC/
fohcCIDAmMsdio9nHlysjzsDpgm8UzNrhsJoPtpmcitRaHLKMOUutniXptpBvztsaVEwLg5Zbzxx
qC/L+aw6oLfkoKZzx6m6nkvY8evOJYfUQHaLrJGOVqvbqyJiLAyyBqgZYcMPLhLwX0Ozy2on3WD4
DWQ54FY07isHvNMwyMYadVBgNaDHSCu0gWSWAPkc2C2FS2Jwhau0v3jhFgjKwwBIv7Wo7J/LefEW
yI7rPW/reYKVTaHtGYkX8RydEVYIgerj2YtVUl6LGxlcEQGxDzgWls6TSehGuVhUl85DJjUIkCen
Oq/o/DZGpe5OWPU+3WSq154a46ZdE1WioG7V1Otp9USD6zOCBPFqaAM8wVi3fkduJ7zV0NKLdfdG
+rL35ktnDv4HFQA8EkpCKot8f6Ly7SnB1sxqvgtFeRr3riHMm3Ueu0pVjh+6XsvOvHFgkng4OqI6
RNyeiSSl4f0i6TrQNHxYkv2xIe43Z6ZS/7j2cOAGMP0PatUxbr2lf1AOa7G53glnkPhdmnFpR7e8
X/nCybc6EE3fwU62fds0Qx7oJ2nlqkpl0+scLX88EXOC4RriNnZ+4xVWgccwvWrXlKPvZCZovbEd
2/oTeclPm3/rzUEe1OeM7YOl298Zmy842b6XerAgCNCkDkBTWYKdjgV7b64tRKwom55TZUqkA7i9
50QK3m7txdWRKSpHsqQM/Kz3QZRodc8qC99KT3rQmXtZCj73e+TWf3MBLbHs4L2NLCJx1dx1XhGC
a6TfK3xTi63xYOVfBNe9m4t4+LOZKVJy0ul2VHARs3xbq4eugGKgwcEgiwPg29NmNFpZMtVUbFeF
qcIQrBdLhVNBO1IimkXC08MIZEI/sZ824oqDW0MEwLSjETT2zlW3VMqnqBV9iYF6IKQt70eXs5Y0
Qe4hPkXrk3YhWcgXXOSF9TgMW7Nhu/xcc0ljke3xrDPjCKGP7z7ozWXL8pIzm8KNHz5tW9XXoeCZ
4QM8Sd6FY/YbUREnEPVm+QfRw1sLQqTfNDl+0OYKAVfzscf9K1D/cAg4qqr/olc8EwmxRi1GjnvC
9d0w5OEg6oM5ATmh0SWZsq0e5MelLX4SlBJ2hCyDleoZW1ExHfBu3O9wZFW06Dt/z2pwWgyw7ZIh
v9XhBeVk4RG9TVKfeux1n91F1kIoszMiPPF6rSFSVyPa7UDbeOgLcUkVX69BAcDVjl+AwPtwBLNy
iHrAfK6zxYX5Jf6elPoSnnOOWGLXhNC8//38/o+3osuzMwDhNgEiU74f5VnEpiXiclEE1KFNTm3w
LOvbJcskrCgtUfTrSEVac0l26wDqY/K+Lz0elfvjzuOvYLnrQg62pSbmNeSYWczZ1bxxlgXHMWnZ
zCCR0Uzg9vEBIC31r+S03sE6LqF0QWn1QB6NH6btp5XkQ4WWe2ElF1kYHISD6fW38D+GwTWPWC50
0/weOvV0qoB0441NQwcCeeBTrKZGFc8IySgwxoGzttPq02/SNQQwz1zk39yHG4+ILJWqIGIssKnV
Yt1MEaEs3qY2aO4lF5Nb3F0xaQnO5556HJEipX8roCoGnq2n6KV/W7sSzI2UOTr9fRfCYVcpkjs8
e95ts516DPX+1ZAN5SqO8/u5IIHMI+HYe9f5WnVL8eKbJFMdIC5fPiPk4IjczVkJ2nlPcaLvpryS
d/6WqNT0CkNJii7O3A8LZUN80tOSRiwbiI4VXkYDVnRBFB5ytPV6g6jPH8nHLMXOGQfjEUhoDc3x
87r/cnElHzL1DVQqT0L18s66YlhlorMKY8tpL+ezKvRTLmpQpXpcHR9rq22oeb5mFALG7dYPtfVU
CmSrNnd2T8bvTvFIWApt338zuzXHcUdOXBAtsMzZbh32b7FCNI0vkW1WCkzpKRsKFCDONiT6q3Ik
IoSHph8FjIioyJOb/fuUaLJ+ZUtGhfaI4PKti0hT6+jfiiQyZS2xanCUAiSOcHQvV5ZmX9Zp/RHa
WuLzt4LV5uHgggBImhnmQZaSAUxgibu9TFcbxCmVzvcH57898EK10t6+JjEpRN5O3LRNRWjlC8Ip
+x7E+Hr5K5buqmH+YWkzu83NW2zQ8lOBVyeL2TD0VMah24+oSUfR6P3HHZ2vjppfVnhjhS+fJMAJ
yQgFeOn/y0ksl+hBiNSd1HZIEWiN8sXMfZPBZipIQ4jYfgNQPaRFzz4iI01QUcUDTy+eR6xMKH3Q
cz+mJe/1FE0W9u4DwuXHeXLeNxZmXoIoErOAX6ci62N1xB8vnOezbJ31wosbRfKHBx9DzlVAFTKq
hj9+8tt4Wx8D9c5d4P1uYQq32aqXbzE3riI+KJZIZExdHLhaDAT8nkRSSSlOCPk67rRvd2GGl1X5
7EgcVYrRdwhNjlxFFc6esyRvkPTCX0PcBHvSwzjr6TZRJhcw41wzpxLdGaxeQdc6dgYok/1XUDkT
L5Uz1P9+g7noBTbCKU1HlwI6b22+vC4txKNYOqclMhsAjjpC0o71uls5jrX0KAJotq2FhsrF6fTJ
dhdWh2/qbwKVn17emlWqZM8c7A95Tn04eC45jXj/KpRIG5GRuPryNF63IFCIPKVMXAzc4vo99rHc
n06NvGWumIlYMRlqsadpzqHNCbbm+ZIQPI7atZQVjq9zxSQOUOugStPmgfOlbHXsWK8J8/5HJQ7Y
NXQQnAqRuuP1eMWd9ZdpeWlemByy+YNre61UXUPQOuWhRsVBut8rmEFow28xtxxV/mH74gJYqMEr
+k88eTCDNMxBnPo3Gd9AAs9fV3bT4NMuuYAO9h4JQTTFWBm7hjenhUwFljfL3GR/JvN53k7a2pww
8EeUM/6e/vcrE75AVJzSkHSXyFOf0187V/saF0Z37rDGZCFUqqWF1vKIC53z3VzjjDNZsZebvAUv
hr01X9HKXmOh1eidQ1gvYW/g+EbSpXa16WmBD8hQGbd7CGLfJkNU9eV9jHsJUJ0HZiu0aJGCxvmH
Pcmp57Q6aojUbtgdv41x3COq/MpZ/7BIed5qtGSsrwO554hrOgrzRXqgADUPJMZS0O4DTjwBTUx6
DqBt8oXgVsAVmdA63JK3BfkbdokEui10CmgSxfvMqjnVc5F2I9F8q84xGhjtFW8sYgWv4tTr7blH
b8TWaHtOplvaApCeTpUPPHzlObrb57+Zmefpd7Z+vEuLsSyQaYD46ZbDu1SrZYH6SZqMOLmO/O+T
kROIcUvSPkWGA1ihy3E5cx+h8FhcKdW4qCzsJGF15yEbRgdFjcSHAPQg9JqWp2mtoSfs43i+CAQJ
KI0QcERP8mmkkBS+ZhKbvlHjQxi/c5OmHNji5n3z8+QaF/UGaVvW4jF0zGoV6viu7ZYUtqX/cWdw
eNC9Xr7C2A+vQGvPZb1KwYe/XozsKrjFkr2HoqXzqM74wIt0gwN1T5A6MWZK2ug8LDS4b6U3BgUz
y+4YQRvjWz0yBH06w9CtWk8OAlWn8Q0vF3Egg6vmCL7c8Wvx/I+c+js8cPUjBmRa28dbJ/aQkH9Q
sWmnfBvW5FompJxOpmWuB84I3QnnEoe8MgJ3tiCaxacDXxu2xe66Bxx74OitmiWhlIxod2QZJeJI
UEPedi7vEM53KEzi3767OrECVF0HRWsnNi6sEMwwef/+6K0MdLdpfxHX0bwfk7m1trfQrlGr9hi4
vr2YlGWTVNjcxRqj/y17eSmC82lq0ce7vjWPcG/vV3OYAFMP+yfR55I/KrcQCJixe0FkfdYSjNTz
I1ZwAvLt1gAhAAOQHoWnd+Kj7hKKL1ceT63BiTO73RlP85/CZh2rfZ9t65U5xPwlFyCzJ9kCnCG8
dj38BGLcyKDOfNnTLehy+QF5fwl/eL8DJfjJNEeqoucCS6a+cAJZblT9vQ0UBtYRQC1aGUcknYNw
YLpCzI5be/uCr0L8v9E1cDvOfxRaUz8fkIcFwHqQPU02RrglbVW82bprBivNQReSOcr2DM7FI3hq
kqK1Pc+4uYkMx5KInf0Y0VcseE7btH+7G32ZdThr2OE9TlsL0PbOug6M1N84ovYsfHMPLrKZNvo/
jpbGFBOWd2qXc6UObh8Oe5doK/xUuAbZvKlw2v09Zn+bVO7O85uqb4v7GJ+d5W8ErE9FJF3ivkbJ
tXf3yTvngB7QkOH1ZzNR0JOw21VfIKTDNttC7FwnN34gWE+SwYrI6R7hKm4+P1WzVEjUEs5EVhw6
WAXCrULa8tsTlCKt0iwJZy5hc0iIlCDnbo2/AQMZCsNy5sauqQiiSIpilnDWwXjAnYXHWY0luWu4
1znGxW19gPijszwQLy3Kbjp8NtebCqbRXvzXP2ltA7EftWzAzXFlrasFAAJf1natK1OOZ7lrf7ar
a0kE86jJwIINraMGeZWayI2530ASwUlMy3Hrn8eRW2cq3ph0YnVwyHbjznPz1H7tpR3BCNfV3Ha4
ZZ4CV7IyyPHr8pNMGTuH7ma7HSSir3fBCSjxeJxHh1/rxiSiYmxt+v0qEBWzgKk55hKLaO15g9ge
W/6Ht2kNu5Px33UrBRX6o/g+aPqanoK1EQ1D+cEYQoV1tH2b2HGzipS7KfVz36BLanZG/Gb7LRaC
RVm7czGsiIcdMVczs5YviTGovnxB1LThNbzmGm12GXf9bOHZ5HAJx0Ki6JRs85Hbj8JLOY9tesKH
M9Bk5yySjlHGEnZmn0tEteN4YWPB9frANp5z2fneDnWgB7Ai/tuUNHPgjlnp7nPwrvZK+J3Nu3XA
rfsmzPPhojYTTE5HjjHdtqc2gjjdccY5oReMda+V/uBQYVJAxrzE+aTJimK0G/6SWssCokSvxh63
CG14y1iXscyyfce6zvnXA9tS6ag29WsrzGpEtuyVrQhUGizra/NWBryD8ky4X6A6PAGaUlQv6OWm
U3KPqwlIkPd7sfAUBx8Q19xHH4HD/R8SUajHBurh7OI1TGwzPUbU6MOt17YZS1xerIgxTZDsk93f
sKPzE/8xTN1Z0YtRiLpLPD+JlBzMehU298e3FKPD/RDcSyjr78+HcxuCb4/eBU9X7qWo2PvNiLBK
dVhMNkzSqskrtQ9D1MLjv1y2eSwxk5wNVSoGVLB0mdWv2XkJXRaNJlhkoOTfC6KGcYoHRCcLeZc0
65/BqtORyVo9g7my1AXMalJhsSzV5V5oMYf0TSeWXqwrpXpPYHaOKQGyg2fGC+SxECrCTdhYlk2/
wHmaagNjRcEds9l9hr8QrXxDgLEgY1EI6uEaEeBNIubXNFMlEN8baCC6P4x3YbCuVLnkUGgWOclX
rOGDiFjb4HwPQY7UqNvT5k92O0Z1z7kBzHO1r3fblK+MEz6Kuf0/5R0JEQn4Neoq1u2f6SpBHHF9
2kv02e3paZQfqO/pzourzB0RF6wBodHhwL6MgtnmRrmPuBKnySK1h4tFbOD7TTRfTEcgBXbhgGNi
ak1bnfmV29hltOsXC673ixfPaLSvYfcupZqYgm2fLFp5Esvot1+gb0MxLzX+gzw7/dyG/fp4Tm8r
D1+E55Son7D9MR48F6W7d5EtA7stfg12cvxqVZwCTP6P2TalsguQx/RI8/VuOqEYU4DoTWKNgP1u
A4MMK7QVJ4n6vFUC6sHQDw5mSs5dOdXaRYd2Bdb3PV/OdLdKCUdJZzF1yHUz9U1Yw6ktrqKdW5q1
JmI7BwElvDKhMZa/wEz7ubGHyJmNyQ3smSCsLJ7UWAdJsfM/rFgltuwk6hONZsON9lcyN80ddC2z
xIlK0jSGIV14cYnBUh+GqtrLy7EUZZZdRAZqr9/0xQOsc9eHSxSz4LFbhzqnsvr/RELHvg5flpub
YAD+6NRSxdVIbTp5YMKMCbEV44+lAP6Gz4uQZF/YWWvxtprsgpVJUHbLpJelLlMaNFO+MYd+AA9s
prSltoxZHLwQGCU6ASwOkVLv+gO3uIuYalU1lkySFL7KFNVfVedKVYHOqQD1hhaFVWdovbSpVmzJ
efytz4G3fJ0UqwqWJK8w1Khkqoh0OhFIb7VOCTxHRXs10f8UO+efqAKw2//LF7qw5rftPLxj1pZU
caFxcH7DiPr7SRpwDyK2KI5zb9vj9mCFtSyhFsALGVxUY5FTWnBE2lfeBbSiRF6tC4yJfsuUVruI
c3quJDjxQqbmRWJyOoh/scR5JLIhh4sC6UaphsYjaB7h9C2r8/MIJ0AaWSZvhOQdBtNB2gt/Rf0G
44SxBpWePd0OLW80S6Een1Shuxl45F7ZJxidgyk+xZ95DJuumzlmPhHF23FY1yfQCuHxnNt1tTLY
atZLaA9k6uhfR+6uD1Qo4Icch7znN0n7MofewJ1i5TJMdB3kt5Xd3J3WRxXAyduVyF5Yz9DWAuff
Qel75Dv431HNhS9d9+D5bKCyuyOzIfc46pEvElqiHzgAzb6vm1ENWXLV0WUZYun98SjZQAztiRH0
3x3+hTmz+MPfd+caGfsW0fNx+KH47Qj9J/Li/+gaYYuIPiyJ1rXohOEx1h2dTkPCm6wvLO83e5TS
OdRP9kUGL1jf3DryObYapBnfwn4AB1ZIyGDeBOlO8va8ckS2rTB/s9FzwYwU9scru4N6keDEn1Om
Wkpto3ztdOd55b9UX+DUfXv5xslcv+4sk9SJ0xI5B23itA0b3ueER4B33R8RO+h1FuztzI0T1WM2
UhMqknr8G/a1AMqbtB/kdthExm5B6d0vIZ0hWeojd5T1ElJof+8xkg2KhfGKROexaH+U8n8HKiBG
UKOzXr4Zoe++27YVZHab3Id4t60nz/uOYDNINkViiLDTkzXwMGtnu+zmemgq4Y0LdRR0AW0nXDwE
j5KfHzo3bd9IWFDo/QAvjR0mPj7xPaIbv2txxXdXjP1Df5ecvgBv5dpvQtPbMNUzVyWTpweYTcWb
jsNQvtP2a677b2QxFky3ZTfpaK0TBOXur1bw5uTloPzJmqvlSUaIVk9u+Csh4THOWEdoh6nkOBIB
k2nkoYNaoVw60/BWuWE/NZmmfNWAUaTfS3UbMO9Mlf+CdlfqKBJJjW0TNfM3+k+gvbpIz4fzo5E6
wcSvkjvlNJF1zgFccww9JdrfqITq80wSkBpkXI94EDYuSPvOUqT72uLmI7ItqEdWEWQnU5KW8eSH
zyJf/6PCV13Bg+y1mybYzHA2kz0wUSQUagBccWHXNp7qRFpHO2KP5VYZ6QxclpwYBlIc7gGZwmWo
7VCtMwxd4pFboPpT9TF5mCFKOfuS1hsg3FP3iW9+m4kkAwDWei4FQx3ninR1pqDiU+LQ3j6v3IBj
IEyRndizYchLgORz8Q+vDzh8fBhuV68QF9ieJLzABWABlbqN83ay/jK33kl1x4z7wpWIplVXFYLn
z+3d0pQCDRAH5SxtB8kdRk5xjofH3louJh1tSxRhT6oapOv16Y32UMUUpSBMZWoLxiDByHTfB1eU
e8VTb2ucXLqtqhJHJ2f8vG+OCnYg5yusw3ge1zJRT4RKLTQ2THypOD05+pDq6eDrYrEuHE/6dA94
GGtX9aRZ4rK5OEHPNEPV+6Da2gUDtQchExMmR+qog7lvmCVF+UjYB3qekoTPNy6g/cErhdgiq/+e
e+67TtEaTN+0v6C7KhrzQ4pnUkXQgI1qD4j/d3PKH8DR82e4pjSsvcMFc/seNZ9EOeon+nChFI/l
GiJ8nw55kKN3EHB/AS4icqdShOW1js+XgRI5x9yQzSQoC7/WLQuaXdaIiZl8kaH9fb75KVluAcaD
uv0Kmhc6fagyBpxRNfkgDIJL6EhvKwNgoTPqIS0TiMgpCEQmCdF9A47wXCrz/8FAJpvIgK45yin9
/70+clYCiKhLVto+doo76NpeEgP1HPkdXCP+p/ujYugloT94H+fOUbIRKhFNoybhLIS57bOov2Cz
Fu/pRrj7Jjo2SexbtdOb34HqTZJm5d2qT61gJP31yALI9fF3UGOkoeHU9LvWaoi+twkiA4KO/3mw
vZbUBaFwow6TA0add0AVrCTcU6CV7Xfvitjzo7fn8D8RzzrNL/A5FK5Kl2y/Zjikv5Ofb83RFfCH
EV22XSruF64CGXFCdOYDNe9EyFq53Br8E2I+TKyWSCMiqzmfIViRSEzH3wHJMhyStlvC3YgwnIJp
UFs8wR5CgaKwjQl3WyrKv4xDJFZPH4lI1gprC2ZMDAs3eD2lueBglPNoznL6CbQyN94iNdqMMWWr
jAB4K6f6GRf/T8wnLxm/ZrlCism/ccEIOD3p/ZPbV5K9hDTy7gf8l+ZFhGA2BL2ERSYApN1jle40
EZ5IP3UepDbiJgbEvdmyt6ybepdyWCp+OLUwWCBE3ZlhNE0V2AtkLqKG3s2pchx2wG0IZYIXZPuS
eoKy6Ncqm9Lc30Rwr7owDgi9LsoC/UdzOgGN4ufKq9htpTLu/nyw7ujZkBI1kc11j0l6hfuvq4DO
ecggjF1UtbQiTDX2egdjKs6MqttozoG4t/vq2+fq+1+hWLqg4otNQCzLjHUKcJ5o2BaAmyqH0q61
H+18KqAcXeu3m/cjnjwWjkF5BMudI5vM/MhlHKtjQ+UrVINZu2k7B53NCUSaPBeco1WMALU3jntd
1hhtYnpPWXYVmY2tIn4ah9VAMP88mYbkiRCNA4D/poDAI0sCaXXBb7BJslKRER4dh1C4tRT1EAxd
gdVbV90Gzsu7LfloLjUYizJdnmrJ0ddSi/RXPA/7aMwc8gwFv5Px0/mVAF3OKjJgqSaTAuvFLEGo
+L0BuyqHQ3zIvOe/ekqJ9pZdKlrKx1+LRn11YoJVJlbJ87AR50bo6MEHgB5SC1R7oO55kyTpYPs1
BPVlADefv1O05g0XZBLeyuFiSQwIUAY3dKTADFHB14V8IS7zu/kMoMnLKbMhAhU/FitVWaAlIN5p
s3/UylscfMjbROy5MBKJlZSBkJZpFr/RLXSUn6CCqZlMg9nd1gI9+SDj2GPXeB6b1YlP+reLjO/O
HpdwyxHdtgoIAhCrgSXvKBzkObUvaL0NeI2lVBLcucG34Rd85SWSaKjvX8t/k66zbgpilNCOLfqs
sUIUTZqHuojnKSOSYDBNdq7HidpM6gLqRtGm2r9jWIU6xNVlJFj+3qxJhDxC7e5DefYgF/gDts/g
HM6PAwGLQ31LlRFZ8pVOidJ+qFCnDAyRSlwaTb1xgjp27DSQUM28qeWzTV4wVkV5rzexWF0oYQcD
3FpxECIWCAB5kBxAv+e8L7apJFpp0wDvNhGVPwSLscpHLCBoBjp/Xl5tKXnLyc7XxwBLRtt1b3xM
4VsIWjMRpl324qDijQMtHIunO3HCKxqGiCX6bf4GPmvqwJ6ABQd6SlOxTqYkzWZowoJ4s7fQmf3M
yul2tcmcJAiLm3/r0olyy03GTN/bMb5s7D67NYRfiwWmuv/Qvv3g9dw88TJMnFlT3GJY2zinlUaw
EDO8bkgVQQP0tvJAihSgmiNvDxbmvzmnfA4AhntWkrcxbQR+uM7vhoW/c0h1TPx9pJMFmovZ2TcS
tQAOUU7Lfc9GPfyJDMHMCSgF380PSYAFodCu/kAeI76/NGfOX9GAGdOM5lX/HHjfqbYGFbjUYO5z
xueHJ3CAnPI0/d1xvYRgdbHAVNrk2w/fu/x3gQ92UmvTz5Cd+kXnIjOkqU4aw+i72+xfFkq4iYbg
TLhLYPAzySenFRZw5Hjx9lgt1wvEOkPp2+OdHV+jIsgQ9GR5hPqKnHupYzCsLA44RLuDxyqIrMpb
xLOMyzVl1Xn7Pfdvkq95CUUuKsYnmOxcuy/2aUAgkTXJUjWmB0BUhD13ncdOaDZHaMuYShuwjNsW
D+ea4GBn9R2dpQu8m6UqTpoEnz0n6wsuw/uZ+Crg0nSpbUmuyHSDuPtZYKhULf3MesF80WMODOhB
84pjumTVZgWO9MwZME+3ilFJL/gjZpl8zOKC9UrenAkxbxA0fud38oZA1rAvqOvlldTe2c3GgI2J
EZgia+WcOwcA2R8ZH+HLEkQ9KmIgYS8LP15pTc7rS3VU04cF4Bam/Yx4vfjRu7qKwRz0Q7rw+qjI
MygED2z3TpFuFkS0mh7e+e2OLYBVvnHW/u1wjUJ9j+0Dax2nz2p87R2CvDZjgFMpSf/9ZINSQW4S
HYaj5mgwEca89wHlY8fe3oBkQqEdBqciq9t1Tkmr5ZrOiwFfAXLT9TY2vWfacENBqYTVORxuYeJ5
S97zBBqisaC87Y8nhCAKSp+FlJj/ZDwjSvytD0QBEzBaCoDNcmQVvopPMc+mR1spYLZCSJy8P/Nv
zAqFc2jZXFZD3c+km/BbcW6IM5c0G8OxTfAAsYbEwbLB99w2s7CYPVec52FDlAVijE6FnP0tRwGe
OFAs5BAlrHpBOEPN9u6n+eR1WUW4/DD+XyN1N8U6Zl+KgOgL9aD6jLhvLJxGDXoNn3OadkYnlDVb
ATOVMV7xKskaSW+aq435KEMt3Bhm+snFY3xUnM9H0VCtTjt/xtZoicE2FMAPETOHIsVfIoJDBcL5
leN0bPlr9pUA6P31SnGmJpmBUgbEPuYbviam1qZ8u1YeRnchIFirNfiV8abcdKdAnAA21CHiQ4pT
Xk4hAFIzYrcA5zZEBPOGDvdFwroWXjRFx4uuQEkHZYb1DaN6BBmybfCZ7JdUc97NwXDURGX0RMbE
yNJc5ut/DfiKvaslAUsUa+FX/QKpxKIX3YHO1xFrM2WKqPCRA9fnt1GuG9GbOYvkqtPfESNlP7Oo
T2tKrpH52gQE6n+nlEPe13PQBlXW7ZlUW9iq4JX81FG4ukc1RqeoWNkPz+uDluFoY47evun3tuHQ
xUPDXmXm34PDYHPZ3OJzB2t/kFFzZ/SgVPlKbJaJQuv2pyIcBWpG1xy3Y8sIjymNr4qQGeT9OUk4
LHAsLUZhYyud8uJ0CyFu1k3799FU3YkuLhinKxF+4LXC9ZiwG2vmpw6PmfxvZSHal6Fma+pUOUzH
xuEeKtsVJi8e3NfIJefM2aneIk/24vyxUceJIeigE5Hnb6OUK2S6mBSCk/r2wCOuIrnKuEWIJA4i
bY2S2a0cD3ZzESpXe/Hy2SFxJkBq5HjKH9y7oyS22hyzXY2jxup9hYC/Q1ZthCq0xQW16tSpKOYP
HGxPyfTqLvmbU8aBKSoB10WP1DjByslYi3mtzh4me1pQ/hm2S+PWmQvGp+m/5SNpQKBTG0nmREVg
6dxlmfTCqjRIGOmqUPEQjvipRmf+XA3ueqzRUlfdjAiSKvU2ok8BY71CzJyJFfd3tn5vNFk8fEbX
IDbnXCeisZk758JBrHM+y0ex3L3nlSXmlImTu8tfYYFXYdDcX4NsueX3V6f3vVS4FkFESzQk5Ggk
kF9GcxQxltGbENYkvxDCMHxE42v3gzc1c2VmiGE3Zm1qESEYTIK7EZJTtMIv5Yr3Gy0xsn8yAUdA
E+3ljdVrGRO/yK4dbnc9n8D9slMD4ju+nbpdWcZhyYmmCZOMKeF5b+ZDsZu1n8hofZZepHerE6Dm
O0ufFMxU3I5qjhfmAaKBLqTkBDYiYrGWrziXt5+TolXhgv7d/CldMMgRrQKJYoVU9kVTWu34sSJc
6a9yGMOHEiO9XSQx79kdH5N/5UIlxIM9pbtialbI+c3l4UbbKu1k8F45PDFUoLXMezx3GjZTxi5Q
pKdEYzKJTqs+cYhHztgWPq6VIsMBPX6PQf4N/hhhWxyYcUE9K9wAYU0KwpvbsiEw6jSdCnXr01wi
+WWMwuVfXSJK/4FtxmQthZf3v/tU85JWiotwjxF3XGesxS9abu8bD8XS8plKEifLcJug0xvDzuPu
GOqB/J0zVCYR1x+Ge/UNuLb7r1UkGAL60hMenX9Xt7tAUIOGdKmepy1n6za8rILKeySUfo68mYTD
nIq7UlqXGD3UaPmFCxWUBspvZGWgeiNLbznk6+no+bT/+DDbQ0u00nOG+F3GTfyViwVitwZmHoZ4
Y7b2v2s0ZznjUC7KJc4How8XdaVchUO+DZlPeU8eePe6UTyEoZ/lNkl8npgl2JBhtslbHdm+8jMw
ADmFTTDHRjKq/HYUMAe7XvjkveVlJs6HZZ3x4d/UX3nyxgHCuW9GZNng4c0k75DZJXItJcenxUT2
c4oqdspmkyaRHQmAcHy051uqq0bywgGVv2Zn24B/GudGLlFB5gpFGWfTzZMn0xDsNY88stPUSxXd
Eoj87L6TlPVtljUf3DbPEWUodpbz+qIakMNp0RmdFIPdeWk+5gyxQa5bBDxat/qpF0UmdVcRLNXv
mxyS9IIx1cKRxdGcymAEuCn3W2XiiHfeYNWPVBI9CHcKprUtkv08nb51DYbggUIOVeUftX4YeUOV
nrN/zmns5vbG+wSixWx0LwdxF9kwRJuOrz+EatFY1gqLcnteDdTx5z40SJx5hv9wMvVKdsxQU3R6
TjTCNQ35lOnaXZesjsyiB+v1UVZ1sHNMXB1DFZQsAJv2r/qf97wDgSgKpY0qYTgtfFLC1mujYnGh
F9ejXfexVBvZnnRJi3hCj1VghX+nrlYK/ZDHYBQvvPynOHD9CeN0GUmO1vPw8A7FAALKTgMLdEZM
EjzWIX8S310+I6TvSoa7rCJ1FE4kmatUMa4iJGjDAI4bE/EfWaYuYciMLjppB6cb6HuIq2bccT3C
TglMW3lfLWEwCkLfmxjAtfMh9v8dfJXsGp9rQagTnsmlwLzQrSTzdNhA6VIIVwTXwcqqF1j5poaO
NLExGm2Lrhb5EuCzE8sAtgI/lVOeu9gR2XFArwvngylR21NlUcjNx2Uk3p9g3N9HMbVZ+YoGdA/5
2GedE7bfm9Rw76PDawWcOkg/PvM51O6fPE5q8gphS4pZowLWO0YABXqtcYO8n4x+Tgm4i36Vpr6w
OXKRbW0jcUhSYwXtJy1UDSYQBuOJV/9C8RN76/oECW/MWObnh2ZYrQ6g3Ykm9P6wzxKdpSjaYKLX
k3DwIGe2JuDvy0xrGc31gZlHHuvZbNaigPSL/22VVbL1Nc8GWp86n9mGJ7rQjHr1OuV3F+voZuHN
db5vtn5aOlDrsxq7m45m9uttvUZSE356n2Kp+GRUPgg3DAhlTEB1OIu6Y1lekss8el0vLCLlZwfw
4wluo2mVPsDHauLmFC0p5X3MYcudGyUqquyga+a7QXYCL7W9pm2Pjpu/RtdMEIF5DHfZrQGy8Yak
rpq4SSP+ONWvOZKEYX3y39T6teHG0hhjlrdy1Z5yok/osnVM1Sq1EGXTlGN08ljWL214xnBJGd7x
SnR3kCZyfg129N29ywRlJ3MlDiAoZLqj3z7GqfFoQFUGGVZqNgCNF327O3JTLGUdoqAowXaaJlI/
Jn+etLybB15iCmftlaP/IN4rNvG/O+z6f2iFGe6sLuPqXR6cdeCZfNeAU6TDyFJ2ppnWCggsoefN
abl7K/0Mp2ozNAm4xIxPopXg/SXZ6oJw7ZzAQFhU2Xs2U857PnHJtHj3fnn3PvyFyeiVcvJDF3ov
obvsJSKMk/APwf9u6YO+ECz1OjL9mZMnbDNiCK8lkz3lLYxaBokODkiVT8o8ui+IsZv+2vC2Hirj
HvpaW74n2ChFwieG9Ge9AuQojA9l7gW73UwxTTwE1UBTZ6otutyIg7sWdZBXe8A9S5shbhQ3hf8c
ka0wrDVtFk57S6t/NO8ABwhhXmSX29Ry1rB0JMU46HOvC2HYLYGaTdKFUZLmMmUzNXN2+ZvTcgHf
R2Cc9i7V59oGIjg/ifvttGtoz8fX/bKgVp8OKF3YY0TbpkSl0sIxrW/5xrlFQk3C5XhyBSwxm7GC
kp7XXwmiH3RGTUmMGKDMrL2gI824RYk+/VAmDVnmjPQrhg22zxd066hXQgrCS0b24HQ9LDJFBbwf
Jyd0u4dGmiAaN0nngE2RzZ7VgK10GdVKwajViK/Ecgeow5De0XL/O5xCqAlGjhcUzJ0iCnTb+k8T
jX1o3Dx+736CJOXqDzGlB3Z6F652vGkCUy4ba/e8CgkA0tUWctJUZaLnEXjPeWZuTAJPsOu8JnFH
PEb3dn6xytfMGRqGSvNhDT81dqePOgqikhuNEcWgzX5WfCebCxHnJoFFH2MVcO4QY/unlZJADJnu
799CdtPMdk+CRZvZcCHRccRBerK4i4i3QGtLm4tzoMU/LYE3eanNpQy7oANM60jykkWmLvH8D4lq
7HQ9O0YtnYaUY4Xbw7qFofsisvZtleZOCp127hFbY1SvYYneD6G/Jfhz5Fy/9FsJM4WJovKuPdo2
X7SMaERFf4U5Cuy2iSl7o4kbEfxtp/OwlwQlDGkfT5Qz4N+996ETNGd1r1UvcyFrbr9B4erndcfW
U7WQF0eebHs8XaFqg1Q+7XnyRzHQ2winFMrAlRhubF7U+652CfLZylWfxK73GVSYjuPqs6WDthfX
ghG4NShrigjI4OMF5CLIABDbAC/OSqkTQ970LESZ6d5T5vOZeWffR2wzDDkDt6rgBGegBN4pw9AG
i1B7CiGL5LSuJBbnTQjdGwQ9uVEnEfqQ7/5AXiscwyt5zUel9KAj/X1aKMNq/G1HvoN4oZ0h0Ti8
Y09ZWvSq7XCDAK75GoqTii9y4WYFKeMNZ9UNlECqw8Aff2j3noe5bs4oo7c5AcFUnfVJAIpaoE4e
gLXKsdmU9hmPedvLOecD1r5ZT3dpn2aObp7uuQqaz07hTwqedJ2Ld/dSwzdmKSTnNbZjU9IHifyN
U+bBJ8uJ4XkRaWeeaZ6T/ZDxNN6GbMpXJZnZDR0iPbDp1YjVktAwug/GnwTVCnyMPVmmoY9evl7C
tpvCT0YKT4jBKgNYJ/RP/Wdv7o+Daxv7DYSXtynwEoXuRwPniMMtPQeTzMd4eLNocGvaN+JjKBU0
DkoANTgCv8Z0UxdLJ05h0BSTenZw9XKKjMeep+BZo/i2qzFU/xqIleaY4EGNMvsqRBMd+vhWL8mZ
KvM+Jly2YqlZAKkBxFNUD5fiHPu2nIz5KmPD6oA3Zy70uquPrsLqJjgGju2uRJ47/85HNea9vWkL
h+3TFLXiRBcBB1pLoyBbvGeb2CM8Apc24dBN6RxDZQuLwLpiFff+XpD8VvNtZ1qCtPJV3W8U9rP4
NSYELs6hKN8VwN/lBZkVek0Jz+8TaxZnESUe8rvJNIoVWL+W7Np/KDxEg35HthwsDRterxXcOrB/
+ga8v2yE0BJF0rdIzNBU6rc07wQqzy+PpN0l2IjN0zZDQGrUDRUgsTa1F2o0Bvb/8+q52RRmRytu
A0H6f1WvhiSFDbxRZKcLFHZ5x3qL4oHGuvt/VZmHnUBmM2J/dmC6ScRp9G/5wE1LE/73Pa3iirZ0
P3Jbcfn3lK+PzRKgmyda6pfDvM4hZQ6/DFUM0kNs09lRXTEOLxXzSkURmmsNOj4NdbzG9qlHv7Hd
Uqm4J3GOLjvwLmJxB75kYMNxP7E6ET1YuB3RH/T7Giw7hv35BLOmRaghYQxCNhvLhxuQ7Htn/KuT
dagcviwk1yt+dfFii2pTG5dMHezBB0QAdwWyVjL+1WFSp8gDKfhuVTEp9rrn9OY8rJiIcWBmhjn/
QNujpcVlmtuqoR0dObzc9+KuE7wfucqUHKZvaAr6vc+ZvipwCOtSrG/2sHsuQ/bLdmNKcjShypkT
3mU6r6dfNdx4+IvPvrchWx1XTDfFEy2nKIon40e8oAbsrnsy+tMY0432Ow7OzAXdp6zt8yoKb107
BpJKC117fpN1ahkZDmhNSwdIouWX4qbdfB3xdaBCIh7SgXQP+77SAO/OHdygZjir3so13XrlegE6
WLyCxreI4BOyLucR8u5Bb4T5qWX6Mn2dkKynm9I8taqeXsYSICD4wnIyglSr7CLxEfz4G8pSQYTk
XZ4ZFmWrKPaHfgR/VzEt+99DK7LgpPxtouwZk0/4R/PJantQNoiXi1r7pyQYa4eEbZR4wEDkV1eQ
TJmwPJJC8DukhkDHgOw1l/CQ68dwc9fRox5Lasym7Ksj4n1ZiExeIhAp5HtItbYVVGfE4QG94jAy
wZ1CLSWFaUFiM/Ew7tCvQ9EGoXsrJgoan3U8Km/K3EdvgCUob7QUNbGngiIPN0gDRjOaPRBI8r6V
8I9etpF43XhLm0fk3F4rVJBBxeZ7AAXMrTerau2+E/Iiah6a7MHxNGsMbTof3lAayzNOmrHNk5cB
+JNujYiI+cVjEWlNuOKtbJcqFhr55qeZ/SdLIx3E8Es2y+8eQUhw2H7rz2Q4khDFFBAcppFzTF1M
f8J6MbO2SM8bHv5Sn+dsDI0f888nm9gb0KVgMV33y2jzbu/LZsr/FqfKX2p0z/bIwhqVeMDNQFzm
GOw00+be1ObB/Nw0mO6HRXNmKlvg9QnU9s1BxVcdVf22hVd/dH4jU6sKEsooQEYPR+656/x6ZmY2
grKtrgrQFsf2vjY56mbBQwi2gsCLSG5i3kCbSBcoluwG54sDFhySxRUCJ5ZTM4Di3n2HD0tjIdqg
17CPHlrYy4WMx99+OnMskiwd1/pGcDKMsl+X6g85VX08eRS+Lx5DinnmJwocLdNCqiCFUHLa0sXJ
jvltAK6bUd2m9MiGg7D1m4io84kVYjlBzbDKZcmWHqNEUrOmSNCFksDEUuZXvJRV/TmjwhCx1EGY
JEgLFndlOuE/LeCbadDDwgIqWkcCI9LMPUQocvrZh5bVO1IB5bIaTUY6Ul4jqg9PI5/9jGLgCtZM
Lh8oRx7Gjc/gnYRsikiEQVFEndWlwxN5tGver5Tv4I77BpNuRsfSZvb/9egLG+OlefvqtOh+PiKs
bnvalA8JAAE7dUE6aBdSGxDZ685fVbBA042Q4Y3h0SKbONyuyqImZ69h4jIzph8kz4HCke2nclU4
zrig8l/gJci9yTxp39ZjKb4GK+xL7cpNOPDja0gqFHC87udiBMBaiqr5giTPfAe15sK3p2vKawmH
rtSgP7ijNG/CjngJG5fU5P5t6DdBCh+mNZU3HsdRZ4iaRdUJo9fL6SptcQSzzI1DbgvqzqR9EYWS
IihEsnTh1basDnqQMoqyJcgWK9wvJFHE2fnWtjoB6p0DX/nPmdxqM9p9BYsXyJNUr3Zez42V09cp
X6TqW1n04j8YXNjHxvsIx2oIClasHguo0OkhWZcPG2S1On3fE/UebtjRF+4/JciKTgrZm0h3yesw
80NGxS5mghm25PmjCy2GXYm1xveMNqGR74wY8dCU29uhtPWbw9fBgsQiFoadaB4703wzs5FwCW09
S3ZhIfYob52/u15/vorz+WHsAk8pjnQ5M48HZ9tB75dUc8GKq48nrMdjJvL6NXDWTqrILzBMtIBa
CZEyIAlEvnE7G7I7yuJibKsi8nV/0zT22cmugtYnYZdlGDlhZRFGRpOiEfZ5hDzIPlD02VeP5AId
0bX1Pos8N4Gm16QTdYvThZsSRnc7RHBlBRVwgSFEG9h1339Od8LN6Lgd6Q12/LvAL4bk2FTkjjZn
71aqn4xSFpsEpZj4JC0xnLbV4noBpjprCHGtHNnadMpi2KaaRlOE3SAdhPm7FynPE4m4SQDrM01X
0ehplEdBnlHNKJagbf4xf/hb6pcKQDn2lU98gtRs8n9IF/tUm1F+TIvwtxae205dufCDFykNzwRv
2v9Oz3qUAp+lH2VSS3+cDg1JBRCWNu1w/TvWfY5abZ+qxrB8kK1QraWqrl0OfKgn3bbVpZx9PvdO
zquWuAMdX0JLh32XfbR9gIYn+Ec7rxhkWXu5BcsJoeZSMID4h84PI+bHEgHnwljOjdOrgdxQTawe
JSSR4UdpgejIwfKSajUEwA+PtYRC1LNHA1CnmKx2OHWzhJQtyXC6CtWJXV7L6I+DoRbpOYuNhkjR
fg79sbaBoYJCpCkurDDwUiaa2Ey0IXnMhPbx7ddeT0gmjALscuKnUBx5mW6fWIHgHwFMxjIdnz3l
Ot3jAWD6baYTxIppedW3QSGXSq3CPCK2yjudTqH25lQM8nQi7wfgSNMMVCvBGcquW0vtA0Dlhck9
m9p2lJ0z25qGitbSxuPgTjDyneiOn9UbZhygoPxdQoo2P630uKSIN3394+2zhFlKvBiy5VT2XYl5
TULksbXy4X/ZpZ76vNeuzseM+ZrvEJRwLrxQgSkC2B/WRDLyAlI9Pz5pmfvOuZWcWbm9aPvEww1k
JcT0oc9P685o0QLxoQBColtygT90Ze0NL9OMi4HTETkSXcLPwa0Ox/VfhmPc7dKawUzgWdbGAQAB
PP1Vsf2i+mQUKVmGB9c+7WevUcT88f9e2z7s3d4CiU4lpPLuYOUSR5e3WpR5m8NOwB+eYJsG53e9
y4CfUkunVKf0mbUf6Mjkj0foGg6TORrD7fvvjfhO38I6LBBXgziCpghpxaecXKDDfGA8anMYrSKj
uB4y7RVKpfWNs/x3wFLSCligmeyrjC3OORd7+XWEq2GFA/xGDh4oaguUpFUi9yLsUBXJaCVE0ku+
cCQ7kXkla/ruRdAnNO53gHP0L+eJBjzzhi4l2u+qaqo5Y+JvWHkk4xc8fRxoWbqHOtt6HbHdkAq5
a750mQmsr5vk9ePD3MgwULuDfNQa6paeJJvb0wvmrWoyu2bMCLHbms2T7ie8vHcJQcjN/FdcsZgp
q3o5sbhFlUMUkcp5yqsxN2NdJ/U3RS7EdIxSSn0+3pIvzVy3IHJrrjZvRuR23Ag83kBi6F+RmlKk
pkC5XY7FAZ6+aOOVPfMn335Eyt0zvQ3HomGFVErqNkXgAIIzwucOJ4Zi5olyHGK6bUlyierU1boK
nfGSjNxpKjsPH9pHJHnYY105i23pRHDKT8Asvx8UElSolGNyvkWYbvskaHXMZiwVT+paPOq2Mgdg
ZV4kj3shx1IRNPqfT/Z4FdIo5rMZ137YyzS97rEl5dl3fyoFuS4WEEjZg1g5wvkFuvL765XFgSJD
lagQbS4D3yegoCwKFQmVBPYftYjEAHJhqfZUFZRxhNv1Jj4PWVXdSKAXUkvpSv4ozXw+3vzZ7jKR
wz07yLZFU+qcqIZgYvs8OxfVUrefzpdTw8oJQZoN6jPlu1Yw1paNx0B3+9pAbDtr+7JtDKna5haY
UBwSgRlqPY1t7TSDqIZPz3/s+MgGchKue7knHOB5NZWY8wQS7pJPPsbiCAACWBbomZ2t1/x5aqn4
kR4YwX1y0ZyqofgceoiRgF96u/AexyTh4zqYXxqhuNB62KnIzYloY8CJnkPCjT1Wff1R31wCPa38
cgoZoBy1YJC69TzA/wuwVAX44Zub0s12B3Swiy+dl2N/ft1wp2/nF5cCS+UIzYldv/cC0v6jQ8dh
JtpNa1i9YRTkjEVdP2hwONOh2Zefm4/W3o8KE/tobeS0CTr3lo2itqsLEm8v4z0Ab60ZdxfXVnKG
mi7lAp8v6enQKpnA6JuW9Rnw2ZZv3FgCbg7LujVIrWSvSjQYxCG3/MBC0xN+sjP0BUzxGwItYyMe
hdgF2KQXHLsXlUmsZGL1XK/PTX+bfTkGfutMkNjWXYciRXt3ayWta4/nImOk4BWxJu1xmHyn0Zlq
8PEwzNwyPVMNlMNMmEwMiIXysfV22MMiZ5oZkaFV9bqVtmpOzwoTyuBfutA2vMcZdhc13KINACoh
lD2I7apgvt+g1SoTic9ItUyovShF9d2C7eqavuigoTlTdL/0xX0Zt1ppp39X75s9gqEeAJSGUoJk
awr1PnE9sDbDO1JI36lYc7VjJmQhLTsgJ2Cj/ihjE61ZE2jt/wZxWDo7HMyi4KiEC9NprjpTxrsd
3Ub0MjnoFLZuzTqOJFL4QYR1gqZRw/g9s8PkiBK1jQeVMt0IQ2hpGZo+17KyrAvGQfrV0K5ArbLD
KXYG2WPVoCJ18XwQa6G+AO8F80VOYMUtsxB2R0qSLGl/jRB0l1hiUheskNDJGlZS2LoA87sEhl1y
q1fF9Beo8fkRj5ICtBQZMHMsAG/VN6U254ALF/8nGmzbE+V5OFJFr2fyDbHa1gOgqHBQCFY1MF7y
bgtQDanhrJkSc33VkqUCvfBNT5It3TpywVB+CvaF8UUUNU1KFZPuHppgpXqruvj6UGV0H8THtPzt
69A8Y4GAXs17EqpDp6Wi731Rpn92e6mmDHlfkXcngQfMKshgczaL2WKgEUr+a/AzVcmkNZ6ZTUmD
/1q767TTtb5b5ionJAGnSltj1GS3FZqRMyDhgx2sZMLwEi8KiUZVTuYvCsNlF8BQ1UTbappms7YK
fucLMIeYrsuJiozbu+OkWrpukrnj/vgZaGuC1Sd1FL8ZsRZGgAyptIh/LOTVGlC8i190tv4zhbAe
+6y+NCzish7pv8s5wH1fDShkYRDAsDIiIlt4RkekFL0K9Ye+GSGauvJkZksTvRVrVw4W8kVh+vxE
Ov7cXB9KAYoI/y2fbj0OoZrmtHQWNDk+WtNDra1WYxa5KqMKDh6kmKkaTqxuY1KAk3ZvihFguJMt
k9CaNwK1EQl+VVlYRuqKcdjrffMlwoKGUuDPWDRJgcBnRajATOkPOwo7jFyYCeCCchIXtOW+df3m
SWAwtQezeTTpq2vwVkmKVXVHdOWPS7xB1lhlCb3x+O/k6vB2R/2uW8Xs4VGaWmua/+P9/wdHBhT2
DoAudT7uaKelKbRnu8XxexH5sFA094wL13FuecnC3dPnAQGJwDwxXtHkBWz2WwooR5UMmWqBu/8K
2xHO9kFFqYXdjHNL6PkGjfuIi3obBzNBByERvLFdhoq7xe/dr/g957T6ur0npfTbLZA/PqjZ1hr3
4B6wnAlXJVCcoAq/B0xMz7bu9JFJtSqR5IIwi0g6d9f+Y1/LkH0Ccmz0vE/UVS9C4S5Migyf82S9
birkJklS0KK3vAbahiRsxzqmyUzPsh/PNvQ32I+iwrja3yPmt1Oqcd0xgYW6AQlIUGrSpjHoQUC0
TmiFh6C/dhODwRGXHSUbx8fZ+AbOFbj/RGVEokN5sN3+OtU2hTGuRQX1tAu1GrLdVGepND8iZo+h
i9GVeSiS4zw9Y9OZRbZWkglmzCXW+3k9HSyHaxMyBy2MJhxuKRbAL7EuBYYMfWzJnH5N4OiZ3G1c
kbYlkCqI9+VioLLcjwiVQNP2SmhJYI/b1NmttZ0XdpeU9+y4U7/pS1YE77UVfljElTgy7KAQL/vz
pn31nq+Q87cSk0Urq4jjyujNpgKglJiByTfEqYVmyEA8jblK9B/RV60VL1OxGvfwqEcuY5cI6xyt
uJjIYB+8qTrhGyKjaVmeB3JyocOxeAHfz+1aN+hUZYagWf3cV3otl0f+M+VP7PESqcWwnTd47aWc
N+KcN4uPL3Y5pLeNU0XpbbpFKX0JpAmeDH9423FhtGoDKb5ULVFJl2XxhS3Lg4pniRshMVJj9H0i
ap6XdATuodyptL0OF0bbOgGdUPoyKgtAxRwVU7Z0K41T6jL1AyRS6DRsZ+Z/yyJ9jR+w2C/e2JOd
zUsSaAQfR2L8q1kwnC2CUUWu7R9rA5SBIpKfEb+z2K9zSFZkjeu6GfVhhhTcKvCgRF+0x5LrA6KB
oDxEZi7fPa1dwL5Ivt1DTBlmbtaQ9lqifBOJuEkswUw9xFOVbid9Lfz4R1sN/lOCpEg8ox6HivYJ
zSt8oCAUs1Qb00rIoMRFh9gJzyFkDmIJZxROkWSYLqRHfA8VDlS5ltNq4+E185onfN3gyAvvuvuZ
RZiNC9iV0lfCVY7uABDNeX4ytjrKV6f8FPo1KkvPYDQuQ6VCoHs4XxnbZQ8aObDndC4edoQDg/2n
hHs+wCf3WJRbHeMLjnP2g4O5b2hrW2k7qGERDEbaTAuOVJgPPEF1Yyd1itY0g2nFFTI0aSqgUUQw
PzvFPnyMicdLM3kjmIzj6KoyP4ZAuSjSOTZgSPEZsl4m5fm4Okk6967goollex4+cWvMftBmQ8Z1
1+hPJHi0qgrHoT5G1yMROGbFQloGx9m4ABhSc0LvO8mVaSphLeNSxlFHdarblESef5QBixAGTNH9
VV+9ze10pb74ncEAyHcnImnrpV+uXaKiOT11GUKMnedFnAZOmRHNuljV/HKb4LfTT3A5/EJ5TLKa
I3KYJmYrxx+oXqjBJkVqaRKUsXXsyGWaBZuNkVQnMXHTA87TFntJBPUYGQAh6VQmYaPgN/RQfCfh
BhwI/M4rca+LOVR9QG4vh6ddLNpVwx4BqpO3xRgre9r/rWOIIq4KhTj9HRXTDlHZqw9UK4bOi+bK
b4V0jwZE1+q5apu5ZEjBTBZcVgG/l8V93vmeZak64Blo1sibbiJVe3mLzzcj9GDT8hLoEOqGwNXa
Zy8EQDOQQqpuJVElFJ7N5MlWvE3ybezIPjVLIMB2cKX+pume4DX60LL5YCGr7Y1yKCruFPpYur/S
MtNjPMKUA15xCJuwFkpgbEuwK7DQm8jfXMTFE83GQT7CcGCXU4vPzsq1XJpz8x6F9GMk6xkzUJEJ
VBXOCZSBwVJRO+6uupQBJwPYOUcZ8ZkC4OODND7tHZUOkuIA2IXVh9m9+9Gqr7qwN27m/qcNEM+T
/vUUeYvDtW3CCt4COjpKpCAkO6dGTwk7uyzJU/LJYBIe4JBae4FzGzwUR7UoW5mM2BN8kQzAgcD7
MXXz8oGMTopIJDbyNpPHLutzFuLMr99r2N0xJIcdMDlos7pRtbCumJKaSWmYzwlK0HCyASQfyb8A
dEJFJFU4dwrzIaiHYzTFcv31ucTM83vByT+YrGgprBOrAW3R9li2vevxGoDaEJprz4j60Z5zzUq+
QoubBuI08zBxzTSha7eoYdIBj+rHXTekEqS55uhxkFNDL9ByxNkk5cpxL3u0MCP5CmQ5HwvUbba9
Vcrj6QK/nuRJvI+tmo+bzTs39rDJOuELQxZPCPbG53mHpZ6tsdyS48Wni0GZkccUCqHu6ivFH2UF
GqWfHH8wuYw4GjUqW/dhLzllv+wbThWv195/ddoHWJUrQ7IegQMVuX7GVDIwcdOwOX04m+zkRxMN
HjH7SQg5rGS22mMjisYfVP1SJpvGbPeEZpjbukGMk805LHSJje42DUUjSBYL0P1upzCPpY6t3URH
eShPMmgfgqN2SQp4AbsYp0hF+1Orb90ID1lVMkwIEHpyia5o1Z3YCvo14YyzXEu8QAXQcBys1s/A
ghVCrW0D1qKKH0GY1VA1LuzlAqWSVV/+1FTlE3dggp9NkzYs/k1xSQTTgWtxl1d8VRXpVdlLYqwz
KcFkQJowZZ9bAArCCWRtZJ5UlmeqzRTIexKg3ueXd0i+lvE91u8LcmtTzdi7zuLvkS+10/pJYlXC
SJqibrqK/ttELTgQd2lnPND3uGRCTFp7E3Uwmnpc7MTS3HG/hGfAL6dsD0tTcaZKaCpzr9laBuQj
pyQKvmH3y7iz686ByuYdVLYOSk2FsSGGrHWp7PSE2dIZLccjnCRTknfikkCLKlKF0IoD+oJiFyFX
wuR1DbHm12AtXB6VTNzKgcP7asR0FIrF8EGw8QVdCPyjle36y/wjwhOhbvNpAm562T3EtH3BfdLc
m+1KiEGy/R362kVqhP6mJwmAb9hMmJX+76EOsatosUEHHR7c/06M5TSCSUQGPjVOsbXdsoDJqBj7
EW20pWTG50qVt+9iimshKrNr6bfEsjqrvcl4emv7v0IrJGox3zyuho8k/HE8zYakBJ9t0ndHIk6W
pcNf5lOnqVTljw59OvFe8i8D1P4hVXbfYnVnJQXSdkg9lv/PXoyqUIzYXHOXeLzHX1sMxfMAJUaE
Zb6pxYZEZnZPSHPPJewmV+7c1D5YAT+sAd/dcJmR2bpiPQ/641qoUVYzFoCEUruQRUwFjWzba8xb
2phgIvujBjdNZ6dzs3Bq7NXVP3dcvzo01dhM8Chb2jBulgu1X2dWpqZFgguwqAJ94dGQPfd1Mez1
jjCuH+qgqr5g1Jf3AJU0UbxhXmOx2lXSeiyppQllhsnhj2f/Khx/ZS87DS5efeFTUYWcbHCRLDrd
UdFQiO7EC9mDes3mjA3Ko9oMc8XlASbaLhElJGRROm/6DZ1i/DHp5hlgMvM3YV7G/kJ+x7MS1ps3
qPnKBDa/YyI8Osd/g6sD3YvhO0sSL6nXJAa9SHbKCwxT+vnuLJmoAINJotbtZ2eK2jNYSzES/J9B
iROJ4HocLe3fD34ubSJBO52nOAZBPhy6g2FZ9oeThnL21SP041a0PA8LubizHx+rk69V/LsEb+dr
jvc/0j2eJQ+yq6W0GpmEHqy+CxpDvUx4t1jnVnpbgr+D8gJDs1pea39FilRFg3jMolFToH80q93t
qip28UF4IvuaMfDJJ0rOIIVVUb4nT4CNl2FVtJr5QtuXgNMQj+KsyetbRvCp9dudaN2oR8rYbMXd
c1Vtb6ra/qymRpWejgiy61scwgCqDX9e/dZUhb+KSrkmwRB46+SPEzEFBDZBI2BJfk22JpPs9qJi
xeL4SN36Cr4UuT/BzLcTSsVcR/l/Qb326rsvO5M0fa6cMy8mlgui6LxLEK6mcz1ZAd74F8VvpsEg
/kHpTffftkSukCQOkc/wxRKwsKE54FUPrRQ0PTdJUWcQMdcVuoxXC8EWFWj6HByhwv7YulpIRzcR
FfT/iD08MWN9lxAhziqYJAwwquFRN2FhTrz4Sglnv4oBL6UmMKwO46gHeoeLVA/G25d3tqup1naK
2YMAau3LBoyPQvtwm//QXzdyRHUX7QWP6CR2zUNS5EDzXwugaC7mG+K77I4NqzrfibeY7hmZcRV+
5JmVnyuepOr0auIU4oajMMj8OIR6kJYbnrHZ3aG0zTqANQ3+Z8z6bmNKy7nuESIJRKRoZQDhqTVI
peeh3zEilKEEAks71TOcrz1vEdiqdq98ox8ebCNLPTcYKCGY1AgzdiAOusvKiW42qzszbbLpACPn
qRuMWREtMYkvQAg+LQiXaAWUDdugggGEScC5d1J+FvSSTCr//Vu8HTLUFKEIvvt6GnNUZp9COthx
/NoUSyObryQKMQ3d6UIm3tnJ/fIitMqy74K3KaAm/yiGaIdgAKh+HxfcLXkmzAlnw4dszaLL0NTE
bpwug6ixRH9DWLPvHFV9ufm6htowUt6maHNiuS7ADY7AE9zREjxPITTUjc9GmhTHckm2NVQHfkKu
T48GitKlSTiUaRpcjuFEkOf3+K4PXDBY5Wtgvsc6CWzOrsbPMWcL7vMXO3ESWJ+e/nXfV9lZeujR
dwyrTOHkY31uUTs+0s4WNfIokVhrartLCU3saJaXWf2YLhFDo7/O+2EgnHQPRGzRn6ur4mVuwWd0
oH+Sw9QWYnn2ljQDSJ8bIeetRKfbLpfYGtoSaVsnhjshJTQ6rszLhlUD1HiQlAone+xcseLZWRls
WuPEUqp9p6pTYYdkubZubord9I9NDbN0FnYf9g9DAeRKdUREAzLOQ17JmtyYqtxjexMRL2r5ATk8
y7ewAx7R80wi572Xmv+2NPhLxps0Iyy/CJgZZY/BhD/GSArwrXEdNvRtP8P3057SUsk4g7aewvdL
q3P7tVCIgMRiNS52woal+mTtKr1QX0rc+ArGR214EORUwtxGV2Jk499wLeoyHOGB+PhUShAOPQT7
0Q/zTWWnWCkHH3nDxEfPHip/3Jt12Ga10LnFdFVDFNRQ1fllT4I6iQZ2AsXScpmmrPeAcS5TDawl
1bCEriHMQ36F/EVfcFNogLzGlk0orKckrT4IThaxdSzqxOauKzCjx5wYu//UUfrcy6vz8nzRhv7c
LvMx6E3K+ND7PVkDUqAGS88zqcG6pdvGi7Ci/u/5BllPJ/S1XqlC+0D1UsDZ76XrXmh4nxtKkiag
Jb+w8MSdoxkwm/YlkaB0E5jHse6bhvMn17tLva1tIjm9QuH06yHQZftPy9R5ApC0dhGFcqKD54xI
DhEdujNsY5300D4A2pYQ3zu0h07bSr3BbfZrTheiuBnynXlStgn7JYBZYkdQcG2fRdGA28ZMHY9z
2xCTwWUOS1C+hoePyXXDtd++jFPGKMTVqY8jsK3gMBTSo25ZBoQCnYGUIkpePE5cWeHDUQl6koYS
t9M24nY0rS5QLeOOJALjdmme1kh2G2VtVSLysbrLnUDqvPfaETGd7r4lbn+ZqCmqUQON6tAnd1k9
qxJM1kyuH95KQnweembP935w7XSFFuSpDlOPQjdi0al+RcfMvCITacTipIDi7MyfvwazmJaehuoa
L8OAtS9eXhlZpMF1tu+NcLoWbAlOP55bwQwJPQZ05y3rzmI4UMpSvleMcNOKG2Pf9Ruxwq+wVa9F
iA/8ybjP1yDX0fUjxpcgLMxL5rOVs7I7e6MJ+2k8dKHZDgtLDYQ+MNE9CEIgnKlDE9pQ/GaLr3EM
3jC5BERFOb40U0XT5l2JyByB1vLqGFuYGaIfR5+kn3rNZo8NZIMLOaSa1HTHerJGdzaGtxdnexbQ
bBXwxw/NuaRXIhPi5gBOC7w8KZ1UvwQOxa9i1eVUBKIthoRWjiU4RlRDV4xEM9tyh2CfroHKftip
23Bd6bfJ7FR0EYCYVbM83QiqcdbgVMwbNEV6qJPkCYLCF4T2Qm/dV5q1uzwSqBHqTpjtiOa/+O+I
FRCWUC1m0ska+OEy0gtgurkdZsaqux4hUdTFVMNzS6s9uaiEDBjcp4phaMwli61ty7eyJQOmL4Sc
NEx9GKkm1TnMuxcMJTD2oMeYoEirKqljvs4RMQdzQTglbGDIUzhuqLG+GyS8AfvS0ie42Al2PTfM
r3ww0KlZahPosb8/rEr8r9ZncXBipQ0mRnPtBjV41kH2tifHG3FH5GFWuBNYvA5XWH20N3QcoNp5
60k4n1qTBHpjJkXMFgyfYGzlVyisv5o8UvRyxJft9QaNSr9VK3biDjdvO32qI5QE5wzZM6N9x/Cp
r80LagMEK7ZhvThVgapQ+QJ9zFL7CLvvAYzgkAMjS5lI5IG/JOZJ1Pij4Voi9tthNrz+1LyIJLFP
/zswyHuv0k3VodW7gZ1C2c6OXPNdzuBgm/p/4lcwf+poSqpSt5HEk3C7AXF0+zoPhtXRp9V6CBVd
jS/iO2kBcutv8MxIL+I9+R5M2LEm6NVDMz1bPwrGKEjC0t11PJfGp7Nc4EP00wBPxZT1dsNQWiaa
1WVCYgFZhBkE0trEQTwJgue0hrHEcSEx4pgEdUqPIaw6wvJakMJM9CG9OkxZBhQX2nkdR81F+kA5
Ra9BvbTDrrMdv9lVh4vUIrLLWRBa5TqXtGuBKQ+kGPhlDcezowi2eNKuQRA4BoOnP5qrNK+3EPmd
FXSldDfYapMEMzA5ocXr3V0sH8j/FOo5/27svdlA4xcoQZAIpACkuK6SXdIjPcVUTTVYz4ibHpP/
b+ecGDUx/GTcdo/tJC3iohuFZpeW5BuD50mMp/LTA3TpTfdwyS2cnMJSIGfgu1WAY40d6C62FaLu
5WmsWUgpEf377sW9MvAzZo3RC6TvsHPSexyxHnn+unMpSebMlWgW+xymZPsN8gUVjB1V7My6+7MJ
K4C3HJahnM9U6tZpFwZ/G1RSHXDkqEJfhYFAiMm20n9FxjgOP7Cw0xiOvPuyn4ukXTtKMAZOUXDI
x2OqtUSE0Y0Nab6L4bEKiLxc5uzF7GCIUwkvHoKWZrScfKzF99zsIva/t8SPnMwqYT/s3INGK/+z
WfpyzanPS19+LxkUe7wtZ44HngzvrDY7um7z2Gmn9e6Y7eEPlswhdtuLH5Jby/jUk/XqGhwbMlkI
SjTJX5PYwpeNmGCypO48AfCdwHGXazhGMg3M+ywgX1SU7Y51slhfqigh+rfzQ79Tx+66bYE99oTZ
EHeNuFFp/FnVKhdPE01ypOUU1xY0SAdO2A44xs9H5lNwt2iumhgekHGWm5UT7V/lYIN037+MtnAT
rmxC7suWluU4spSIyYsBLZWOZgnXvfZa3opNVt6dy8K3e8A5mg5IYWFsteMfIh6SJ+/FdF3jvorA
dbFKjBUciZ2mCOQwugDbhRRZJsEKZ4s916u67lU01R4N88Y6GnIT8nZDjQy4hsCKS/NiA/BjChnG
9GQbT9f/FCnc3f9j3f49ifO/Z0ShOBxqpxCeKv1CVK6rQCZ5wlvzr2j795Fdhe6TL8Uy06b6o+/v
gz/5I/jxZM13MOMB6mz3oBWlC5l9GX4Hd02SZPgOWGaRKYCake9mI+E0g8ec8CfmsMqex4xjkSHb
Potbk9orx9/CpGe73fkuPmeMITi1KT9bQrYznvhe/AOIyIl3UDR7ViKL8WWsHB7Nxu48DCzk6t2a
IiZfWolnFOwcq5Dvahx3WWPaCNjUQ8z/A+f1WU50FmJnTFJueIrmnM50DcMLWMA39rY4cmFEhvuk
zjm5mP8DSbaf8hiBRf09GcUkUEPAtfkjgN1zcv83tcSFwmPkp4B4XCG1XqXeHvYnj/W84Tuh6hyL
zR+nzcIbKx8ivhyY3bXHVI6G87vd4pmJmDnPHkt9YfaPDKBQISJYtPzDQPygdgJh9im/DKliu+UL
JC670YesmPPpdBAcDSmHwdg8CFNrv8OCrmSuxVnknNfs4ETk38hmKZPY06poVqw7MWbXq8fN7Osl
+ljijpe8ENCIxq4nMvloMIigFe5/6MXn6Qbts1bcJiPtdpV92JRpIjjwPeYqWvxGboAt6LNdB1ZQ
4Z90InIBhFQgKr26RpYUxZ1UXlUftQrVHoWVYQKM0yFq/O29G5PbWO5QlV1fDFH1G5etIGZBRb+/
GfX9X9CGxuZIPb89vIEnGv16BUVRgR2iO9pQNeRSZAXCWyGeH+YJ7QDDPTJlyJrXshhdeNQgS34W
Bn2FYRPBYHdWIUk9VjVdTODih6xU9P7/6ZVC5C0dQvAlSSQtym6emEqceuC1roUvaoLs0JPIIUIO
c+6dbrI9UYyxlbdFNjUh9lAp2qnQOSmBdqGE7HuMVvsl7hnIXbhn9YVDPfDXjjI5PSe3g1h1QNi6
ylwH1lklH+Oks7G71HT+pvX3fzTVmwD5pp/KMnLAXjnkGuOypwXUwZG8VLmyvjuIsPUAsgypsroz
XmwVEgrNN9r/ZlDmvEuxQgdWv8IZyhtympc9xEpTFy8Rki9XPb5JHIA+rz2NXZvMQfHMAdZvZnPc
1kvFf79z0/Tcedoa5JXI4qLkhtgkgcqExtr1DhyRjOu8l6mGq/AyNXbXh5MMYOeWO/ONYQpRXwz/
UttJ98tw6Q+wHuXA+ZV8nGBKKM2nNU4QROuu/HwGOytNoetLJakTFUa97AuJZc4iJ0LEqs0TG5Go
Cf6hJL/9c86lPXKDGkpKVJo1NAmaBIlmpbHpaUPlU/5FTJi67Mayv7aovKs1wolq7oUaTm0zx6lp
MONJ2nwoqsP8FnwG6E2OhzCRQ9M491+cNFJIwqaPX+eKPrev/hlIxbnxsI/d2Nat2RihaEDgp01l
k1y+o8QZPItbndrhOIt4ebyukyhP3gb4auDOwyrMvu8tMQTg5NlYHrVVRtl33eLMg1ccnjQGBI1X
NSmycEOwAk7MZ5XLR9BxL6n0qdhTN5DdumIeK/lwEjCmw9sLAyUjiksNjwDkee33A95Q4tmy3uP+
I0Qj3RCPxwakeByZYG055fBNO5aKk3Hdc4QLpLF8NSV/vx76t1jkKsHMY976UDWoNwDRYVwOxkY8
0hlROc+0opNZDWf4ukFybqS2a0hFfSpmAqKDricx1umy/HS7hhKsYSCtLxsvkqeYcPbaJJZ5bLW6
VzXTtop23fZZDuA8Wkwt+V3c9Zqa7AjV3LLY1gnTT5hkarGM9wkU9QUU88XxdloCw2a5CnJaxYDu
bkfxbBoJVCWLv+0bdmjnYzNRayMZ7MFbHoJ42XfN9iEJ+b7W8JNpcytVUoPHi8UrnHK0PKRfR3ly
IFzlkztn/66d1qHsh9WZNWaIxdoDbjm9RZQ/NJCXcSce7xImmP3XpPmHesLIUcVNYM4jc+fwis2K
gzjdShJR8Im/qlnpPtv3dbB82Kr54IrteFUvU/5OIMknOEHwddREFbMa+ra1q9e191ZtyGb7pOhH
1cVX/UnhUWIO/R6AC+sEnpAbr/o8vAySHMl5MG/L5cOlO1VQvLEYD2MRgea5mXn3MOk22LlSVNm0
7vg88Iw3Nmsn1gXzA8jvE40i1u3bNKeBkJbCKGglkj1T7fdsd90GK65AsD6gEf0aAnkZZwIAC3t9
eDTLQdDV62/aKaQziDJmHYsfrsxdoWW2qhz4qKT1CgxdrKtuDBic587LIbcUGFnGD62K/56Yg/HM
07NW6Geb4pDgzQEx4Egl4ScpVLYF9N1mJiNdLo0PGayNqlKnnnpv1COS90k/I3igmaYW13BaBmaE
KbW8GP3noBe8PSse2k4MI36amig+HH7G5syJ4qPytSIgXRc/U1SX7b70DtXd+fwnnnnuFyuAgv7M
yxyxcHO/8hzzZ788amBFNNsaC2zg5/GUIfx45DIwb311feuNjxt+iJ6MeuxCmHJP2RsOnPe26oJ9
42NqiwrAx9eJ9xpDe7vOvnwAMc9d7hzaqiEpktX0/UFLYgmzOTx/TyO4BL1X6tY39/DAPyWUaGIr
Yu54PB/aCq6wartr4BPGws+x6HfTbRBRsP2jyUKUoYhOxbhkGztRMorCi1Wp2VrUVUTvFF1APgEw
J9/f71WWyIuOSWcgwEC/T6eEf0J0N1NwjIpV2IDEd7gSHsAYFVQWYvBp7H/hI/euL5IAcPgnmUs8
a5T4x9I577gKaOr50oOEhh/BmHX3iU/l3jPbnRxg8qGzfTlfo2m/65hEsR6bd0wvN2EnXXboJXVA
fBCT0RBkwr4N8kfeTPpF0k/nD4gqPVCw531ZOUmnrX4q6TQ/DeI71UAXARFTxHsoxf2a2Pxkl1LX
mgtUdG49B50RKfDQK+FIQhAz3/MckqNM3Utdw4S4JB+jfmBTcI3OCvfCDUIUc5eFhsJzFfiXCAmH
YKuW1I2XYYN9AFAP2KcZo1YEHbqd1g9YLavzqeSrExg9xeE1QICM2U8Q9XUueyd+kM1yBNx2OZJ/
sWdDGtMCUy0HJR5CN9e1ejTBOB3eNQySMWxv1NGWVG7eETKpWjTArQGpoTmgf9O8oevrocjL3gDY
j0ufxWLPxFR82Kl7GA302BikurlLzlGJTXsEn66z5Ltx0le6RdmA3v4eqMrmex3+5Ks5bvU9+VwN
jopgXDtT53mjwExUqUD4To0X/be4/hB0IilbyZEUhkIk2fI4TPqKM7dpnlmHJRXzalB7uii950yn
6gsWQmgRWYa6MDDEJ1z23Zzn9LMoLELJtMol6F3Qaiw+JNtNN/jx86D6pd8G/dQcFBzV3J0FiFLz
95t3+sdHeAqYAS91cE5zj3UFSC1JtnlDc09MCg4GUf4rWEboBRfvdfl+QeZBBnK0v7i8lJSD17AN
2q/MutIfA9uqzlmU03gD7DqcGuphZCO3CIygTCExyzFi1PcTXYlAc7XDokBXHhjH8H5EJwnyOtlp
2RFDj43UpCkpWsdNPiZDKdMJcP6jmKhUgQt4XjHPb08EQ/iYoFHXQSvfIRYGJCjeOE6oBe5gLij1
9jVQ2AL82XUdfrHbZpNvyMl0DiyfwQFxYKfj6vqIy086TZIrf9UwrTle+S5rvc+mFLs8gpY5AY85
fkv/W67tt2xoe8Rio5JC4cle9vNbA/a2o9cGV/gbI7INtExZz8eM4gOaVPb/Jy97j51RQCHyKcVG
gK83Jz00jBVAGRBaZyC5rlQBYUNOmeHKi5sWCzsrHlE1Bmc24wFT+x8h20TEtLuKCS8nH9K4tWkP
6eukcxXMe4/UyLEMlCY1cz1jPkOryVyigAY40lwBtqi2NwAB+kxiOaUoln+tT5ZcbHMcp6EFpT+T
+jOs8bxCk/eH5Qwkuc89nqr8vuo/zzqcHwZL6aawgpzU22K0Nj7F8ou6sWZGwTtK5sUh04sz9IXa
s4E7f0/VKc5TdwTU/hKuQ75x5Qol0K7LDivcy5mWn760E3V7BjKICwshXQ/c4v0cSlVQpBs03NUW
Yj8tAj9dYeR+W1N83g/08r6cc8mr50UnPi64+m+mVfFSIH6USnZezb2EgpHbuzQY9eSK0V0Vl1AU
J8eN7RHnyXvMAn6+ATHbQrFwt2LeGSonN7ncdiinbDvIZrHRAHy7Qk1gvygwAOnO31l7HXeLnpqi
3ytcK/G4yV8ErVipTrEZG1dolBEBrHAT7JNc3TbLLNDaS7MIGApkMvL9L/3dUzIkgpwXCeWKGznT
Kj43FamhBRID0rRqgF/zAi/aEb2W1PoPghws+enxpz4qPtbCK0SWtRByI0J0RarWKbLMj44FSoXJ
8xaVWtJHGGnkxA83XCMgMwjy/kgs8Xb/dv1a66+El8EO7au3cnEBq6L72zPtqwZbvBXbqyiLQpDa
KGK94d7Spk+Omr2Qw1mx/v+YrQQhpwZN2RhKFbiUKqyfL6/X6q+wv9LYUAm0gnRwYfVqMP1cNZbi
wlbbx8zG4JRAlUiGwpW0eDttlpv/KQ3/TsQp906SF9J4JzMt2xFveEX6hgW/eqgRZ3ioaqZqC/7T
cVvfkUpC8YvYzfAGLq107Dezdj/ytkl281kSB6ZG3FKzgHMyBzDCO69sPVu6xeOBpZ8UArrxOLqh
VNwxpT2ADEUnrqXMhDwjM57oP4QtqWtzn1cX/cQUOtsDKAzTCDm5WM3F3USaesIuXsQJ2/85La7l
6ScNap/uGqFx9aoEM+dQzxb7DDYh5yRn8qwhXnvZISh7eOnn0TkkKB97cWWpRGDLM0NARV3w1LeS
ddH4MqrwKa2GmdZwmXXgF4NL9Ixgsf+4kOidGYLTV6JHEoB+ti7dcxLJ+UP2NW/yHrIyO0GlwqR/
6+704f1qd8jOlWlWUkhWlesElIEQ4pw4UB87bhZlp+s+BYhjP64fkRXkxNE8a9MVu6selXXOD1sR
3+ENlQ9YKqIJGLcJz3cgyPwgV9bQX3sUg3TtJ6+W0n0MTYOncEr0qLGlYyUwxwRPeCPbmHql/ONt
DOBZen0PpXb8Ai8EU5Bn+F9S4gKg2l36dTYKmEwvUc3FaOVWnNsVUzkvYPsrJJlu5+KUpupLV1Wj
U4T4nMoWuuXbhRRNuh7zLd8PcXaLu9XFXDklo9qWqJdKyT6rc761QtgtSYEQCk6sCMLW9p0Qkc8y
FiIecjQNeZxjtz1cysPo4U2jPQCyp+RfzDISpEzp/oicpt1zxv+RLrgymup2KY3Juv5pePZUc6Hu
Aak3HfPS8TYPuDKwqTfd4gTkenxJS8m0t/yfHPq7s5wiIH5t5RUGBHqfQXzOFH6Y2IMVly+CkasI
gm6K8Iw9vbNVfDABXv7Yle8VQJDLoHXwIZ1/gnXjhbWw8oo0rAFMYZ2sAz59NDzvWOiD4+8qIRzK
8lKQ0jJF5NK0wP0Ue8bu8UO7MYSOpI3nckc574WQboagCK/5jZ7mqgG289IwcZOitfPibXS8er+/
4L37B3TykH6Ojt5ARgxqMcBMnWe+VIYiBuy5LDGOMj66rJZf28c0k5ngfN5X+m9RvM31yfHg7FNZ
NWyPDWEOvHQjr8AhLXtEgRosywLnpqWqPIaP3bB9w5uqQnsrPEzcypfuNsXPU4YQrON4TScwuyeq
ly70NYlP89CCVQ9yjkxcClDn35UwkHeaadkjltWhNnL28kNmjgb1d1DUGwVcYKYJrYR15rf2H44L
COMUPreFRhkFDAN4hiA/hyW5BO0ABSuuHIi9ApljEZvvUpHoy0zpIHs4nImU5qpqG3/osgaCrTEk
0uhiQe3onYB/pnv5gvyizClLDMcx1brbfu0q1gv6P7B8k++gVOB1/9/5Vs6C5DRKyaJvkBX1urZ9
NYbE0sJ2iHSbOTYhS45aJWd7vdEJKFqN5bZPGsXF66zsmn8Q90dVbG6JT1axoQsFQELegzTOIPLA
z5eU+HeBmyYDlS4jc2eyoiRSoA9HgF+NAJZODWd4T1pmWKQo+aUfQhec7B7HFrOPlBo1taFjxS8k
ZVMBWZdhLepSwrLmZN3+7OjElHPb3iU4T4hxN3dD+AMsPCCLdXFf8rJozS4mVdA4oxBSdSMLQdpA
APNdI3WHM2wXM8n/XxhSx8+tyr/PNskPfnhcWStoW+djkbbNv0cG/YG9dHDXyKtmb/4Zxxl61/ld
X5Gs5FcfZ723TIdPCwvRLmg9h/goQsL/7wLkHyfisggqiFez9Zo3AiEi/7/zEGTfvs2l4l0z7wy+
GHPCcvjorw7XqJBWV8QPZLKjyvoXTIpOe/1pwvuS9CI5PEpcDYyZBYoUi9oRj7RKOyGO/3DLVtfC
gS88kqrhsAUyAugt+yLxaK27AiTP1chYhBCjxhGqUklbUASegsLrTu4uwmJ+8HjOlpCkNTLM7Qxg
e027CpjtGX5jaQ3fbq+dEUWKN2aCBWo/10CwToUncBtz82E9Hbab0MzEX+OXfinyWBkRCYLJf8OT
G6y45vsYUJI2lRkn2sCNEDKIjtKAoFCg4DSVetCKDdxQE2sVgjQY/q2ZO1uKP2HuWEzlMhY/hvwp
94eqolDJ6S/hdiABAxuth87q/B+DJY/ORyPmN2FJKIpTiLFkjHsMf9TTmDcvacrAsVMWH3trwwHZ
N2xOxqylfbO7ktKBeDDH4zEFBYIgmXGbsRaKJDzv2cnBOaZK306Jm3t5aUnfQpLiXbpQAMubFFGJ
HSonCzMwa/6Ck1OaoZ8cpRCyYe/hlYizWKca8cWBZq2CAAEdyrXEuNP7hP9Gv1fl3kPHg2RKDlkS
PDjUjepVZQB6YqMZFIG33/TwL5CBbulDXRIlE00z10dJFOAH226MgZszCRSekd1J8hOtDLdA/Qbu
RmhN1ZeMra2at51WDJ/6tZ+MEdLvVDwYMU4tQVCaoxirUSFQ9aG9cSmBTAeAFrw8c548s4zXKbX/
3GD4wZm1ui8ExcUv73oiJGd9El1GDWrMPQ+w/9EFNqKS0Gps2ILHCANKhJnQK8UzHtOQBddQG1lR
923tnB/bbCxYJNqOKIeMND8pyME038Yty9F5S4wqCqGiTE+hq4amuT77eYFgERTU3VSeYh0G5xaZ
N7/abikFmmzJ+YkI9i/zvRynRgcbDe5FBdbDKWnP0RPvy2oWDW/cckgUC7dhKoNRWpwmlnC48PzC
hHcvAEoica27DbKXpWkjrgPrHguzir/6cJNmMBeNez3Y9c54ote723oObf2DkKzJ7/ERkvWIDAxq
6KsqJnoqoOSyNs6Y1HxFY3jh2vUygL2DKpLGAgPAjyzQcPJGEUVO28kWQ6jhJuVT7KS+WmMUwhxE
odnNZODXCWTpIGkn67/O/YSr4zqE6KPhGbJetRyjgAjQsPkkMEm6zocd9yDLF0QZCtTUmI2l5rVu
J1/1BaQ3FhdwCjlBzduPZK4Z90N36Z8i4oh7TDJpJv0OZPhsUMz/XGaMXE8XCfBbfzLLpU35zw9R
Vr+jdhfLlx8WdPRrQHPSlxdr87/Wgi/t7LBJB0Z8OnIvXm+iJ/7TjtG3+gYZS64GDVt1CF9V3dWi
gADggK0/cGgGGih1lquAlO1lf4wXo2Q0apaN8+ty0NHs4ZtaiyeJQW/Oj7+Sm6dgdmMRO0U8kqu/
7T/dcqVearTWo6fWtmSGavej0uA90BKFj+wz1tqJ9TceaIvwMzTiO+g0hKoDxl+qlX4bdDtVbwkr
kiSRdq3KBN7xrkj6SsMjaFRjSzPpIuLA0NVwEj4CFck1n+BEijBRGXxh/LE0eNbyBZ1++2D9LkdA
2y7RYyLWdg0l45E7fnGXEl6eQADjYlmhrgup5Jks+3HQch+AsGt/LCi//fWttic5p9pvkU7fUTvf
bPwCPUksql9qSn0hCg/vmR0tfx7tSIagTljzqdBhQlzvSFPlcLXI54r3YALlGRVNkiP7ApAlnXHE
9vKU463bqKjdFARa/fNveMX4W7CvwAGw8u8L1m4kkowCTTzvOfRIQACm0uEz7Y1fROO1ZV1tp951
Cjr05xwU2VCQRCZuXwiReDQk2yjRRZcUCp+CiO5+M4V9AMDN6f0Yx4np2Y2vSOHlyiRvObhBRkhc
4Aa3WLL9369Reh5lyb/IP8YNlR3CXbZvDM8JD0vuhyocW4sPXnL3QwbZEKDNOU8C/8yJeLsXSMS8
FODyVA8/j0gOrV+NMqe8q/suPukdLyjVtj0ddgP6oD1jurefEMECNHck11i0GnXD8NehsgnrrmRL
klbk905l6nyz4yUVEZa65oaOvCH0GqNkHyumc8tftah0ZgsYVRgV7Y+nzjAw079+NIv/2xXHgvxT
1DTzUJjdsFM986znX++yaOsVqs5EHDFVNAsP6u/RJSxdy8Gl4RMRAwLrX+t2ZN/mZU3DiQ8jAVg7
X1Wg++gjBG1WPjssvCRtfBfIh6dRv8B6R5arBzK7TP2Ydq2RbJCaGwC0o0aKVaF/BFw161zhI5Ew
58tNsFLmxky0gheBuGm06+PehCQvUBOAqbXihJ6j/e612anr5ZTwwWbVKlyHBHqFoodkAl7wuS0z
uVTfoo6vcGLjoMuIIg5nBOo3G+0vmHq4/MdbhaIXtv6URCFXOL/lvxZuUqaKyVd5/Gad65ZN5BJ4
QUPh3PE7WBx5Q6TEeqHZN8ysLFZ650T60pVF7q00l1dD3VroKqzeFRdPVSu00txvc/F0nkhrqLJy
+TbhnlpzYplvrOOOrGLOZqheAwNgZ3koZiP0DYYbRVsPA8+icZzVXkJMCqWt3H6drgR+iJEfAQlB
p3JZdG8OjfTFnDi+51Vq4Ps/whuzcwhOqnwtiXkvDnIrcDV45LfXiLNTW7fyAKym4s7ObgsaNPV3
LdhSFmAa7e1Lpk7ZUjjFL3reUbFspaWnwg5L+cjPa5J3Vzn8HkOx+Zi2bd179fVexkBnPdJdigh2
V2VGKMGcS/BNDq8yJ40BoB1/V2RV10+t9ghbu45R5Pc8IyqREQ6dXN8x8j9sDFvy8lTPOw5ztcnK
t4n9XtELAVleaOLDHjkOlgSGFjp+X8gUNuZjKLadOWikroVhQN6smB1pnkvjtRDfuelvvi5bAbA0
PHp0fScPGMJuTUn8lATI2UhTaNtxznbl7TXluMMxEsircU8SOgBC+Y7yL0rZCTE7pRUWaINu3BOw
t8rNR7eVWe6U6mATZy0cVGWA7DrgfRkeKdaA1zGd3yUA1Qc6o0MBX1dX6AYcdxGIqfBvhxiDDvJH
nuhAReHMtaBtukNYrBX3VycrC9tYi6aO9TFbS7f8xXTGuNwb9Ka9XqX7xmmKVLtL/yLBCQAtBO58
+58S90aG+QBg3o9zdggCBgqu3DnrGpejaSyUG5VRccrcEDGH7GCAaiS7gXmIUq20kqXhezlFJ+Gd
+UUfLedC7WFB7gqIhybSbQbc8BHvIkhEmZp7CKecbjRGCxfaC7X9Sb+2TVU+G/xi3lD5Ki9I9nbE
CYIYmlOwR/f3aJOQR3rt1LuQwNP6GVzd7/qpqmye/C5xSq5Az/+xZwgiSS/BOSDfRPHmUsRpAwla
mobAST/sNjAPGIyuTrELmLv9JpeC4DcR/OCu/GGvjnRvAl90eKkmX39/2kHM18kCUuF15NRHZKxr
Ser3IqAnmL/CDX5ImCGv5ZQ+aCxsDHzwx/P+P6w5miy6QuWB1Hy1aii4rFq6USk+dSr0Tj21JfvO
q4aavapzLwoW59o8OpVncodu7E2p/TsLe2vpEPaksATRZwuwFG47qAnICM2d/y6TZ7xxbPcL6f1m
9A/pk6F9XEEtbnWKH9YnhahdqmB2SIW3tbN6SsCeFN6REvLaRCuiCGwtZS/dLY323p+kwaHN3j/d
5uncAObwzUPC9PDHnFHZ+Kh1mFMAUbMYoISxwYZZJxPYTGefhyBYaca/XVe4y2LhUeFPmDIM4XDt
BrH1whNLmxO3Arrlcoiv/Gguhbgv3wSlraNqU/NWk4ItqYCa154delpMUZaGyPKRpaPCleNLu7Je
kcoriWb8Y7VaQNQkSmfYkZt0gkffCf7pRHpWmtb3RfRy+W6UiQyHDKGpJZGY0citjIr7odYN7mAa
nMhu+bdMuBsMcBWwcui+yG1uingTfnODzYZKFa8Xk0l14icozVWwUliF93tHvLgzT76LTSUshuAq
GnlAF/msaOCnr4TSRHctf6mWTU1s8d7vdQf/2ZOuOyZG//EIikDEyXwsMYtFhJtzAt6spo7nbQyB
2RMl419IDXHq4lksVT8EcHC0bdAIJe3sfkz6B6JcUVnXEpnopXWb7GStGRJmWJAwc35U6mjNGiyS
tOml8CMQJ6cg1myNwqXUDoscIVXLmsvtg0K8NdSmTt7fnmliJFpCWGrK+C5bEAPtegHmjowo2547
sULTPy6gm5dqBtUHvTocvi1t6B8O2Ay1ZX1Sk5yGPcbX3diX3Kbukud2/Elw3XuHJOlT2SVlpvlf
YPCa+0tsTBU6Nw6Zl5k9e8gqyintmmV0uValBwLI2x+HUhEnEBOoD9OkiPJY8e+PVLA3f0NN2dJs
cS2g/G+0PzynPLNAvDURsAfZ1TDjAAQHW0CpPdC++ApMNdMdZ0mrsS0EPN46mhQ2UQhCMOvGR4pP
2QGR8r1YXyJ5vOWaArS4Uqcju4fmKA8i7kTZc8g0SpFRzEw9jnGm/zAY6QLFqzSSnfrakLjA4Z6c
pwmxOhVBP4BEx0tk2sP6pK5TOVO/gwyXNDLlJebSXgU9PIwjuBwBn47Tp/KW9Mbdx/PrMI01TYeG
Yklg1P/hLHjvXiLki+3wiLpKLM2tJsahcoGtz+mq17MKxGelNJHeWYtDsBC1ruYinKNQ+Bur4B1d
n1qAAyaR/QScw/vw488CSytn7WMAX1gIsemyfGCA2i7FKy/J3Yx5iCxBf254LK7XiL0fdMjGa9P9
YCi0HhT622TswQ1i5p0c55uiKuGV+VVtvWWrU8rNC1IL+kEe2e2xbZ0/gc7IcTn05l7kstpz/OnI
IoLPw16/gpyXz/WlFxN0igzzfp5vqjSxKbEwBNrjuNcMv02VZXsGwPe7ReOhdOoLNWD6v9i5Fhel
yW0evIcDvX3Un7JFq/ldfdlviQs2B1wzjZUx5Bo9AqDcK0/3t4ioT51ckPMFQH06NupmybDLZUoY
426e5QNCqwdGQ8dRTi/Cq4nlZS2ekGBLJg4N4n5lLp3LCXjiyrZgrnWabSah5mtqS+DUtviZ7vIP
mg5s/izANv0In/tMfNMfhaJSo69LMmOBKQRgDIynXh5Vs3mTqobZ4raG42zw+58q7W8UmeMaWYon
v5mh9ok6qImcvDGr8XKRZtD1jiAY8gMJqUTl0/8pDCgJiXAXcql4S6MVAZV5FqIZjT2CrA/8evBX
b4nmnHvHu/4VLzZkBBHtCkTiOyYn4zrQ8YEBVxNVaPvHwLRW8a5X9/RAXyygq1Bwm3SdHnn6PEdd
Lxlj6ZuS2OUpPMj9JoFcLtPVmc8+lv/LkCcUjx7Kg0Sjl9FAvgjKY7mFbBI2B0SKY8oXp/1wxwSh
O+cfhg3qxm0ehDFLtsN7eu27IGM+ppf2vY6XZox9Po75r2Avfl8frJZGGD2Y3cAvXOpaAaukq73d
+CcLu+eATW3ig0BN6kelc661Hi+UW7rTZgyHgfWEva92CWWdsberRg3xdm6m3OgZ6OOL3mmV+rzo
ILgj6UjT4gYNHozWHC6UrIoI+20ZpjJj985dAQkp2DuFS+WVcaHXsCMfj/gnINX65/mcq8kuZGkU
6fTHZeg4MJebZFQI4J4Ig4DBZ3sgPDJohGgxpt+CA1dOBnjQ8H2jsOj7D8vsPgx5gzDMVCnQC3gW
CF9E7f4soWBIgMtd9faukp0kPPykuCABn3tNMuq19waOR50L4Hra95RGqiGrL+UeHkgPlLw2BUka
yW6c7TD+sy4GmEY8V8shezGE/q7qUBlt+Gae3bQwot5ZoAyKD6aXDUplZeAqoCttKgDWKtwOAvAr
Dxru7J+p9FRU0e8aXxZ3Tp8LzRnyH1dgd9j7xK97JK1L7fLaTKl6lbXxpTJu3+JO/qmaji5cmFvd
RFC+Idj2oNKDI31gFAmz8kp6RKejvEgR4T+GlnSK3+v4vRW7dT8b9v4lolYzo+kWFQg/9XG3ICX/
r2Kife++kCvjS3EDQyh98o9I8tg3Uu9sbGr3qbzMt78MEJJ+lgXcU4Cq2p/W+C5n037ip4nqv+/X
FbDNziGaJpIURQUFHgk/GrSwszhH+xMCLsqH/vhs6j/zCf+QSqZ8PvJ0LqOBvBh9guz7SMo8qiHh
FdQpG8SFds1T70eTshL6pVdbr/dsDJF2Mwh2e9tiLljVjNLRjrlc6XdK4wTfkzmuEgT7JiI7T/P0
+taaMzVG4dF9y0iSvOzEFcYGKhTuBT+oPAPld7yUT/WrLdRfgq7kKEgUb/P/h7b/sXHdClXjh3k3
ihzPx34m/mYaIy0Av5tnubRiIPxg3dokK7N4/axw9SifJtZEgDSq7wnAYSrl7w0fYnRuZiMrraLD
ocuGXXE8xsowVKBOMM5baIUf4K8EOvtBv9S6owsnBQ+KaruPiFlqBLKEviWiPJ/fdlFmofj6Caoc
/aJx4nGghH1KSXjkA0IqTIFMGOMavpRPOPgL8EmuvOgHqF8CwGUkleDwWzjUqLNKXgJYfBAsr2UU
uelfclWAvoV36dM4DyA8A6fWWOEArhG0gu9aExce3xZAPkTRZgUaJon7cVkT3/uVi5UjXbtPLIIn
z6e5zQY6MD3/+SCn7S7gl8LEL5eBGMOLII5zTqk5OMgGDz9y8KrqFkKQBDfyuhMXJ2VvvBlPCQN3
uG61yg4my8c9unqahuQrSw/LMKuKZG0r32/y+ZGmWIADVdYWOfy/CkMH0jbXrZd0376e2VMZ/5gQ
kimc4P6aqnCc1UZEnBP0DpgC2ugXwb8kgRa6Cf2PVvxuHnWasZYXkuLyroXYmJz895aE62R3CTwK
W9QAymUQV9dS1lgFvQ0di40NxafNwwRDdEPZCwoGP/oZOuWHBrL9rdR7whocJyFaGdZfzShyt26G
NHKFErdoX0795cTIA7BMXMqXDCLDL8kGYrbr5ULjs7mmZovxMrikVw8/oWvtqaWN9oEJ3qnp5wSs
U1yzfHLFkstv+Utx5xcKdwD4DdVAEnMalTfZAi0+06QXJg7N5NKJ/1n8uRWUWR4RDLghEo3EUYL5
x/NRlda9l1uaCNaJ1e5nTnHLqHiYgFmedS8fUxnM5zszB7RzuejTv6To9PJ36P7sSqCOTp7E0iP8
ZqjX680sq7VsBFRseh8E9Jh18G4PZ/Mf9mb/Rak1ttx41Kia7tk7RGZ0zgdbsEOPrbuYsVJQkYtU
DFzN8a81+L/pwE62Eo0CxT6xJfiHT/2P+5wzAbGppISbh/1zZgJ15O8TTf9ilrhklbkkZ1/Utj8x
Ub3nsktAA2YWhUJ8INe2XK5CyY1wrgGffhsbcznOmzDAK4fsMz0379h7wZWzdsK0NY34ULQlCob9
SjGyCbueyK9mlfepSj/O48OTp86NCBdCJmDLd4hcBC6AtqbEk9nfXPi54oke7D1sPao3AnnM5M2B
eJvbdNRPSIGErubBo9FwsPO5TLfOKtfS4gC8dE3V3UquJW+v95MXzAa/9UNI3t/uakjCBCXUR4+7
JHrLTS4ListiISQEXqt7HgNJ4dG6uaN04n4FZRlhp8ZlOsb0ChCvazRMzpS2+okOJliQOy/827iI
pr4HDo5ZurmUCSSeRAGDfSRAv66BUmHOfGsYPWrCV5ahVBzSOUCVBLulBNyeCr7BnfCtK9oENULf
JXTz1uqWO6/tIeLamvWcmvOnEiS6JrOpO1OH7CgUZiWkzqsUe1E5evC4+27/NHg6ET9XwBEI35tA
IjvpRJ9Q7+pFK8EB3VfdUV17sLfR2j0BsEzB3UEdXM2zZhOixYuc32rSUlZujU90/tVYsq2pZ7MO
gZEqcgYsQ1DTuucEh9f7+SsyOC8qDgI51nPKnFRdCtm7AjwOWSMb3yLCmXa4ZX1AwgdJBFg3t5GJ
5XPxo5Ss+Vabrnqe3TMmJ1kYIwzmKtx2fQe0oLBL9HoY5KAJpM/asSikA9HYjMBYFOl/Rjh2TDqw
YjJfGyELERuRz34xsTxbsv0Wv7Jt5n6fDjA9cqq8VewS6fDAucNistTCWh97nfSCDDAq54dF6bdu
MyWGIS/3hk2+kOTs2OxysWZXOkto/od7JL4Jva0K2ImIn67wDYXxVIH8yao/GiVg9sJdHGwebz2p
zJjhN5a1b1TUdhQ/dExLy7K2t2+zYTWEuZKDnJMgLdFs8zxUS3nFmpJVjXbHJTnhkT8vqRRvIRUG
5SOQ3o9yhPsfdMuISCwIHRbRYgtH1tmzlLG1CCKlnBY2U6YyQu0wDfUGURkQn1hamphznwH0BxQ7
MH9oI0Qw0haLusZpjcG71zMhhX8mgk+usnqLEdRBZXoorrlD5VORdx7dLe6wYs6XVQSYlQROK6O4
QR2PaxudRJ9CSlTG+JpaiZ7XFy4+3Zekpj2vZPqIr+R1QgyZICcOp8XgLDD386Q5wKC5FCa8J1kM
JAUUc511mnRgu44i27G4nOUQfDfGMPvb4Ok0ryJEXWdtXOd2bWnW4jvS63S1QOxGvjP3YYYW9eUs
TnvLE1CoMj38JG5Nz97VnzJCfLUBFRL0RyLQoWaFmel6aPPLGRKckIEzMqZVVpj/9709yajL1K3j
McWr64tvfyU5hPIPAJy8iiRYWldbBFiEl+/flOUNIvx12ZLS5cpkHI06D728DHOPQa4bMTv+eeJI
MD4QZEZCnsVzb15ai8vMZsSXON/+nCZcjmIukYYaZ/ovm5Rj1UsR3c0PVZ9mA1iK5AyimK386W5m
7f8ABF1ZSkGt36GARX95F/ErU0JDEy5M1W2l12qB1gHT3xzDek5gxXh4HuwBlsvpo6r2lqR0e/GO
LQYn6Abkrz/iQ3l2I4LPJV8UJK4e7XiENkdikbc2GzcjDJ8JYTRqDJLGjueQm1/WMBa4jM8/eNkF
Qc4LIb7L13iNgzmhYXfxmJE+vD6mHxgh42mwc6tfcJ/hjMhuB0oc7i29uIG4xKxhZAjAB3LhIWQb
ALL4oTGZtjBJ3q+9JY+Yi5u92BCCX+2iCbtugnfR1cOF6P8uO6mbjvL12i25/ewTSFuzrZJAPqby
0vvfWGresAOJocEBFPTKaf5uSrS1gqKQ1A9C0VVHrDL4T2x4FCMALustARcq54Dp5OApUQco6gxx
zYexZGdukiCtjozw6kkvSbK471E3v7KgevQolGszPR/YyytTBr5bRWL+DV4xhoGeIpUkWEYSbEzx
HSDcEPzxLIDF3JK4beW14j4REH4mNLEUqqsLxWwYF69kkpvJJhGEeW9e1unPC0IucH7yKPzB8L7T
ThBhCVr7id8RZtdjYwAWNv/1S+3DR9GEArcbriWsbH3VFn0Tnvo4ZdWYZa4wEK3arb0BatahPKqV
vUkx0OYAJCai8s1uezqlni0WQKvjoFC8DWzt61Z7FSTATkRv4guESA/4YyHltajI0RO5v4YxcyCx
0BOQpaUt3Mx1UFUQ1jVvcVKdFNjWT6m38uB1Xk+o3Yok863omBN+SqlXfxIGivsCubkitmhgru6S
R2Fs1S4vDuoSUgC+mIGUe+Z7Hb1XIYIxW4PXvUwJ/CE+sfiDjcqcskaUzeOf1j3gKVBf8pDM04Tw
URvsIUNVvx+HUGjtF/7cvRRo2H1a3W2heJpCC98XjR3LjufeyPYVkrTmuAcxg9/qXWDV1usQl9qt
CGbmTvYiGx6KiZd79WcvY0h68mIOzFYY28vCvzpASyT1xfQ95xq5R2O11Y5Gg1iyYC9xjBlM2W6s
yRjT+mC6GVK99ecwwpUqBQYG7S90NAmdEc3yrP8fpMZqkEfoVzjbPW6NOo+vhu4+efBfKK+YCHCI
6wy/cgnBBGYp0J1U7QglVcJVm9wYWNYzjn91JYrb0m6W+iv36u4e37pqMHTRA//n+BsjlovYYos2
nZVjCGHaBnltXi8w9NYDdm0xmTRgeEnbkfVoR7s3h5hijzZ1A0++pzt2LFWwE1aLCFLo0AzTmq2Y
jTq7Yk9+gdHxosgT9yI9iiyTK3BlVUIlgHj7Dix7E7+XDZEg3kXyMOJmHSC/o2pfEYmU11bJklDd
fe5MC/G8GE237UHvf6lQBXsG51DHqJ+DoErVz2UQbuQH9SfwJKUONIV1Yw1pEwFgoICJccic5JDA
a98JIuceZ7yHObfVpTj315q3hrwqQWC59MuvhloJSz6A9BzFbS9JQzNK+3HgFPNHISjnrW32DsJC
53jpgTtQ8c1aP2ZPgsUCERxTjwEXVzUosgMijYk1SEyjQYyCu+l+O6vuci9reb9J1FdDznWjMoZu
RIOCFTpCaCyzYfw5wKu8f3av3h0mSJx3Oas6FkD5DHlWx6sFB7pnFXxnIBF/ffLZUSDgaQZ/5Z2H
J+zswe6OllcKr8fF6Xk2i9CwzC9zTHC6a5Eii2NLborZjIih4925fD4DPTyUaO9t9Qma1q9Q2KLg
hFSI8O39MHDu0jpMf+vSWBTnqs1DS4eNW9pKxrxJ7N5grGvgTVLKM02D0SWqGJ93UZq03nuDxKk8
IT7jTRaHfwjIodFQe/Yh4eKiqLoWkFYsVE7x1oMy+fS2cEf94sgOM+v2UXlGYIjl6oh5ezNJzuEo
OqRJZAu6VwYFZ1JnP5fFr2ub5+iBZjr4namawCCdRhcpMxhASn3YHHD4bLsaAhRqh0/tvHQxGv1L
TiY2WREGqGPtAOVD8RqKTW+WKKiGnLBybNkIebHD4hl39C67aotDbcqRboIWDikchs5Ap3WzAXV1
490NaOgpTlHHGSvuyGEdLPOrqExrUYmFkv1Xr5Jjj4ZCuVhbT+oCfXjesIQjdQJptJAUXlivgVgs
nVQmC0Iu7SeTKSe+6S6U4cyBEbG+ygLhkk5FlXjgwG8ceH5Jrmp3/DsCLMnjZJlknNS/NjKuLVVl
YMEc/uOeP3GDjRr9hKd4T14p6tHK58FWi97tyg+ZHfxzdJk2aHODwo4zWLOKfeCsqk7hlAmAhmA3
8MmX+0MamqHQUyTJb6oRROJxuDL1vyjM8NuHs+Dlj386vIu/GyKONdOldP1XqCLdDgDW13m9Lm4Q
pKucV01H7HP9AwHeGOnRbUUwtk1UkZ2WHDArhkA3vlEEH2jKz7ITWrlIYPEs6PNvbZLKFiWeJxQe
Q+VHTnmd6BkhquFOeObm+EpBJXe2viHp39nw8d9BTkUUerruqaYPaBIDTBpeLnbU8toiwUzJTTyx
pbp9z5ScyNr/Z+90sPGdtcgPTtqrIHfJL1DAhfeyokPGh56FqcNCa2DPR0tFvgYr6PjRH66SXVDA
eZnv+wQIysb7DunJ9um5Hc6pysajZRcgrbiO+yuz4xpatV34LogM2tUSvZCSyatP1NnUXojxcPjG
mRR17toO35GU4nNwbDxvT/lyJsad61jw1oInlkYOv0parXx2IkPlBzSBqz4mFznZeXcoSVv9rFDk
C4vaUfa/a7Er9YsCfQxPDVOviiBbydimDoeW+ehkHeeu6Gzds/8BC2TFjzvd2ysvVWYxV9f9YDJb
UKYmedzdllONoU7G0KUEl0vmiL5ayyAjLEQAynb1FhUkvq/OgfTmLptFe91B7PRjCGutHu950G+C
DCXDRnf9PXBkQStkp5GvpwYIhccCrw+SWibPg1ABkJvkAUdYTmNO92ZzZQjiz2BmRceorVLJoaGd
FuJPVkmmnK2Uf7vOumHdEbCf3fvXOGzclrjJY4dE+uvntOUaoMbHQtk7nRgpSg5m2iy3VPkLdtKC
MbZPDqMGLkLxfZ/1b42zlxAf5MqPOnCDrH+YUd0MqzesYkAObjYESR+XtSTuirraC/SY30Yj7q+v
y7x2lq8hmedRC8MlBqUKzZKz3ARSuf0kNao1R+xUsSVoeq7ldMYzk8+mT0zVRiqW1+xlpwblS1Zg
qZkXNIGuulVz7k2aEP9Hg2QNPckJj+RaUjinctFMT5vGqQRBXrfXTW5KUZF5cYelSavyIO/z28g5
D8p9B5ZhkBOkrheIbz8GYjdY01Tokd3gQRsJQ1IyBe4eBe+qcc2A8ze4dOgpky+BCFSw+X76sJQZ
03/P91ZEJgClb/cyJtEqY/47klusvpe3/l9ScnhvfpFwsNmtlHE8UHHDb+iFR4pyIrOv3nEXCItt
rHC/HFdp77luCJgtCt0Lpwv1c+i2K0I26FV/rnJ03AYg4PlbWBwyJLz2ZB8y9F0B4XGUU4aAMJqE
ExLd1aoX0sY2S5oc/6y4ajI5JR+cdLH1IiuGhJSH8RAAoe6v36i2oWeAhfhrvuF2bNDGA7PYFCSo
iVfHU3MPguoejfZo9wi3uVD/K4difJTuI2qb+tdu40Ktx/97/1ew8U2XayBo3rAYDbHpDHrCy6Wb
Y3oEMPDAJZgf/DtX6KLxiNggRlR8Twvm22B0dnt70tNB90VlgQrlm1C6TEudFFbA9vpAIQYLCphP
j8JK0jr0WUsTyWbah/vjUYZ0NnGO6Sv9hvip6m8e8d9WyMS1cYrSgnbe9/KQaL4LepkgSTYperPL
dKlJKn298doZ/AXKMwdli64vzNf2SNkIg3+Q2KBfSC4swwXXn2QtgrSo7RroQdj9LFO6sW93xrRT
OCIcRu5vLHORoqZpUj1fEcPeteKQ9oWN3qQf5Xd0m1h+0qXahdU9+ZWnjOCN/KTV1Qn2j+8MJKCv
3PzH70FEi+9wRD+UmVu43bwTLaPaP1KJxP/1ik3s45N1DekLBnYJqHl0YyCkpo3RNjWlWURv7/d+
NByyfqvgwmSR2p3le/nxOe0okQAiptg2PqorDYNOtB8f8jY2d756cKpPXKNPW++Cqr+C/rdiIz/W
3W9lmzyQhb30Bcki5c8QLndCgKjsJlaSRZTbIovjbmhDVpe3G+R+eNDP9gfZGpoReX/2nQYwRteJ
zbU0HtWPsNu/euG6cxEfg3TM3Pac4H6dP0HdqY3D8X7xXjtSehWn1Vr4SJAHeS1LcbvbjCJQRuhv
bf3sERx9hd1nNhl1gSTUu/HuPS03Tl1XYUj11Z1nYCXZpDHknSYuoqsMoRUOdDNRr96bVvxe+eHw
+3eWVgvKWzL2gXXQxrvJD09nttyduHy+QFV4GZ5SRwqbAMxt9YG2CoxeCYZpmCnh9HUm7lX3q6WZ
KYIYvcaLfWnnvS+YshgKaizEhd92AN6FRfULMRBIhZoA3Bl/+xMYpaZSTD4uTv9/J3JDBxzG8yG3
YeqdKhEIlFlt1fV1H/aFlXkET9PENnFhHPNF4eCnqj4E4ya5Th/TIMgif2QN8csovloPiN43F8jh
CAmS0t8qHXHKE0y6vtVyevqGIClZXDUDPgVophEF/suKWH4XU3cMCrPT4PneqVYL6Yxh6HGiL6xi
tqm98RY6qSXLzNFe5WF8hTXf+HTQevjyaSYz9b4yXK/fa4SuU8Vgrcfu6m5CTif51vnN6PG0BBsC
Z06bvPN15/+upJy0XagiBUpPwF3IKD+aBS/6X9AIsvtvJHFqTky034qbc/QYc6ynwuPdLqPthAJt
rFxWcbjMoJig2GGqE3BPFdHZvfc/gsaCXKLoObNTDMfwdeTN219iBhrdegaX5tjPTTuGxrvpE6Ra
2gyZnqbs1M5tZe6onftcwkWUIpIBGsX2m23kAQYtmRedkymdzdY+SvTXOEEP+QvHp4yivKDClsQQ
nCbLOXycgo67WaqgJtXre/ZOu8Qo09I/MN1iy+PrOLpMqs5TVoWVOdlnQzexfFYfp0pguht96oKi
9eIVPU5UjttcEtmSSnWt0feVtsziDS0bbS6Ao0ONNDjQqRqOag7cuuS/WNkjX5jlWi5EFeIE/YWG
Gd1CbUZ3WEw+jcJyjt+vQSlfemObfsLlxrLgZBhMKoujJeFKUWZzbSPrcAuSD1re+EiPvCkLYHoy
dzoUSvl4XHYd7UP7PzdBkG2yOLck4/MIx3XmvgEwOG0zcYmgbljr+LmT9pUep8xzujCQ4B/Ce3w3
bM4zww6bxGlFKhHoGiGcZSHOkoFLgnelXPcTmFpeB0g9SXSqeNKjYNGULvcn/uM6LR1mkr82v6T6
JXuCtRroTQhre+MrzewxynMZ0nOUFdDcaT9l6Q51XTNqicKQWbU867d0mjDSAqAusJfGkcj4kn0E
qpGD2sGSly0H8piJgP4Fw/hLVu3iZj176aC90dwI1xlRXdsvUg64Z9DgweayYf8qH8wT7x1LovPI
Y8QKX9OXCm/44MTVjMOQSDOSJ1DmiKYh5JFx6HvhvjoXgJFDAO2nWjsCgRnuVthI7ngwjyBDqzXZ
hK2gDfYxD+p5+EuFkmziejrfZkaxIaYwJ/0aZuW7n59+0DqU2edBqALikdaX588mtBA5+If+R2o2
IF0CeilI9bprcEPoy/ulmvdisk2EsK+klVt0L7yN/5PYt6AzpryybqiDZexDNbY/mfROlIjp49KI
XXlSDtPlT5GhPY89I/dpJDSS6r73xCc9vj+vmamkYVr0/GwJSJTNHDIl3Km+bl6adH/own1jDhVG
3BTGj499Jhg6xqgnzoJr0uCfHp/io637dwije003Y2DzucK10m3Ximc3vZN0SSdDE1LkGjMvL5of
vkY+a/S9wZOVXS+Q4djY9JWws+NmjkPtE+0xPxFfb37sm/7KyUOFhBufaCaoRKHVX+aBXTMaMsaZ
AncKZCAgah4nKxe6BjY5mTQtpAz5azhYW3b96XU1GsMGCwx5JZMKQnJP56qbPzVGeeNKf3JtnuVZ
Finr536Vhfk9V743FJNNwAdCzs/VG/OW/pTr9uiJqvLxUdtgKhQ4DhsDoGIbzwJmVWVy1pijckNR
aqaWc5FQdd//xLCAIqgP6fRM0pZZqrvmruKlyq5Jzg5kIq9qk5veR7WGwvEXhfEW+VvarpF04qJf
ValFNyvjbZ7FYhvQ93FRlAS7Lqz1+G7VJc59teO8pheRoJM7Br2G+SKl/vk2cuFtHah4FaI3cFgy
CU0nn72TJiaPJ6op5gbMt4bdL4B/qSWKs+w6xKhgSwhhA4ZmU5X659Ibw0fl3M7QAanT6w45NUu6
EcmKpK38a8xXP0YAdfdcDCxDBu12HNBqpNpdRvnF5CVglUh4MuHGkJUcWh8WTjpxg6vIynfLwWNe
I2F61sYxSRMWM6DVXFOT3dY6vbYcqnG8ceAG5BFQ+RtatSWC1GUMVU0vlrZukAAjmlXNplgZfJ1p
VkIqftJD6EZpqrtm3aLUSqWnwIsOLMKSANwoQBpKYwQ+ZVeY55q1FY2ZkqUjwB4PbDOVViy2cxYc
DX0111A3JbvypBZHjyXhRA21Oqyuj3UNuIe6vN2dW9SyI/PjUL60KNYGOxheamqtMI5+1I6Tsfs4
GzLvi+Z0X19hBNAblk/ONFXTjDKBPlg11bXuapv+dnWKVbJ7hWOp3g0d0YeloSQtDMENFFEQzgtg
xZjsYNq7jkWpVFh2NWWBDFaRV15jXojPc5H8GpEJ1YbZfLUoPj2LFGinRB1tGJLAUBVFo/sDBxP/
n6Dp3X/urcocCh4ahfvFu/l0HKl0Lj0lj9dt/50zkOISQoAmYtroA5gOS4Gw3lsDXHc/Hd52IdN9
xv27leDwHbrNGEoIGnzZbl9OOu6IMLDIkrbWknm0m4AWBHZk3A0H4EltfJUpiOPiRCOIgJMHRLTd
MZ9Xy6/9nlWXBT99I/t2xQS/UMb5M4P6CxfZWwXYRZjdgJOQngy/KAG9SAHan3VegwJ8amZ9lmXQ
eyhifsTORhg5JkNQzN8/05vIPEbwblLzjwgkxYMF5asnHtDSuU68jFf8+DAL2MiZehWteVZ4mLkI
76zDUmU0B/q03CgRRxiqAGkUuouprDSObq+RuRrf2G/Nhd++kMoR+uKa5cX61JLN2ytqjNU+pkuz
sRhir6M0VJO/1cPGbU0UdG9o7QaCAx/ROprz8OsxQ+LUN/Y9Xu8M1SfJnSIjCIuCXlMDKMrJYqmd
iA86EqZaO+h0FhiCDPyVTEJRCMIgl1iSzQvvwg0WWweURbOFZiYatqR59CUSiq30GtraT/2wkGEB
hWIoRh8784gAgVZBSrDZ7PUceRy3rvPYizFqXToX9zDpPGyZQusWGbmRlxqgFUHOpB98tNUEQdDD
vDKeU/tChXnAdLdmSbehcz7+PBUvCbr0OFi+hEZCP3geVtYFavpj9kgcJG+z9pOsImLKDGobuYP4
fRt0SQ6uw/Kh2wJ010bnDq3pdM1cbj9DckxpCOZ8WlhifV94vUUUOUPe/mFuUOrX7uZfJOZwSBl2
xsMDOOtTeomI4z9Y7DeK7zOScfO0XDn+Wdw5G4BIVoOcn0JTTFdoQFGtYM8aDC1wI7290qvnqssw
kSOwZzymX0/srjtO4upMvx3vKfEBxA03Mz3R/wFtvAVoEsQ1UTU799Bt1TP4mNKNweJcAmxTs4ge
AjjnfJ/E+ZsDZgR6PAKurXvTMxi0+FYkoqM2ZR/1jIan0kuxDxs0ESFY/viaW6+cSquIu8J/Fcpx
WsVMC7UuTgHo/0wcZhv4WsjAdXYBDleu4Gg2k+/hgotyEneeWT2fU8M2J9XsOLnZBG8n61ylH6k7
rkMGrYsMJqP9H/Aull3ipHuE4dUiSnOudRwb9zmN2nCFWWHOb4yJJBssXY4kFwAY2nfJYJ0oLlja
jw3BOI1SodfbGplL4wdz8/ntmebMN0N3nlseQ5ZdhqFgCoSOjFR4ga2qkmmG/ep7fuhD48YbzVlJ
8RsVXuY70CjYx9W2MQCg+QYGg7SSiLDx+sKhqh//oNdnawqZDWssZZLDru5/e3v3crymN1IsDroL
G/vgBg0T+5TdXxIL7XrtaQhGYS2kXHujb3ouaWbbh0XxMaukx8Mvs/G1/Se/3mBEBByYbKqQ1xNJ
kJ0ae/hFCah3cVVRYF+oMZ0XLTrLMnXqdZ+zMXzQjyXIH+oLpIhSBq4eltMXRI2dIdRFy944cFzB
h+nnN/FU1PqD0dmkmPXuXtY+/YoaJy5THVtqiaPscDvQH/Lom0T0vg9c2yaSQCw+y0AsPeIYr/kt
+UawDYS+fYbc8JGFuRoYYx3Dm+mDmS80OVReFX3lk95v3CxJqm7T8Vhj9Zig7nlY5dq9GryyZrGq
Y27swWTp8J6Vezrz7YBL+Yw9fdIO+WWbvNKwXMp8eM9zTej4K9ccVGdLZK4WvwPRBne7d2FWd0uJ
tNfvTw5Q8wRyeGnrKb54cMU4fv00QQXs1EZNq545l++XPIFHnOKr8KY32mxx9k+QPuSFGP+efskC
38452pVV/aBRDLcoVa49yD1P9iQDtJc+A3N38xWQ2mk++t8p57E7EV4ajYUhT3AAUAvfi45wXWSP
3yDXk7LmMs8yz0K6oVdCO1z4RjDXJNQMggMx1n9AUnRGpxqA8AoK1RGwFa5qMvTdaVuklzhhH0wi
6JeHsG6clE4NUv8SotJqmIjPRy4Qbv/daHp+seVMeqMuTjW/VVu0B+gxv2/LXgVBdvE32onjT06n
AhEXhe1BH8QAlERKt2/RaRHN+kRrXeyWvSkQQRp+lvi5AX4OLdsF/nCmmdoHYQkRzZjuBOfcnSVJ
DYftwCqA3+B7v7cD3vM3RjA7hopGKEa7kjjih7LVhGgJIERqNHfUWus7RnxGFcwBns7ncwmGlggt
gLgq5P+c2C7fLPs/fz66UiyCTk35/BPMgxD+9Cz8ZqZivT+fa7U4JEqGNWWzDgo0AlFYgUk4+4Vp
cgJZJGL7ovOuhx3ktZ3UN+2nWL4axlyqZJ8NiT5vGoVfMeq7wpJMfYGb/RXFjhM8BlBF0uvRUdx+
nfo87bakuYH4nixX3QWsaoAxodmN5GeH7oYfusY2tltvU7YTmWE+cyvMT8Hs0KxpGcZhZ5QrOZKi
EaSGVmIG34wIGIOJ0dctOXctbSKePf3C2kvSIv4WzBkFAmh3SfPBJH60rBPPPHuBWaZX4PFeopHh
9diHlgHL1CvjmFBYIIQswegtdZF6I+bQ6SIV09FuhNEuTnnAtxbZiu5E7Js/6UtAVDMHSv36tfrA
1p4/gunNIqposSxHgni+uZe2VgbPcVKbXZ9J6TowlQtyBjvr30v2LGEEssKxf/QDrwO+hoDSHTCp
3yMZLmx9zeu+0wBHBestxz6Yk1rnrMFqLCqynxwErrahrLxDRIXi300zvUD6hFnSJZPnB1lVv4sp
5yCaZnNue1T8ph71exb7zqwShog8r38Z9VZFj8HJWZRLVJOrDpl8Desw4zQxBrtohBERtQN5w4at
XqtciO7CrY3PvYe0EN2968i/uBrxdHdNcIxcgWOW1+FFxTiGBFWniEbZyTEpuM53qsubvDKa+AWF
aAtfCc7JqDcdjo4Qkm71F3yjH4ywLHTDlB9AeCorR9s0MEulzc9CLTU5Mcph5+OoNoFrWwwiUVni
DUnjdKsFCziFYYBmvjfpvQFjFdoXFZuoIlQ7Ej+SqWqiwESikna1wLmdxWbNcLCVbRLz02N4KZ+/
6LMLfTOnfVlFF8REazaPb55YReGAwZ7OXzugaXpQd7QaUq7Yq2xy5XfLX5bTdRNI7My9T3c7Pitl
D+B17YGVM7C4rq42zMpIcLixORp+IUgJ8gEtiX3dmkUoma7oO8HHGw1gzFtkc/dUJ2Xga+gWJSKz
Pky5L33wOHCeafGE2F95gX0J+ynwttktmSt/b6dFgVpmCXmjtepcEODEtcOxom4ui3vAIggst33Q
cjNjWraGhqSFpMSMT2vGp6iJmnDhPv4e6SvOHohD45+6rrNXGAuMeF7lmGOPJ+KqtjYxhK+NFHbf
sfrWmm3qbrdZEL6ez6JOmlPv0xz2XvZxO6RhMKXlbJE8YNB+ztRNmrJTDmsG6rWcplWtZW7ejtMV
s/oo1xqjSUo2iyBHFY/ROmy1ZCirpRYZdCyXeAHhtw9uUPAOzG36rgFzUPN1n50OEHt+uDLd4qNB
QyKP0NLT+52EJEuR4d/O3Z7mJX+EjNG3oPeb9/dG2eL7TWfpAj8yp1K/mjRRRTxW594LJkzUyNdI
yHzaaVOCe+hNpLbUd/17O8z4osQqZfd4rPWP1O8LUG6B4fVOEEiNwT2FSEZ0EurEv41xvRI7ZpTC
o2swQzKbTyYXce14xIJiNME0fVeG8TulzpS/rpVYZT/eJbq3FBm22nNxapnDv5G/YGSqVeAKbITG
kWhHOV7NRUNZhQlU+4svDM8WwNEB4fYg7JF4zLC0pRF7cq0sHHt1Dc3RLPBXUXHmcVO2QE4JfXH0
HvPDm5r8HqeyDs0VnrO+TPwEUZ0ne5BNubIH9uWPbGOA5wbdEu1FO21+8aEeNAngiMQVA6Bv/1pu
JTLCcnF5qQipmxXRPgRI7pQCaUuQfq8iQvdQ5i++0mRXDceWjJjGHgwLz/HHvET2+lko8krQhBuU
yiquozwcZdT9yJaRBmVKMeTnP4/BAngsxA70Shp3lWbfOlsFSnRAr27cOc4BVQAcPN1l9HaD7DQs
aIBrt4SXCcStfXSJWvFpXoSeP5DbyehSUDUK1BqrlIx0FdGVWMBHEAsOa8d0s+3d0OnEPQiGNM7q
cIp239dKLFYUYEBrGQ2TjJtVPeSHaSjkXBQk6M9uIr7ET+tpnb8B1OAY8UI8reoHXSFpfbGauaEc
WhodS5/twMlsdY7rk8ONg0wFsNOjKD4GU9oQsrDflfFnYMbzM4bxVgUIObNzTvgQFFwxBAPyGDWm
IL6Sqw+p8FAFgITNa2hn3hiUUmTAKwVG8FGjyma+BpvrDnxlc4VVy7EqVyd8xprHQ28cH7SK5LBi
6XFfjU4gkfl9SaC4Z491wSC4dL1yADweSFdQNHGb7y4gnoxF1OHzhIjFJhfPw0w4p+bBoT2qypGk
006x6wXMsy0iWa+6O7AIoKf8EH0NTKNaLBIH9jwG9SVB9LMQhllBX3iKVBYIpXtH1R/ipnBTbrAn
F+0z5gOuf9/5mySuwoA6yAxclTAO9NqKSj0LZciH3I9+DysVyQs/6DZWOG0mQz5Mxq8A10LYm0hV
jURHnzoc0yF4zPuh7iK/NoZRUtlPQRtx/mhtaXzszQdLNTO7TcDcvSnnewsoRooWM1UIJqVU8Xds
MDpPzA2D20q/ugeXxJsbJtC63NJIlgmf7H6f9Q1F/bsxJsfV2X96rSHOCN8Z3QXl0frac44jstf+
zyUoadg93u8blZzWFq2dQBYAuWCqLCc5cCJQvqg+/BaWncWlQi8lb/hTAHSEXs0wqzOSal5C79R9
S5HIEIeRc5tqQ9oxIyUWAau+WOktIiANUseuy4f766GUbPpbsjmknDngfeQtLxMy4wx109L03awQ
mCebYUArhdJqTxG4Wgy0QxCHmQok+7NzuL9mxjx3Wdkk0oPRRHOlwQ6b38gQTTzovZz9gPeQVVBt
3uzxvKyWTgzTnFTgs0DK1cOS6kz+PDqwtOBb89bYQnt3lNnpMU7UTrqAqOOMJBHDZiwxvRJ7O426
WtmiFpN0Y3B4wY9gzMrbHda2d8KhnzryS15v3NcGDgVpMDCBzEmjeAsbdjkj5apiRuF0QEbRQiZy
tKx+PKaF9SQ51ToNylXW4RjPcnklrnSwoj4Qww4uzIv3wggmmO37SKhV71P3UvKZDuO3dg4yF/lO
eQ2JjR7Hos06xTjxT5Puuz0XRFQjNYRTKiYfi4zc6WIcDjh8ZOwohesLQ2kC05bkNeP6JRR+1r+s
4a4GkUGDojGfQW53ZKELsTdBBftiOxWmpvZ6yCiD5vY3nxZOvo8cKiQYjb+foqgGrILhkEP7IgVT
GQSmnykTmUcJZZYrPLpKtAummVldPxgIX2xKVTjP+7l0EUhUtHtT1w9B7WLqGeD7UI9HZwp+IeUi
VM7hwy9cnxqpFy+0/NeOfYccnVV5cHQXyTgDvm1vZgPNuIOPJtZvLM77h5i4/etHw3ZZlxhm+oBK
XQmRGsWCLWQpA8OBcmCQJMEjAWQ5hiBLNyUjc8VGOfUksbZf8ZA/QdAHNCDVmsXnr7Y3VU2RXSTw
tDpCfGhkgcTjqiYazNxQvzcnBE0dsEBEqzgKGFMem2p+E5IQEt2AuHUFsDJFRvQgNwCvD8tkGFYc
ZNaCpTD0cRYWs6Ga0tYwgT2QvtroNTF8vjV4U52etzSYLUqInX4ZsoN21fBJyx1UovQa6lqBw5Mn
3iOuI5vIquiTcGfl7+JEyC1t88F3a26G9ldAcOTQ5I9xfGUWwsH6O6T4m8ODEKQ56+518Xco4Yzr
rIsJE/OB3Hn+afeiw/YjkZzTh59WTmSsU74XiG2eLlU+kWPVRn33+9/HKMbFreX+CgXoolZ15wM9
EGVF3vXUnqd+Ub76w7BnrKcYj6hEqoTwB/QcJezQ/H2nsbBnBf6hLw51j8slaNWsL3Gp0a+0A10P
HuHIQGmQ1B6P+NmDGFMK+KJV1F+aL7AUVauds10j9Wz/sSAYp4jt2IVtivoHmB71EBPx4ER8HofZ
5yKnmU4pfeumgJveppJn0vA6Hu+DBahutnFEVvrvKO5W5Fy0hwafsfeINxvhEoU9wSx3Km66ocpu
CrlhC1R4ah19ePiXbp/mMV+DOsG5+PAlbLm2yrC3RUrTFsFzqYhh4E+qaZdg3PV1h+PFv7gww4JS
ZaTr1vF454P0EGY5HRBwSTL/YvSs4zEOXODtU9a4IP/z5o+8znWifTEwWI341fvUxp6a+7+acZtV
vxuZ2foQYDI9X5E65pq/8Kx5BRe1qOzWKDXM4zGLS13mA51dPte+6SgsHUkg9zVhCzGYpCN5RG6z
71perxndtHUH+ZzaycClkcc4gsdJrY4WwXCwlui0rlYWimdFJDkpgHddUK84S0b3aLmUY6Mhj60b
h9eFlLMeJVxYoo8ZerJjoarOsH8OUO6IoyEs3IGTRXVBwDZg+NHp5aboZ0UybJ5l6wFNatYhcAZf
KiOr/cA3A6D38AEEWQbbOyiu+QmKfvXL6L6/P9imCcCwWSWUOJ0aCz02s7FRiiaySJFCfrfYcfZB
bIhPsM59/mpl6FEF60FzXNb/4xW1L1JkNqaq6evkr5j7JHqTEgX5S64c7dFI7u9qixENFw/IBelZ
eObHsqJ3Rs4FEt29X1TbaOblb5+O+lQF1b44eFH2rQUE8joW2t32xIOmW39ERsDjTJPpFqyD7k6W
Yjk17M5kXe+ET/e0CYQaCjBWiwWeKDHkT2F7cDvx0aqllL5W/vXTz3BeUUvve+ObmYSX245BpHyt
eGeT7VOJwd0CZM4VaRnswLDGe2sJ1MkhrihLNL+n7sPkn3xdosd33OGUBcImEZ9J+AyiIrBccFUf
3OCu2EifMPPweyuk4bF8JO3fxvd8SsXNygkY3LOQBELsIskvlxLlsF4zbn4ijlqYYKeua+sXAf12
Xa9HXiOBT7EAkQIG3eIT1WPiWWFFHvgSQR4Pyv87/zk6g3SfM2jpSsn/nXggxKtjZsU0HhQisQKZ
gmtThe40z82T5+JDlLnWTc4mw1DMCjqodiRZ/i+Lr9xMJs132qRxDzX4U1W8vGVHADTEFyM/weB4
POQ93fcxnNUlcxLuL+pjw8Oy+rGvLMICmZxiujRGL0SzEiXRfRN7af53CBcZSW5cO+5XyicPuYTR
nxrMYovc9L7HUXL4sfsiKHrYfBwfAg+iAqed4rjV9sZ5E+YZmCAXLQhchqTyaUNeni0fPeS7osW3
8CP5BpVQhm6ut0mHZSBNJKcYAfCIyRP3NO/8Y8njemct1rq7EycD1rcc8p6kerotF1cIfkx8El1X
MlE6S4yCYZ2++aVrP4v9yp29pXOPUyPhGPei9VZm/39cVil27l4dcqfc5nxFvHwPeZGL1k8txb1e
HETu1Tm9Ie5E7MTC7TjZBe9abAolfiInf55XYx7BdZBp103PkGbq9WhgU3QkaQRb5LIQ2B+K4RKT
ANyrbcfifHnIksKP33tk1grSijtt+dFcbjGGjtie+AWpvFI8X74tyujCfYD1+VRTOKwbxDpxXy41
X6N68zUYXlvExZmR6zNsvTlUP+Z6Pc5fGqY+oIUXnJkINL9WfMx4faPedjun1mdRuI7/U5tWuwUo
JTjOqxTAGt/POKMRZRio5jdsXJtktyIYq3Xf+KL1GOiQvW4vUAmuDBn/BL28roaGR/DW+mPpUITE
EeNF9GDM/0BhZW3h1zo76Sw+KLcBBxfS0g/4NWqoyyQZ8Vs34Yi3S5J1IbyusfaaZZunOYfoc4d1
6cCOPYU+FpWOnOCr276uSRUcsFogEwUPGNlj8BBU1L/HMRVaafLUes6JMoDFtXpPTWxYwZLAKjSY
rW98EvUx8BA9o7Id+CrzR3ep/GdAIQZWdbTIzRViz9MNRLoa/PPCHOMjjmkkMXah6Pt8KFTpTwBR
iBOq8k1CNYyO1WA8TXStgp5hMy4xP+uCOFew4b+c68drhYqeML4CSmCew+zFZFzZu7abpC22oNm3
dRjpxCERZmJfAEeunfTp0nykHAhVp7nLErLRh0ch/+2+wATHtzm6m3Ieot97V4oYBwe35hx+XcBX
QHA7LIZJoi2FvBjjmK4BgFc1WhVXFlsKQvfovSrFVuB4VBTAc2n2EkVJhJcXiMMY8yjcq/6sNQd3
IsD1qcZIWtA6eq5dEmEIi8toynkA/4FUEahVIE1mb5zr4dJRk1yvrIyZDv3iGapvV+4Z2j2crBon
3z32k84w82e7l6uh2QBrcQF3IxTj6jwWcz6Z6/YF4TSJO1Mr+PcK3Cten3rSDaDEQ0xWHDlnYZ0T
ysKp7MFEmWJgn5xGesaYcVe1Fws8zwFVT6jbkbQNbf3wH7B4B8mHR4fZQmPMpiM0KFns9u0wEeUx
GsjvUcpZcD8f+GbpYkf7tf2JVLagCPXj5AgEhs86XuL5kAAp/aYsq38MejhiXk90kfoGIZabP9Cv
Uqi9i8/84gIgU02KZO1OD1DtCwkQvqKwk8VHo9+Ly8saWl5z5xCJwKCogyYejEQ33EK8PzfiUJ6H
ZrJ5J7FDbVykPopW9+G7Xv03BfJP9yH9uQS9M6qSk5MtB9kqmnsjPQa0QLnG2XVDiG1Kc7nC2cTl
EuJrnWhIZ17R1Nqiv0SGidQVEyybLuLUeQ3ENc9Qx3/kcDcBRj73SOFNvQNmfBjEiUn1F03yCU/u
UsZJKmHGqh6TbMQLJOfsTwINwoe19N0jSd0bhTmJY30ZOOq9UI5gXNeWYoiuAnJGcdtJl+tctz4V
xAOyOVF9FNEVX8xjNeTGJJJhhghAyqSVbCuiBVPbXPx8iD4f0koNIkt+UFTDmLmqFK8sZI1aOuqX
MIEhwzyIlO3L29uRTwjseUvhL7OTV+ZkjVt/7K6A33SOlpaSWE1DxdxF2CnkDczmERvBskQcNGPL
8VEZx5xvnMmvDRkDJu/ywdOSTwLzy198WC1h8EIVfaavOckpNPLOLP+k6Jx/J8maVjuNNXuyIyCB
WwqKt5xi/k6UaOcfo37qv8FvF0je0NoInUQjJfJb9sUnItjn/iD44Xi//Z74QFhdI6T9LvrVps3S
nupaERPNrU9VxqmCK+mft8CMC0bm1ss4bbl07hoqhZGpofk9hoO8ZDL+V8Rkv0dwoUrnF80+spux
QkTVfx1rxSg1vWsmEDu3OagA8N0n4dLYVM4nk0dVdEXIdwpQpZyYYyhWpX2CBp2SIlmUolntLBOe
vxbnKPwUkZMnVs5uvZQZwVSZLd1cZVF3yvT/5SfYBxvdkZU7eszDaysSlK+bG+abfcSYNdibHGBy
pdX8huVwMfTLvd36F1g0YCRxS4+920YbXeQtZuEqj4TI9UBVZIAR+3FW92twshxHd2rF4yppKEUQ
Is/iGL5V/gK3pd/4QadvhkaZOXyxNgrC4VPS6AlfZANpoeGfmuV5+IS4S83MNQXxbNls1U0Dwd+B
TCvene2wiYWPsIghDaLUTOl3G6l8eQ5/KSH4cNGzdUd3eg1jEZJsceBzudSA+DEQdZoViTDkgwM9
7BotxiWT/I+cpKNljI6z6OicXF0OIMlL8Lpp5J7M8eps4H14Nm+zWtnZ+yXOLmb1slms3EX6Y3Q/
FuoZdbQbD4fMOHxC78uTDbvEHg/KNh5Ws2cN19Y2tYILbbYt3XzQpW+5xKVWmFk8KeOf9/FRWOdg
H5xvVyiUJyheueVDaNgtkiP/iX3QZ/UosdNzoJP22zXlYOXhMgz1VVzVo3GUGajlYMr0+KpoQb+s
hPbHIbQQfVffWh+UHtC9D+o5Mnkfft4FhaJPAgpXtKOI7OEMWfVvWWcqATe3ja/UCUIJkfHrii5l
R5wkqQ0haDq3D14uw3xlprriby4TiNNy9eJGzBQQ2Z2Phvn5sMGIuV6+Wm6Kec0l9H/RmfMUp6Xv
JuGPopxntmj3Yd0jmeENY3/iGi3/7lTAaQC3tiW8eEzIM7CoCFsig6IHWP25RcOG3F2r8Yh5WzQZ
f1WTINyVl6q2TMsxLOSdBY0qyBFskFwlDPJs5KwCPMXxV8AmB92IYL35SU6IqZurjKpjWR9wRJkQ
2ZtKbzfjkZTwNbR11v8xG/bqIjdSr7g2tpQY7AkiTDguL2cPb5Xr+FrwVlOUZAnYKqUFNguHle//
k7K5NOKTCyKf8TeK7CumwOwjQdfZTfOSqYQoTA0O1c4su5v1NKcXTF6Tt5tFT2mxorZVYxDImxze
I8TroCMnY80+btZj2X2YS6mIi/3Ycly42kXIyOMdM0JnzBu5oeCVDUtOEV179edzWRwutF60Xo2B
7k/Wc0ro7HOwizbTKTB6vgI4cg4Zx88YZRIacfX6cQ9bNVdMaRov2mlSqqCZ7rbA2M9cM75A53he
AwX/CwiEZ9ICJ/PSZwLYiJ3kHvZ1kXdxLobdrlzkUtVfMyPrLU2djl0tZF45vUvjEMc7zObkln1b
2cLoYd9X7i6XetIel8ctyu/1lG6rL0jX4gV8jhDfr28OsCVazIP+Mg/wgcSNr2UfcxmOI+n873g8
MNuVs89PMqsBeh6nYDaOoPcOKx3ge0sDCWBoJgRKmR0bTIYBqoaSTTEEJo57K7Ej0xPPgpsyZ9Gy
eGpc5ErIe2GFH711cvNUUHX7/Aq/hfcr9W/2fr7U+slubSnuH4Aa5nw8xeW4r+kU6gqZ90xHXAJ1
K5U2Xneg+rgUCqhm4hN4gW2hhPHf+GD2lKR9qsLU9wK0jk6m8KcZXAE/wJhr0s1sJAILQ6u3xQOW
URSvLnQLAD2xWE5oDbXHTjaBrOb729ZcQV4hMxwOPBXKEwOztg35hcDnxusdBqeNtBSbL4OTjgGe
dZaxbxjw6ytbtCLnduHtPRQWCN1ijYyVxSmp7xNx/EElvj01xJ0EBX7rbsqWs5+6c/4KWSviOnzq
cDW+s/2wU5/oHV7TDfUM93yRrq064IyyKoGz3Hyw3DI8fmzU/xVYYJPyGba3TDQ+1bv4ivuw57iq
D0BAqGzBFaRYXZyNX32N+ZJ29YpQGN9ihWXG91WSRAFNgXtQddTLNo7SjxLoAjEM2Ly9iiWlHtse
+x73oi0qo6GSO1zUopgVnDBv7Sbby2mzvgIRYbMhjJiir70ia85w+iTEBwsoBjsxH9lVusxKYUft
N5B3VCxmcZ9F7PLa/inGaTV4pV6pnpatVDHEm8oBwltTPVQPsZAxDUJggZPGeDCGx6+B3vru2pYR
VG081rKHfC4ny13/iwVeh/LX3OV5GbfQzSeMKlHXxBPC/+8wdKuUjpXF9xw3vZTk6UEKRzFaVv6s
CPQt4sjyTVOYSt0e4xxsEsUifHyPYHB1lhmpLCt9XZhymobFQnCYLcOnePFSu4BF6PymEU3/1Lym
Hyg3BCpv1XdYehbrNcLPhzCNrsR47Pniau3zWg8qHSXHpmilKHdbJjoCZV1TkG4uZ2HTfAi30SLi
xxRla5CLdxUMwdW6yrYjaKtxrrb/wA0xa/1ikZb0AYkrFYm9PaYUS/pRydWRBZ8n/Vn1i4J5gVCL
BtOYR1dbPFcTYrTYz6MzTDMsNzboiCd2lHr8u4yPpadk++GHT3Deu25sVX/YCRfQDC6yETZ4VGWa
XHKtnG4R4qk1SG3zS0DSp3Iq4FlUSFqsRzi5cAT3LDol97b4a4V8JrIVVKdZHgmSpLUb0l/x8u9H
ihP2lpTO+ns8JvXdUEBIvOErsrtUbtFQ7x6wa09sGb2fIoUpBbBHqap9+1nKnBkQJ9jNbTZrjPL/
JlH26NTjDo35B62Z9T1fvcjQ4m4eGuuD07+MzzLMoe4IjqlyV+9+POH6bZ4Z+GfcbIb/9/G1LLCs
Acrtrj1u+2+Hk0mQ3hdrPbkIGnFf+acsq1jniOKrHbFPoJoIi4x6Z3NDTmDhTielzsoDwNkJplFW
PVs9J9LXoN3+xpW++Cn8moacdWRsWUZ5tqoz5tK7N3egV2r53VeEbZbeXF0Ok0r/V2vl8EyyOER6
+PEPlqLh+/MDnWntcMdNjbykVNcOuFWGWCfe6XYYDYRM/ENSgEjyQdakQkz73jN737rcTPpOSn5S
+PUH789sldclVlv6JrNux77wGp2nVmBhAKrdhT8J4I20F6cfBf3xLG5C+BEbesdH5xfwwvT7vlLu
IuVk6P9eP7b8u7Hy4QBXaHwsL3IR6HY7ohpQ7CB+JvxEdsLPhVe+e7PMD1A4LPQlE1nndgqe6nJX
G4kZeFdQa+heLPWHSNMnGkrvSTheLRsZdtUr2Dz6yJhHXsiTzyc1jhvuJ8t7EBjMsCoKOMfBIsYo
tr+4a+FB1FWOxU+b+HUq0ctiY83xzTp47jEpCv6mgbxgPaluO8Rt/bFTGmk0uU0G4VFspLl5FZQq
4o4H5L4YLsnhJrl0lqqvi1ZxPh0lgLxnu0BY4lhh7SWfYNyZeBCjSdZ07DohMr8x1zdlNiAJ8+Ek
vGMFoiiAZAi4RBAe7J9R/HLfrOGtWWtB+PgKjo73CTVmIiGkRR8ADjG07qOo7T/QrGpBNnWYt/N8
n6RPkZ8SuL9jr3Ztv2yDjmpIBHElDUuJXoiMCHwy2tKg4+dPl1ZAipGBspWzd2Nn3A4Fm2BwlxlW
U4G0esFVm3Zi9Ap1GXgdX3pI4tWWNbdx+GJzTtE03KSQlGPdp1XA68uW4RYr0CKKEU+G+CpIZ3NB
sskwqy+U6v65BGDxsa58+1vsR2Zmbdtf+FUUAJS/+5WmJGYDY0hhIP8b8Bvi6ZgGzCIhsXX9kh1z
gvv5oYMfm9vR9Rm0flgkeSGmpNz7oVdFdS0CZ7z6tvrhiOQPyO+iMtHyC4qrmRVVTplqgX4P6/+b
ayGhtOXIHzl3YiXTWbtgTp6WzmHCCXrmKuA2L4C1eVBxwDM1OBa6cEvGf5S/pKyOFmRECvdkCW+k
pzPmDKHEMiojo60ORMivVy3oImZxX7ac6Fxr6c83A+NT9V7Bs4G9Oa8qBLQAhZlLoLlD72OoJO3K
UfrEs/mMFI+3uu6R9fUxAmcsKu6RhWzfW0wfW8p8MJLe6EdyvygMs6aogiULMF6VXfxTEhiRV1Rf
ySOT80reZ8TjPw3Q7s1BajMY9N8dN5a4ja+Njvn/CsHRREtF23pZoIqQu4hV/LcpeKWH+WSzGO3W
rPND0lP2Q+0VXOoNReS9INKfAwHYH1PBnyOy6H3CEOW89CmZ6XGD5t335C4Np+ov0XGEwhyEZdPU
eMBoO6szGqszMsmoLKxP4TAz4e2ngo6WtpuXQtKv3xYiVStLRlOh7o7w5oGWZiQcg4R/vvSM1UzX
kN2V2cbBamzkPrzyel0Eh3YAcESQCYSjof3AAK/RIlrN5FXjApM4gCchUjbiePoDZ0uqueAkEoNQ
KjCXmBEXAOCR6huQ/D39OOr1s54ypigbb8jbNvw5zZzEZoJAMWkXHO63FlHC33PwrDttnfsaCCtj
lDpevrhdOyFyNBPgZMVE9jQqjUqzTJwzcN6RmCLHhtiamttkDxhxzgZSSq04OfahHsDKvuuPr9AS
SifpmOzl7x1qc9VT4PEjJPosX7ur9MlNM7V6Lt+Df2ZxgyqlnvviXDyp0ypHptR4RoTs5Flbs1yz
SUem6GbCOOZ7k/aJbFzIZYFLwGC15CjoaZFOo7zcSlSoQrhlTUpp0xopF4G5XwFHs8CY3foNdAfE
QlWlXzZa+Lj/LHV3yTdmfrwAF2AJt/gGJiylU3wk9YoEkf/RJGWUmI6wiQzFIknM/MBbsQuBkQaY
Mx2KL/uq+T1E/jd+FKMuCeCpaQ0BR/4k4ouSm3pCnIVZrK5fcRRU6bNX+nCEww7jDljr2EssaM4u
02fes3ADMV3xy+XBFeKHpA1mf6KC/f2w/5I1rXOqkNQVFOnRn7pw9E48ElitGwnwu/6xNkxLrfbt
hzIrkmJl1zKeBsiGCoctCK/CUzQeLzN+tGkr+pyL0FYUnV6X8bWvUTbJ9OLcN2bqYsKhNTXlvIdK
OEdfHmWsw0lM7mjKrnrGHPcw93rQL1pwAdkKSfboqs/FsdAAxe0hXjHDfgeTStLQ32c9Iu2ZeTX4
nfG1sJmuvrHa+v9OyUms7NHAL5A7vN+F+T10XCgQ1fKaFN+hsWS1RsRfVe34UZJR5Xt7qM4Xxyv6
YhVqapAh/3dzMpqoV7JuqFq+T1sPjOuLSXGvJCH5AX7hL7mBIYmPvSQosG62o4P/yf5m8ui5kzH1
GFTZx1xIiGqzsqAY5wqzbgD/fevVdHWxzVSZlYq5CYq/5oD2FyF+PbSxokf3+Q5RldUsiTx7F+9D
bZ1R6DMq+mT+tJx1qxZHN1S00rEaC5ascV3tUeayinIOqPd6rZO7BzTLoUtukXUsPlD05AU2Mw6k
uihanQDeyxW9NnszHrSqrY7saj70LrNdk1NrGqNL4pl0Ag/IEIytW1b2wyOrrNSkZcWi0l3ZIKyv
jRR8KAQJW0araxlpxBl2Bk0SMIAmoEfdKSWqxjOGy61nHaXtDbRgSqV2v2dDZZUoJR70aAB4PB7b
lc5WupyTUviBCnNGRaNHx1Xund9kxLW2hTR8bFRURSV8ygIDCPzmz1qenVBfjRxiCMV8XDiCSl0W
M8+8RPcM1bGomiggu56ilF0ZLfSrfuziyEmksvHYg3XpgeAzWrkg3mMUUN/fOGijEhsd9glO600s
7V1TCDv6/Bgmsodms9ndXaJlq7HdbTQA22wUSEHsSrYtnQ/TX1uMFBK5Nt4qNt8g5hAmakiJT+1s
DXJuZ5pZLqSa3STa8CqlSmqqpoHgBnOM7/G8YGe5tUGXqVj/5W/KD4uhSLDYfO1rCKonZsMyH/SQ
/A7+9j/6ke31CecvFCfDxrTQtBUpnmEFgZvi1mzoT3sIAorIGEE5WcuCN4KOjUdGLLar98CFDMkJ
ZM30W3UwOQFVEtirmymx2AAj5DrI5hn+gwabRFNygi+9cJcz3GgOH6d/p22qvftCDZJ0OPeeJ5K5
ZPHvMSNEGlYwcYL6wP3qq5035+sImonIUdrIr7uooe9DxmhCnM6aPUNfcYqy3IP0BEqtNK38MCuz
0W+ng1Qp8lwFJCRoUW7IwKBlBlmAHhddSnqW3pKtfBWDTOPaxM1sacyjtjEZLNEVjtbMTLjnvdZt
aRIHvAr2h/eB/q9nbkvRApnu1vY9UNLJVg0j7m2OYFC2gwUYKj2frlRiiDY4y7rQrzR8a61vp5cM
S8rEyY+BZVOqU0qb5eE8FDr2FPMApQwZgDxN5TmPcch00mVZ1Keax0LwEScIwih05KPk0PSbhj5s
426U3ajVX5Yudj7wQYE7zAfSvdO8gyBEjbBx0P+WerBSNkpgMCUZwVc5Xg2q1poyAM1ioM/Iiojl
e705T0U6OcggpzrvVgTYz04b0Qa0t2BXU0vWjm/tH8ynP19kseif21cTcb1IKzKPeqbkSvDNNjHI
/Zm+PjAi8eYOcxErpflNehRV0T+ESLlIoul7fHPd9PlLKJJza4YKV5n/YNCSRH9zUq3Gt0rN8cRs
WHycB06J1AofIF/6pKm2i3Ouij1kgethtCgoZS3kPPyRqVIGiVHzVZe4AkpR6TcycXCzvqYrTo0M
hSvYqRp9LYkKRt51KxwG3DadaX3z+IH6in0kyphNM00zZRry6PWSKM+mIYPerQTDc+SOF/qD1EHc
TAJnWEcsYA/fHIzILvFPGnQKGoWNW64n8/XPLQTvEG/q8YOBbxY3se1YFJOqyoEz3v7nZ/5/uhgP
KaUiC4tWzp+D+IyKJ1Fe4moXQVy4/QPp7cNOfPbcMnv3SFgKoR4/zo3FVD4KVxZesAYJmtV8swbh
Cb2Df0zMIhmPo5UuCsBivPBag0I4O38FsGnyuhS2zJb3jpFsoZpperZ7FnFNdrTCO62qUKGZzXdo
FAZAnon4QdtV1NitFslH385RVMp1vetXkwhRPppQxfNT5ppdSM/TWj+NCY4Jcyum+krIFInsg1ov
JDgmx6fdsYLKarTkAWbuVpIfYsCh5xs6tWitSryqi9gk6xQUiPqrQCzhUpDGeUP0pGlAtPoEIEnL
mPWJ40qcnQe/WGFcasovNQOC/Ug4rxa8JJ8pj8FCOic51yERl8wRao+SvysITwrdaWV/ejuMiCFK
WDwDA3A5n5+tMBsYKCvujn28mDJuX1WhaKJzr/53gqOB+OkTqnWMD5T3YOCDHQM14cgQdgBpNPUf
23L2ph1gNn3rty8ynnsQnC8mkjAzIBnQy8z0WlgYud9Tzkg2lTpPGwun1AQ7Zb+YuLDiAVHN565B
BCb9Me2EOzZeqZzpKB6Gs6yhvyFECa0WxqYEMdMgiTkkTR2Una42qCJP736+S9WmtdmzESTeo5+e
XlHldbXZtRBDW14Tp/3aBQhreZH5vFaG2oo6CJeN6SUIWfp83IFsYUji23WdHlNtBQSFBxe92cfY
/OUxQWylj3LKPgVohTE+Alh9+EaZIjBDNZzW82X03HufUDITmZg/RftT4RlirWtsfZxN+pMj8Ru0
0BSrwCql+gMettHl4ptzMWp0ZTKxuJ3lJLjhBRQjqC9QOCwTrwZ894Qu1bq3+Cgqviay9G6HqeI3
/c2vOJ7gFYx8M5rK1Ssm05Wrn4Nr2+ih0X9nrUI+HHWRpsuPHpZeC4YNeaJ2ip1zS9v/s6zcnWsw
VRQZgkvGPF8g9P/BAzqX35DVXTrnifPhi1WJBjHM+3tTJ0guRHBVZOTnYYMKIlM379lbMCfdwWLZ
AFoY9zOGSTQrC7oQ6JvY4ayB/RnVteyReDNWNC6Ib5LqJbauV8oryaZtJmBwglx6eGwButzIMPBL
pjT+lqeENAcHWTj2LyFzpKfsL6tlzzmqE1O8D+zjRmsfLNjX0msPdMf1IHVpiaaS1bwxq4MVzQnV
IHamq+9pxwQT+wQLDvMYN2Ee8Ec39z1Ly6iF6ivCMxrhVbk2ryQUZlsmqQFvrcRBW3BexBvOkY+S
dlaoXpDKCArcuucyUoKPwJQ+3X8ypk1ktdOdV7nr4m0DfIYHHCWU+nVnhrkOjhGIq2XpHkLjbIxB
LId8/bKeD7VOezXoC5Sr9RBwXe+V4oFjwSzVLjk4eERJ+Qrc1rPgRKNHaxUkHkcdQrOsVpIPUPxi
/RCWofoBhSxHW/W2zWV2Axeb3M9/rMNZzQ5CJ5H7A6nVHS4dnnhLYfuD5vQjW0guey3cNbQn8r30
CccSCU3tdqMu83SqOkkMSWHuuGxxnW3UOBj+WzVJOKuBVSrkRija66i0exlz2QsU6brhVpWSmXro
7kjNKalXqehmWAGO8rOD+CZaqKA+MQeO434OU8DvIaB1a3jIeo6IW2gclnoouVx9vEj3O39QXapv
Q8gcNAxoWhrod7rnW3s59mMgaekLXIr2i2tmKpapQRsj/BlWB3KZ4z7zkSBAtBLkAPYAfNXR8eap
/0vSlYfCLJuyznwxICMgCtXSMKsvOdMrsPZ/H2njFgvkQx2A7G1XGptMd7owDw1MxG65eOW8kEuv
UtbAB2nEYydUOkgNfI05H3k6iX3wEyULpFmhrlwVj63HZaOGGttgmWiW8K2UbrlIKYn+1Y9LiyC+
7wRCkHus1UWN7QXBuE7R6oSvCQ/NlhoAXMDZcvpG/lyMRGE4pmT9zrXaneT04kJ7kq6yfkti3ehx
yOkFViA0WDuegsnxXuSgeTm94QXzSJlrOyY+yNklaqi0upeq3JO8vQ2reOsHi6Muhwh0iNqOm55s
BPmopB6Is9k0hfHZzPeAgzsDr2gRmesfuUETLipvxztLTID7ObCFbIBvcj0Mj/DQLmELO4GyUgSm
CIO0QLey/2sgYakHebExIDGr26PpfkNTIkSXfvt7yg6lzbeDsfiQL6mdpMQoTUQqYG+7ooXcUF35
CxeDf3DxR/ycDX591Gfg8qL3AnrYDIALMj9rO1MYVAE+Mp9K1fXmgJcL2yfgULjEaELRWCDTzMTQ
vdWVZgPcryfq+iWTZPcwegK05lchSHU5ABQS/f4MTWh0iPgEBtEXTePS3kpQ9iE1/FOZcLjS6O0F
C63HFT9uWT0BtKKW5sM/JJIoLcr6ZyuJwRCBb21mInnARucqJVWMzGwbj9qL4OD4Eks1aSWJ98dy
jH2kqFt8Eyntm8UVvkxCdw7N+lw0/WGfpMHxJrBdU5oAGvDBQMg7gKqRQeKIVGQuV6FPNLq+7FTi
bj10zZrAA1eSUJPe7P6hWB/twXoEWCk7aQNSwM9WoQFgkOyBaTnboDFPPerZRlCzcgNyzD1Y9wkD
UpgGsyzCTQWZbQ9DzyTg+Dkt79cC9eDhQ1yxy1ugVZDzrhf9G3tLJP5aeI5EL6VZv7JC0HwV4HXQ
GEYh5OUPFxJyWxYs2khnPcUXwGSSqoocgsrpGAH3tbLoiQK7tBjNCf8S+wLY2dZ08fbkp1jp5Own
hUhvqcNe+4p+dtZl7Ugu0Pr67fHaY5FitTKCe+/fTaQkLjj0g0qKJ19pw4Y8eQc8oBbZQ+zA6Sak
F0Rd/laaqcp6EOXwVyFjFxnCruuvVtj0IMjgrDS0qLq5sqi27y53ibeJKrH0eU5ykQ3vtJj69ffV
VgvqZ/RqGrVwHarKzaAjAMbFm/12dU+VO7XFRuJdXfznT11XDXeowlS5MKUDEJ5Cyiw+U99fmwy5
DTph4Syk5SDu86oMFVAH8m0QBNSJDHMYsnCUySnMI7mzMb5QqUlVNPzFFyOBYQuomue+V5FRLiIl
cKZVRQqWdJZ/cDThcd+fwnYTGSQsAP9knfL//z1lada1KBMPyj3PUr8XneOVnjLTeRK58aht8H/0
24iHqD4uIINba2UsH42yLLAvxA5pdQQBrC6X1hS91+l60Mhq8j7B61jJC4kJRmFZ+ZgJzM1wnSbS
NWDGOK6S+96Lk8NHwieb2ZLCyeU80gg6sLTvKfAj2uXDwouDE8Zq1mzo6Um5bOe/jDhmmeeDpk0U
SkknjYDxkayOvLlBUvX2z9tAio0KBjMIrbN1+rwjLk3NLsOfdhqMNS/89ff9qUtjcRBisIa06lE7
+DOMA1E6BKNcG6GG7L51ck+8FMKGTjBFDuqavl/h4FCVrovu7e8G+cvVYuK/6U/1rnKbYI3+xYS9
ud1OFvTN3VsPOxIxkZKY4mNgBknXqKa+mqmjuXX+Y4NoeFEyoeCltP5gFLWE/d3RJpvzMuYipzsh
zYL4mpCctVKPIO6c3tjZrzXXhs65o4xfaapUg2ihkBSOEycIitZ8HQFVB1+uoS428Lp7X73dtknk
NW4Ky3NqQBPANOZKqoaPID59z25nmPjY/qUGan71BoqfaAV6TZ4YOfAPfQ8kh950iTyVcjV0ZLsJ
OW/F2VEQQioseOp0ovtWCYj+XEDO3SjBjXEP7O1957nsg2bWX+Ff8uwoCe41jfRAUPDPi/XyZXIL
jy+gPNM4wb5Y4CyMljgAHaY/arLNGhTSmPcM7TmEAYFGSvy/wUrH7RHiiyp9hifvdAAHxc2M9kxt
H8F/sZ6UF5vs4cNg6mYwYPDYnZYkmI58bbXzuLeYIrmlvfjV5Esmud2q7SlA/LKv7+15Mqd//ydb
VkIbw3VMGSQhQ+NblLyM3b/KkQPNbGDyqdOEX16J1fxT3zNQNmeYkURj/2x8y3MTJB3gLF51BCy/
BWhgxaMckE7hIVk+m8DdacL9Bwr9mIMaNx0TwBw9TPyLQJIMH/Q4YPLYGf2RP0N7k5/6FH7+mqk0
bcbAzSHaFALpOwem/p+i+6gXZyfsLm83daoR3XEnlhtJqkQsECYMLFnZt1S2Qh0VRLFeDtPFFQ/d
gMVG9LQMfq55WnJcdOsfkmyHQkG7zGE+3XBgQa5RGtBQ6a1q3rWE3mJ9Jc/N3NSIyuVVBXtCaMwu
pHV9wcPtNfyzV3uXc4pdTUZk7Ih1Xoh5ydM8FhehkaZlUY8xiV8Jbcz/HTSS/8orr8UUATUheqfD
VUWSFYT+Aet9rSeC4BT52IzOFAE07UP6JD+X/EWviiilpJgJfLYy+RnO1Z9BVXOonTiyVdUQO/uq
1FO2g1IfmqxvZkHCrsDcQvgXC8KraUxImceRMiladOOaaiX0xqOr+ywQHPkVyHEZviyDpWhh7mOx
2tAa3z9+UKSEJfLKRifxdEeAVxWaHOism9tgyhWeUIburyALm7i5lClUl8JmKYSv+k5XVaabrla7
TaGYInoU0C9ec5QWVt7j5Phe8OcOmr/GQekJOeF0qat74lB2gG4inT3mzQxyzTU8gWlSGm4mlEtV
1XQjggJcKT0VNRkcrJSZ2IRmarxDrsdwhOjcZyv4XGTgEKx/tebC7ahejOukepoCdaqMFRnmWVut
bTK+AHNo1HSTYnfEv++le33YranvUMDv/ifEUI2CrxVAxT9JbozopCEvv9ncOExmBB8JgJBzHbfo
7Dtf78utPyOXtV21rmoYSXTYZ8Ui/vCHsmdxFFJo4Zk602RpFkONnSvYIplMmGnj2W8fSpYpm0xs
fIekwMOR0ti659SJMla4c0WZs7Tho6Ag5Tgq6w3xlZ433zs/2MyZl0GvFttLdySBK8X+oFgOQa4t
K9rdGQdqE8sptSm+pPYsgwBTs+GhGxx1en3JrQSGLm+l5gujCXHHneREInXYf+cpVrZ7uLxjs5JF
HVkzjzBRos2TnZEXZFS3xHX4MqF0XFt9+Jj57zHdQ04V29vj8BbsLyHmWkrNJUIcZp1DM75ijFaf
Ds7flfjQzvtkdIIE27fdC1fso3ym/vbE1/l67zgvVWhiTQZvTPbVcptgtDS5EiMiwTkKHJSJSNa9
s9TRK8Th/lPm/bVLJBTmKV4+r8YF1CDzD2sPIRO+kVDh85VX1mc6XajGAZwHWqs98bIffB9FqjmI
/0Ps7MoeKgwmbsUXRfpkJLn1VfqIt+Qy8wpSRLFYyBv1CBLSkkTGbmNy4UxAdI58qKxBwSNDTFvj
CkximfU+p8rYxNUtJDHhYISANsUzZu7xpjnGL5nR0K89Q8Ja/7de8epbMrBKcxWCgX/ZL/EH+3ZL
TpOczO5obu9/YJ0lACYsJHJBOC3iieNvw1GJdm9+vuUOnkZ1HcoUKOoaENR8GV+OuJ0T6g6NKvne
wbR1JiqrGvbh1mfYdJfZ+CRmNusluaTOwVN5eA79cF4/yOkN//eCl45d5ebH6wM/nlNxUqYr+uXz
3G7+fS1wuN/uzjTc5xtlFuR5EQrge8z7nkxUPZWXmXvuSbujn2q79NA5dW6ndi0JlCCf2WKkbZTI
xwTqg9GFQYyasGlfYv1WaHJSEf801HVzpgWRmadVlznrjpgXP+9/NN0ZV+0XuGK9+dvNOeT7RJ2u
KCpLwSmj7Eg3+CNa/trrRL8qD6eK2N5sWn0iAQHS5zCtB7RY/9E7wLRR1ACQ5NLXtIdvlbbbWNQb
B+U/jUKf/9H84vEsIP2qkzXiKgbBrrdUf6Duy+D54sgfEn/W1tcXFtKtCOQdy5RVhq+lsHwYNNoa
3LzLCKfgAqLBwGOCll1jHGgeGsX2ww1RJ4mrvbXzzISyNxWtk6+z0bq8Rmpv2OpGz+wU6CQL5ICO
qX0iv2xE9UyN69grisUYbSR5ULkHKu0qs7uBw/1vFEQwf2NZI8cwMeEae9S0/GzVXCGeZeDvyljB
pN7R/eb3D0JgH9KrozS8l5jjDFZ6pCpvof8vid9isSXUhZkCshyCvyllSmZsUrQRh1fqoUtMI+II
ez76bvz3hJIh8jieEhJ+Cv+Z/BSRoT5OGL3uQuxFmsRDEwdI0hHPBQyaLziLPEBKGOJNRdmb+T08
dZo53O9zL9NUBiId+skTryWh3oQRk04+D3xmDxh7ac3vKyBRfvAuwJOoeKIg5nJf1Ws6n+9wRNIS
zdInU2eSjVSyVccAse4shPv6/1Mi8J5heTdj3zlg4J9L7lJDHNmCGb//VXRbjjcjRb2Hb61v5LcW
gMSKorrBPZ4qUHD62oR1QGVQgzA1g2z413ESxCIEdIHliRWbgkU9wzz5k9LI5sApV3Pxx5n513vO
eE9QEbfBMiliY7AYa9auMocuHKKS9fSl1hC+e5NkBMYMYWonABzkswwFfFdOxmubFVwCmN0ItgRJ
xORv+0FS07VMYtxuY2o6efQoZrFgHCQbZKJmAlauSgnhhRTiSectGcu7OvR/bAaqdkK7HLdQatu7
puBLM81eHJJGVFAAc57Sb9jqYLs23Rw5ZNnWxHsugjQWzuABVNXqOjF2nY2E9vbcgICZsCEl9pDI
MDz7L3lkzYcg0uxXO/SNJ3Yl/G8cmAIf3xi8ZAWVoOpwrNopDfjtYv2SdwfPezWaR9I/XI7s4G+9
h5QumQFzU5yyNQwcofPOWQXrHiXoddmvfUicWyZEOlhm6dASzyHabXRgEm7y2Rd8N+tQFRi6o+ep
Ygn+XPj+nDnEFCStlvsDpsq0iz/EzFzcTuu3HFIz9Eny39KJ+NxUwFScdRjQdTdC4wOZEl7Iw8zX
4NymgKYgra6EOZx9FIQWwkvkNa7NV2GuTVFwbVl8qXLgzlYCjKHR4A7hXA2UZ0VieYVp6ceK3zc/
FAYKLYUryooiIiqAC3CplOyBVXbqJ2kzaHm/5Nb9jJowgQ+RWl4B4LV2VHIaeFSSz4/kqx0zycso
eXoks+lTpcGhaWW4ABIlZdSyXOk9h8qutuWBKjQlO/Sdba+NEjfDDqVqEV7gnWqc82E2n5tarovH
o/quOTbwefjuPRA83WPtju6vrHUcyL/OXgR2wr3MWjEJ1ispRQ6rTnbmuvxtuLIZIBFJYd2RXh0g
6edVH6vfE1v8WbGVyHnQsCEtzk9znxGkoYLTqHFkE3IkgX+Psm8y/Ps2XDOzx1ZeiPyv5jl6eBR1
iCUFGkr84Xzacc2IbI1DiMaflbbccV8OcsEDncUTTGswMten6GkaUsmOFkOTtE95CjXj2HhO3vZj
fh5IH/qIwB+iOTCywmW8AszuJJinelmwE3vQtVJLyYZ+xLJ59I3mZF8o6BzYahhtOYgtidVhMrgq
o7IozPNgHIzSkv+LTL1vUEriPXSeQanf9HCjuHqExsCjpR7e6eHZ3iAuRW8ylQtBfdVbb/lA8c6x
CaBh44N1IQdD0mv9GI0fkBxcRbjdNa/WNq6HAjEGW1KSb0hV+BrEUu6g1VHjGCSVTD11t3qv3Aay
ESoT0Rso8pqtes349SuWYJrjth88Uuv7A2SzAymgSxEyKUWeoEeRVqfLrqOhyHfqg1oJJ5iX72Iy
mq2MnKuBYv7T19w9hwxN2PHx6ZU2CscpJf0AbyJDlOsOL+S5uaVkzzGdEESHDBxoffeqJ2X/W5A6
sHbxxmopoarozyafj0iVZGTrmb/AmZAkis4ZPl+7VtleQAhYhi7/DfFW7L2sXo7GhDn+lJ4xDUSz
njON546EOVBDfivnDOkUVOsF5H4xU1i2BljUUiXG/gllLc5jIiviq3U+Uvyx3jD99w6gPlzhrKIh
CFDkk6tJnV8jE5oiNDRMHc/kVZdPgBcdHQX+XgN9SDL4SE/GV+r3vNN18ZFbPDXGh3Ry4QMv0Hsg
XeOVkUI1BVxV5LPYZ2++fFhXYXiILd6O65tnCXmrVlR1fgh73eHG49JgGOGzy6IZsZfQqKSMg4bX
1Nvm/3v6DUdR6rtivLrQiF/tSe138yjiCiI8qZ+0EZYsPTCGafkUXZWSPEyx+Ir2pVpQ1+6gI1lb
PShX2csA8pJ9qz+S97tk/phXtTlEMGclUNEdn4zZrxoJiEQvFnU+qEnNbNs3PBu8woR+4V/pFZhX
KxaUP2RA0siQ2kI+c/Ycx8WxdBTmN0lTgzoNM3WglLnfirQsph0kKdzBPQqQi0HOacs9igS9WKv8
GtLeCc06AxFtKQIPwDFd/6Q9aYLXVDZhl8EdvAk0km2I6WRpoOL4qNv99C+Z3PaLyv5WrtrSG4sg
W1ZUwYZeGRKh/jQDQ3Wl4xDHtuL1us75ydYJzECF+gapCS2pVxOIOdjzi9VeBzFmnf5IF7GYXt91
2tMLoP4LE+aVL6ShA0zb6ub6tHkLJQcm/0LVS67fSTFwcYoJJlUwiVXD3XvoWuLTmPXrtuYketSa
39JeoBvMVPk5ffkH76rtXGgVWp7rq59MRcb1uIUMWT+hm2rCyvRctUOr6E1Z9QQhvmBLZkoCBKip
n5ZWotqKAQXoBTbD8mnXsAi8IVyw1+mIEOB89aCdNM1CYycypHnBV8pYgBLtNByNRyx0OOLRqInV
tcv+hPIyPMMIIejYkM/XHuNQYiriHimrGWzIJxiyR3TYvel1ZxIYluCqmkYYi3QHQVZ2FtfVvQOm
y2Yal5oebJWcieZ+Tpfl/Fed1JCzC+eHQB2v1FkrgpLwZvn+HBuKgEwf3UeZwwMd7CndxebM6IRQ
n02TnLxTeScoEycLZPNGLQPdv8vHzAOWMzrmsemFUAHARl5TwLqxwvjWAi+yjraUhUKPB6tz5DtX
cwbZhiIq6iZMUF+4w+Ef4UoBT8FVTGqCZBswfva7Qmq+H/79wlBcUnM7sIw+PSyWJL+B1H7SoJPm
bSsq1RMIgx9Zfd5UdBsHl8GWuAeMnvPczGFSBC2i2vR4jMsuLHGuZkvpOvu3kcjiM9WA1AH3oEtv
8IIJQMW2EOsSyS0KYhapRHSZwGeVVD7Or740EofWaSdX99djodPE5tzzSD2VV7JoPBm/V8KVeZWx
DIfQq0MH3VMoVZvDTBZh5fUBrZCM6xb3LZWqLOF1Q4njil1wzmJVGnKFelkrGCrq/0Ef3diN/UMJ
xX1toYZK0ZNju+rbmDSpQ4mPKjzUdcudHIVCUmfLXoVK1Y1fxqK+m2KpGlUC0ZcKqStVnNECEldF
wwXz5JvHxbhPuPxa4tNg16SiFjmDMg6dcHLB0VGt7EFY2Jhy2j5vnwwarFw+XO3WrzsZknHZnK+l
6/WhwKIvYifR+08mSZVrfG3LATxVVVrnLslCo22aJ2A7wDM4QsO60MEIax2CVynYvcd2dWafILkz
1xRp+1mwKdF1llIlGwXOeKETahp/XTFeOrnHSada3cweBZzOAsu3FNwzUMSffZcIfyVyGpFPVL3n
B3t6CDWT58WzYr41bZ12TX4eOxIrMuQ+gZPYbCx+nXCRwcnOR0lUgVGtFER1NnN4dCIWGv20XO3R
eTuMnil8WlyidJi7PwE/5hUDYjLBN5L+SwTmegoIhB/cOWgAYyKoHjHIhIP3UV5xeGambwNoGsvA
n1MVvtcA1TroIYTpHzusIe0RvHhO8/YE4DBiKgYqRfOJzv4aw/08MYK7Q/G3AOKg3uZ0hNEo/swl
hn9TTjurJo3t3JhcAYMND5w9OkKMNajPjr/tH6Ss8O+eeecsd8IwIzalxnetcsR6UtN4zyjYEPL3
PanX4mQ58485fymwQQxX04enT5CIKZNHVtfcnFAr9MDX01IYOUg6gZSM3vrHNZncN1uhn5lMkb6R
ZvQAIjt4GHfWqM0LcMi6BRsXmedLV6eegzWbCxYwIFpQr5+O1DhBrpCHTCQVGYYKV/cUF4yaD1MJ
3pfBk0n/dwEVgi6XRVaeaiyXDxhvWlRlD2EBA3E/mUxjuw4Sy+Htn6+AH7tABHefwE6Xf5mQiim8
lkqigxZylp1IVttyQKFomU6nLWWRzmeA0x1gPoyhf2B0DyEHP6rfFWOaxXOZNtJrUVFWCOaFkP42
H8cdVbDaA+32r1OaIDsZE8RCg97Au1LuOwcUeY9My6BeiaWwFULeilLmlCjQCZibnD+I0WbnBnJO
Hld0ypxdemycnvZ8fXafUUbCYLqXS+GLDTpsGSEFLvu1yS/vv0IabfCoyBNMzChwZ1YK8kgEP2jS
Jdh8eaLnHOzY5lQpGOdEPooTmNfBP5CrlV7wVG6v0kP0yQeWDEQyvKYsaY2FoGDPhjFxH1Oe2rDl
ibzOsS66G1xnVTKXeiybDkD3QowaZ6tXODJ3hQ/ja5C09Dt1lsZFflg29UIl7jrLmzVIZCfn78EG
28aEP9lD0zsBewNIDYuJX+fWYcSMJEAGy8kjkXrIsnrIGrf9JmAiohNqdoTg+ZLtCd1ocKfl1RzV
0O5LuID92XTxA34RWGNwyGHGCBY59LLR70V8gdCyyNecrBxFspp//kXozWqWmdKlxrafxkVVF/zv
fG9P9+VBNDmKu4wpk6J9mnnZHBhm/xAlV9v7FjrCwk3YPsQdLuvCDB0+Ma105E6LX0nUveqrA4yc
oVc0ABucdgnSBaCIviIXF5rF8OONYPpt9floKlAivKIsa8tgGdlj8Y887t9faXiPwdjU/nzqeK1y
KUhEEXWPegIdGp274qKi1vrf3RthaaSugvYHa6ZKjL/wYuQzHywKrONQkX4PxZN9TTy5hAnouEHv
9wdIEUi/cqCJpk2In5eyFg9NYhE/S32ht3e5iJDv4GX+pasEeeAzkNjuFnHPc2c6sjP05qGxwERV
FTBbJ4sa/RnzTrBlqHZakHEWjx/jvHSsErlMrv3/JdzRfF2osbd4GZmqegkoZRMtZD414fWq6LZz
8PQMsAgFNomYDnsW8gNANQJbvAJNmYDo2tePlv7gwJF2o7OPM/9ngmDZ0x6/eJT0QwYLjsmUbvEw
ZW9YfeOb+f8EJQPrSy3kLlRPG0gkR1yuMmoDVfIrmk94q+oTK87nQmF1coGdzfICVjQuhMH6DEjG
hgGJvEpcjaZDMTyhm9RVUp9unIKArBDrJoTvciX9B/QqDQ3lxQu8zM/gc1omsgsx2KoI60rI/Xod
IRnXgrbgum3HVKo+YKzRpplXKpMFILI6cLyV2Fn8YlGDaE6vUOBY5gBRagq4+InRrVf//LwqUzlq
Gi0AQU/z7ZEF/BPN2KEubxiw/fkOF1NkKsLeAHIf5qO0ZBqb8jNVh5JeFXAglzRb95JPlvetF2yS
tdT8aQ0F1pv0g66Nt+BWNRv/T692PJ/lXduKgHz41pzN1Ba/9iVUGfvoopKUsEZ4YP61pwHNPOmI
f4KQtdezapUocZEfy2WY94fERfJikBDRspznl2zOBnkBp95cXhgtOq6E/fF7zJtVoCJWAhHMFwk7
LUpDpTgALCZRQqOIC8RQ3P0HxnnhIrO3t/VccWLfEJ/LDw4I5x8OpfGh+QRb3FPScrUVejMy0GgH
gHst+7V4nHV3vfIffwFWqJxLuWqwr8XFgs1OkbKDlEZkLT+fIFZIDqwzzqoJFbwFfTphIBfcyNXR
bqWKWIEJkwgSUymd6H+ptDKX9QrsqVa0g5VfcuPDBYZUyWlmH5qe7/gES0POlfawqnAw4EviMvg6
ghpOhVhvLTCw3ybRE6IUwaTf9CTOwH1cJSf2o46CHG16rp0DEzm9FXrnK8C54QOvVM+/jdKXPwCx
UeOKZDo0vo8TM4ibES4skK/rkfRuOLDRMwvlvTzDDqs0SomvuWWzFDIggE3eRka4kk6WgE7VI95J
uGUWGHeU/1p2W6ZsacPxmnDB04ABxbKkx7XLlov5U7YTIMy6G1RAg/vIet/XPCd0YcM5c3E61VHG
DEe51QS6E91WmEAdnNphbIJm4BM8O1V31YTeIFW13cHtkZGdQRrxAYrTI8Ch6OYq4YRxigUMN76S
SAJeyl/ViMchlbgb3HA8Nvhorklh28BVzp8BXcSEh4CpPmouDOs3DZ6y0aZBXOB3010xDTo78h1v
p8oowPXjhZNv6Ph/MHc9Zi7nKKBqcLZNpX+2YJLlPbazbI8b5tWlREwCdqreBfvXpKNbXbnK8WcW
9yo23pIF2yo3eqqsVPM/XGp9OeqChgDfGfR/ikTK/WBe0izFE1gK9b0gJgvb8iZ7hYoE1bwLgQF1
cCxPngGD3XvqSLpmC29AJ6Ftee01WfgJ7OrhqUMlfow1isHvrnDPVm8FrVFV+a9UZFVYuoUndkpX
sEl6p6d4SVKxfLl6mmRMSKETujrcHaFWpJgQ3eubEChVrPabDUUDs04Il1cuZo5wUxpAeXFBjiIl
E8m9LmDcrZTF2neWSsdxux74LEej5UYsXBkSpSGpurtrDazLlj8v/wiKNtnX2bw6Rlt9ngW+9g75
hurXPfG52NqCZHswsmkj9vP8D2RqpMqWfv+UnOZJr4ZeuAmTQ/iKQ2gDRbR6QtP4vAGTP0lVWAb/
gnrmqCbC+4smGzjE7DcXaPdGDp9jt/7FJXF1zXmarWCaBglGwh9SsWIGicbxOXSyPt2LutmZ8Jwj
YKb82lbBumKbXQ0DFzAuleyf35/42Y8zIxFYCRaGBpgSQmvNRc8H+c9ssI0aYupztoHixL9VnuGq
DRboNPmDvjQF8+o68nc5dUd78VavrklEQEt8LEk3r6bOl/QDKolehvKaAjmAQ1UkrfSNORzQdxnb
sn4cxMx8I+R/znGT74FRuEUeMpV5R2NyCJNnZMpyELS6uh1CpCcOBv3t2+3DqHUJkvF55S8zinKd
NJRTK+7m5VpWNlq41v/1CZsGf2EHOCZ8ZSUFe5LyPiOW4V04sT3GyXnacjZa3i6Y5BK/94icgayw
9+V6BGeq0wq4Z08ZZwDu2DLFZhqXajScrmf6/1+2GpK1/xvv9sjqftUxnujZwGl3N0w/nFkHwaul
D+9YzOMVQg5+1BCe8feuH4QW+eYxh8USoaSNADFLvFvL0ANiJuuMFWLpPiPrTIYy08KXPS+yHsXu
HrEq3/NvFToopssDqmZJMP8pNxwhSnb9qYJuEWbVxxLaF+fiIkNUDv5t0pFG4tk+1ajlCZf+epat
NYf7l15QWlrrN33yDQjY/GAjC9evs9oummdzVAS9Kd/dV+CTMEfBkrezewPqakAXN8JFKxA9EXCx
bb4AnjbQXjIRjdC5L5YDSc9QMTvyXFjupXGPqWeBz8T991rIHOBCyq0rHIDP+ATh7z13GB+gQPyd
okJ9SLh9jNBvq4bi8jb+hyjBgQKy3GC9AhDy+QXVdiGBR/JMaxhkirdltPsBNZUTU73PvpKBwlMU
zFUvkT0yIc0iP21vQE0JLXxTsN2bPaAM/Ouh1ZA3qdpjS71ykjpOM57R+Xijl7SPewFhkve/O9BT
/cMa8pcoaB3N671SFD489MA+kXJcWP/boOmdlHKRpEsmdxxbl3w2/MrX7RLVKP03t+41UYw8MBKx
1PgAM6gFdR3uVGiSkIpDaFjm+N1Cku7HvvBLafGdpq+jweo3+ZybvTFUquvGjIgIhhYeoJI5rqqy
8lHFWrP4xC0nh6TaJzZXWsfkNHB5FTvFYNY/eLykj/xEg9o/Yt2AK7iUZrMIwgaVy4z33CpyG4Mi
3dahOCkBf2tL7QayaByLgr30Lfwkf6ydB7tiqokP2dJw/RHdjenDHWAtRCBoeJDeeT8dM5Q6ikNk
xWJd5k16/0UtfHJkAjUpVdO/J4JJ59A2w32FIOq1L1TOE9ChXfNUSjC3Hd8XfAYJ6Q/d5pP2WFqr
3bOt4AMGz1WZZ8YIRnClUv5ZjNvcKG+qY8JGf7oKmK9MnT5snfxJJ/Ofy4+FtdZNnFjCny5F/j9s
jZwlMCH2WxQg/quxagJQRGExlwyZvz8EjZKIgOLuJR2TMmmN5zqDRuM5XKSCjpENsWnymCej4r1o
iFi6i1OjH7Fr/qQgrp3Tv5I/Ospz/eug4jGxoK/qAS9ddUNrndp16wN1feezI4Hpr93108aQz1yw
MlKGBbKvQud1KkqkqR0b1sGDkQVJCi0BoACUvPGx4TPSIAm8H+dATNV0es2dokhRUerZDJlXFPJR
CkxcqEkj7qMXUshY33m5ZvDA9rwpkE/Tzpua1gMZYxka1y9VPw4oXdVUNjPy/A8vIzVG7u+bu/FS
r61XrjNj4tBBYFBeiIQfG+hx+6XgaLo93+oaIOFOIJ1l73SyG35A2Svrm+9SGqHt6yMlCXFVl6di
e2LL76Q3QRMmUImOJ9Gtn1rXIkPRwmDqdBG3QEnQwq3ezlFvFEnC8rwA/z0LJIwzytL6fYgHBvlp
+0Quank2ICu0II+txny6LKaDoI3reREByorKYBDE5/qkxgicYgLTTh/4ANFA0dpQdB0ptg+BjTiu
lCm3AcSbxm9ezVRCP89d5HO3jetCLHcHLShkJ6209zwKjGcYXU3mYG4dWs/hG5kER16M9kHjeKEU
rNXNA70BOhuwCn16UChG3eBkJL3Iv5YfuTp23kShcjpkb/LRRk/xqprUC6uiaXxhYqkfLuf1rqD7
zS35Z7Ggh+07oE8Uidmibiypauqzdgnz21an+ar5c5Kh84kZf2XIMuD8KTXK13h8W/XtDbDv2Yai
Pxw6enVVljBna5KVPc9UXe25gLNBuuw4ghVSSn+tFEMPZ4/meucAQes+kMln6QJnbYl7PyzRJDcl
2dtuej9sQ84/4qnK8WJWFHMHPAwVDPIYRudRnck1I90V6IIq6GSw3WWXXs8/BPoYj7rx6IB0GBD9
Ek8Y3d14/hQYLMeUuGQLrd7BvF9uRsszfItIibCNseiScuQIccPAc+f2h6juwm9MD3zcMvhpyLFr
04BULbMn3Q6gzMiThtoOofGw34PswrXTJiy8KK7bok2hXNqQoVOPJV+WikA2iB0R7aN4BW4HkDel
MGbSkOWieKEvBw03WJU/h9rXuTXe7ZzfPpfqGcuVPjXiwVHzgLXaljK8joy37evYLYaDVx/UpE2J
UfDgrJ2aACwx+jMy4EdbnGKEOa5fdkU2bge4oabs0wz/O93PmWc6uKjyK7yq+Cy/WBAPifi2XQ36
NqLLyLG6hUd+Cftb5/jGVoNkPj9wK2Sr0usV4UyuoUB6XQVFo0Qs68F4r9GedLBR8exIc9qOgBiC
RGhnsYBQ7IvB8uVX2aS+QEDTd7FPU+i+z0tcn/oXG+jwaeXSDdKGKYDeIyZGbrJGl0Wk3RldidvK
AsvE9r7WjRXsi+Nywxzy705ZlIB/Xjo2NwHq9upcFUqjqMsgPbJaeVJGpvGnkc5dU8Hd8H1IKRv/
GgVuLR01EhRyiMNgQHnPMtfd/q86iElIPM7bl3368CZ4Z7FqoBEuCE80zT/hPOsEK1aq2Dd/DPFr
Y7r+9+K7EA8AvdFYllkKwdQm8v++Z1beLMjP2BcZJrHDh+RxApBFpwuKCA73c/vSz7SU9Tr7sPiU
wAqNgXrDRHBM7oV4lS41CXovRZ9GMbPFhRKnHv6iIQ4VD+09SJyr4jaumsusjFWaONrsswMn9izg
TJnyweCEl81KZIxkWVHq3Mlk8tdI6fLosyuqDoSFzDqedPKbWT4bQyyAPZ0OPQFgoO1nyAfELcaB
pS8NxxhCcQJAZDjtuZJvjkeOAO7TAwGQY5eDwrZHZpyHwZ+rVxorQ/WlXnYZpLvbgif83HNSIqnF
EslQxIHNeUN0APj5gEROf6hMNEb2ArcngO/zfOqP00ZE2xQFb6Fk4i1brWRIpThM4xkzgpqFhEjG
HCdQ92exsOZv50Tr8HvsNE+URGEXU/XlsjFHtL3vHj9SRZ3lnYX5EDBERBXxo877sDQ9mKtZ68j9
QnwG3hus9o/I92ux/0DiGYJKj3EOMmjHqdq/H5kP2VCDmj69EmjroOM8DtkBIZ7cvSL8IZOsKWQu
Hv0KkLe8bfJc32cJBKzCRJVTaYutcsYSZlMleMkuux/NOCGPAN5JymJZhlzApOHUF/XI7k1yB5b+
wK0PaOIZmKXlV5x38RlBw8I7b9IoeJIA6TzTMXunb7iOPxNMlxZI+NhhzxYb6GjV+ARQ+f2o3hag
qvOkB2TudvsBE6+UIbbiD8KBMPvVlwopVvf62kOPQe+tz3/ccUIQI0+8FBq0HpJ9CgVUJUdX6BVT
kzDQpLKFNOZjRrgFS/Rp+wSZqRaOddcVJvb0eetzLbdrsGTdKitvCkAQJNBdtNtMCMbV5yw8P4mg
X/eEfMtH2wRYwuY7w80UZTz2Nj+FtgvFWH0kNTIiGls7kGe/oAHD3u+pNHXN6r0NwYcq+10yAWbj
p5YcAkXdyx89jB2u8qD+k0zr9ynTu/ma7YyPXBBGX6budqcG0ycZs3APpHW5xQPNsz3VcRMAhKBq
zfCyuTVD/UdBqoGeI/IQdcMTK8LdidzyGWKBZkTUATnkpxSyUkjioPh0kblsLXAVjLOzsJrTN2xO
uoX5Myl/QDliOUJHNaEZX6ddUZY+ox5VNC7mbYAtrsaPFiPzidfz/b9qffIForskP37hhhGEj5I6
rX3V1NvlbgQPOIKEdM1HHU4Uvr/0Qk7uOK2ZbAW4wk87w2xfG2lUDb6IC/rqQvkoVbBdmkbq+FOd
JVmv8T0VFU6GnfMFNwwPQgBs2fmR1rqpSApWo7KtEmeJmLEkOOYUjO3RNNz0Olf8Thv4wjSPMasR
ItG1wBoHzgTeldd2vHFb3ZQ3g7A7hUNPNMOEzIwC64Lyzk2G4TVi4Of8ZyIVywdjOYY9ofDZlC2q
EvwcxDmUR1Hypu2DKKpL7OxM+stkjyuZKKCB3tRtwfcat1vGyhY8Fv0W68y0GsZOLzGyl+IZV/pC
SQbKn845Qdlz3/XTal4UgZdAKgvrvwxCkgL3yjto2/xkSAUvvs7PTUSfS3FWBs+RZ9SX8XuvNpz4
sbTJvk/g6XnlNzRJp129EALB0x6UkCAsNKGoi3CzdKokcr5fF43STViHHFUcjLRIBt6tjZJeTXXN
fqEq+/SUMcLCwQ5CbiVHHTdRszHzOhOzoPlJZqRuHg0XN4zil/DrgrQMiFkC0Olf5NM3VxVVaQYa
+0br7VQyef6++glD0mLlxSwSy1EA62Qt4V3JMVTkK+1jkoWozSd0hzY04WUMbRnk4VIFlRaJNZuo
s1FF1iPmw0yMdctCNEkShGAdaebvWEWje/ZCu3iqSuBso6rHxLL68UwaFxXLw4rUs5Q9J5fYnKvI
H7P1993tesy6/m5i/UTfQ0lvgf6RtFbaNwzDiXrFm8ePpw7vskVVeajKC8zMCMAyUP/RJpLtiWsI
ziQIqG8RMf8/339xKwnh7wlkt40qk5G526g4jjr6lBfEKTCr9ZAL+fwB0imFzA8daRf2Qr7s353Z
1cuHBNqqCMxFZuY/8Wp5xOE6CNdbksYMJIrq+4Jyv1GG2sw4qiOvNW1bnjpUzhARQqpgFDDdpQlm
DPCTxdm29AiPYt0EZeoft9M2hA3VX6Yfee6vfjJE7tzP6yIRfPkMxx0JWWHqq715XBJRqXPj8zdo
oD9EuDQ/GGG351ogMxbu2IBKVTwTgszEYMQbDuEUB2+Eh6s0ktSzXwugjpBOu+aZnaOwHNeKc8AG
n1UWaideGzxxa5wyGu+gKLyjbSfS2TbLqKUSQUwejzWSKDtCJSTkK5hPx9cAMHRFmMjgAiYUDnpB
noX/YhZkQ4LPglfgx2ihSAEn5WazN66PvMNBTphBCOMNPH0cpWdkGYxeAGanEK3otosGJQV9IG1L
U/p0jNbtrTc6lx13bMib0GDUVKL2At9R7JmP6OSZceciqwghlXHjhKfDz4YL0d/uP0KBRF/EJKfU
220u4A1B/+Tq9ihQ6MkEmDCYqZu4XVSDvP8Wh3NaNzx/GJqthMDlj37Xzpg0Vlsk/b/Bkn/m8Ft5
8qoAotFTf5aSyanCYqOdC/LPc0M5mG1Me1v+gufe9FCMd290w8w6qdU7zbrS8GyqmQ1haSz7myqK
ASr/BU15SpW13PQYJ1BH2pqNd01itoWEm/32Fl9J44Y/4/dKfy23OA55bG/h22nojzMzQQAbwWIM
zKMCPuowyGgj/YdpA2j+XyfE1EDCEQ06CDEHooSwrP9BOTIZXq5fGdUqa+OaLJwjk8luXEWLZSMv
6yCI/NA4RqjQxsSP7DyOFNTrsuC9p7UqzsQodQT/fQ04BNDY2fv1Sr1gp068u2JpcUht1M2I5T8x
+p7YNmKhPfDjd1YuVQiiYuAjFuQmz4QN2Z8Z4DE4gtD9LmjxLd2C01TXOStz6JgkJ+qNE/YPKVRj
DEXsS2ebMK92fDYkr3Z6NcWj5ogLM/B9+a7jCkl67cbeP5syj5OlDPrHop31mmfi1KxOhnQ05ljl
wmcpvTwat9xGetC+k4wbrvEiVuoWVHcNicCS6EkIIlQv38W/seIRZMlfC+gNZW9hJ4KP24G3cZkG
k9x9+tbSWJ8EfJhOyy4Y3/JRj3akiEaSXjVbIvz3pguyHsqYZrhtORNtkMg19hY3UUbWQteMlKTP
X3QyV591DsMm8SnwhZA05pMLRMC8BpCHc9JyjnVRr0CZJmNjyG91JITHfakTaquGPGmwWYjrRMol
JUHoBZlDdVbuPHfgu+e3qU4xBCVaquurk4OL8kJ9rgB2XZ+nNNodfKCfEPVyRcqeRmVvIvaFZM3M
GPn3p01tKofcS89fERkeIqHYrPjt6CmAdrAJKo7Xvu2boSCpotF7A4raCRQtZmO0qtvQ9xdhk6z9
+B06+R2lKxpJGBCQbXg9hHhoXatR+IhpqwQiIVd32pHjBW4TV4PDE9OA1F3aND/DDCRrFNCTOHEe
PGvsKaczTsAsLBL6mDfQRIwhXAMesBKxqdKmyZrz3iQl+nxQJoAgvNxRdP3ur63dEY3WdYeE9TT9
Yual0K0jjlxtWltE/kerPmRGY/9L73cDpPvrbSNaTPeruxh9CZIWYcTnQAGIsD/XUeQ3YmnrPPp5
u5fr4G1WoRBs8itrA9ERuCHLi9yvfNF40QrHZQzz6oixKRaVYm0su8eM05rh4IUkXCJKFzFkhMjE
c2bV20FUgXghq3ZUFBxvZQmXcufzggQnw8i85v+0N7OFGwjK7N2kCWs0MeL7yaTBjOeKDQE79e/Y
bCBD7ZGuB1UkIP26uggSdcRNieesA9OtQy+tlw4jGRmIhCu0rxdyPdb2vIR7JyHq5tCmqe/1osls
sY57vMo+6D0+Jx0FGt6y4roQRetpNBESqLadpW3Sat8cFojqexp0EaBuhAQGjOdhW/rY2BEbWo4d
LUCVebh3F0gY5TMcLnHFId+NNENTzF80UbpeecB7suD2kkRZHCNXtyYc+Z1xR+/5atdD9LZSA/wk
fWBo1fJPWZhSjM/dh9pe0a7XE50DV1NlmPyZLcbkF3l+oSAYohD6b6E52ounT13dWj5Kiy+9PAeI
iZQporhiYnu6ZLYaDI638bKfYE6632gc3LNaJ/lbKud152NDp5yjfeNMUoK3bbTYDZ64o23XMwX4
gEaPYzDu8Has7kHGypmkDJApbksVW/G9zsIWYZVt8+lZmPHmFr1Te635NGGQdxQUZNI62YKEAVJ2
6tmK/w5Mucbpkp5Cf1lYkeu/xWNbVTxCUT17Db8JlqZN2gFHegob71Jd+8M4IqxhkilP8gVgAZE4
Jb07Net8n8mjXvDbpPKONnuE43JBmcZ8EfUwk1hNvjl6HvZpeQxaIS0491tSRUFt+toklf7e1HwP
eK0fJdc0uX8v48ZTFDDabk4YSs95cEK0sqnyG4NJVhrDjN+PX2DpQdNp+06qSY8xupLtQ79Q1akO
g+UZlcLNnLP+P2oI93eaxBC9zgU6Rz+S5rbUeizC45uF+MvXaxcwV/S9FlYcxbcW4D+foknIr8oG
594NtWz9ICQg7E1qijQEebBXxPmreWYuV2DY2fFqkzhLe9+nAPkLJbqCGAzw6DLKXnA+ezNxjLVc
HRxMO6EJrBzhzTzpqCtnzaWUvvE8WwhhyntdLr+7HpVghbyhT/HEwf1/1uK2bkJBOTJ3qgBg0rAS
6YhQEf4i4yI0E6A6Fw+d2fvHtsMsDOdO1m3RNGkx+hH0iqWYrHpwTPsA3nZunA7nin00EV0bQ2r2
K4l9S15cQm00HV8vTNb2513onmetOFYBwdzK+uoRzmQeuWH9qYXd8QHUXXOL65OSskxhnEejGte1
5vJGnJfwgcHqZD4mJBwSttVv1MKPpNoweHowFZHfVZhlLL2TtSdcI45x6WXaDGOb+e83MPhE4Bje
6lQ6UOARvrHI5pS7UAwHlVuGurxJujc3wqrCP7hDUlOawp7m5wo90OT4UIgIQpD357L7YN/ZOU8G
Q31TY8o2GQyaMy2R3YW3ksd9IhdRfLC68/W3swPKaSrJnJ8GDG9MrrVcUenZh4sFv/Cu1y/Ag7LL
fPBnZjwsz1vUJiANH89Wb98D9uQ+4vrifDHWm691ihAfSHjO0W/n7YfkBM0rh3cDpzVwiB5otHB9
OyUHs5qUZUtYaZSJWlHJi4OqgtBZyRaCGOt1YSmzNgkaSrxIt0ciuZHaTYSvnGRV3UTzFuUZOKor
3SDioQl+I8uQN28Xo4qOZRwlRekxUtuhk7NNVxnHC2umByWWvaZLpAYZ7teOZORtxY+clGrMntyu
zwdhGam73SloUhNNThwCdTz7AUpYiRxenajca/ribZjltzsiz6nkTDJtKqjGtrMLUG9jGvMqO6r+
lNoY3VgKODLrzXp/YtCGGl1YemV7C3ICmafgzmZXZtPyy4Y0nvEDTlAZSLSc01YiPfrd6HfhHATg
iazgityUKrBze6xXIIvRAgmMkk0lpvxdoO9zGKs3qWMUTgkwhTlE6rAXa30vdyTh8JK5m9e4IDIg
DV0uwGoybPhHWNUJQklnFWILbV/CneIFOceXHazNW7XmYQsDF3K2bbT1E0K9eejAesn5AYD51Xze
Hp1GpXNXDLbCRToP0g4twHpxjwBFk4cQYLVewzkmOCSqiaq1a4ofD9VAoaFdebxIdMXgzWbVXI5N
rwbMIf4OV+uo2pQSdxHrW7+Bb1atuaS6gnXnKanKE7RroVehUD9Chdv7lTCu99bts4As9WsFCLK5
BRSP2TxbWQkarNIVm48CZYih1nB/Hl5G7jsGxd87QeR/VzIaQTswg/dYJ2EL5glOT1X0Y/JSDsAo
a5Kk4q7s+S0DfN2TD6LCudffZt33ANRYnedlkKoQWWFv8W1DVvkL2qFS19z4VMAnemn/+fLTmHim
E+X4MC1QzL3KA4m0rC/BXW4rPDczcm0bG3G54AWooFW4Ev7I34EuYjPoYlGVrJZyvZyV1ux2NNnZ
+aXerZGf6XN+HyEM5fI67fQW79BgPTH27n6dP1wzmSTmiyzFKdaRltsTGmo+YWm1Ci6YZpCAgDHs
uvw8VLPJDF2VzgISOb50ariPSeGvWIlK22KoKHYBR/AJfJwiJCkULIzn14ictDOO5d07HHDWtpXc
/DpmL6pQXrBv23NlQBjzbwPivudBP8Fsjf6UbgthEeGXZ1+gZ6Jb6fiHLUWpXMmjRS4Pyp8C0vrj
zG15HGjJsfqQmt8t3do52xNIf1yiraHaQltSxvOgd6SLQAbuw1pzlTdA11nWi5J+di+lcRU8HkhO
69tt5Umsvrcr/BJsKAHQHq46Xtr8sdqoyQ8gfLAXehiLAW0/jEUMB/nmpQt7Rv5QzpbDwPGmqNT6
vdXDr3RBdF18OQidfNz+1g4NZIKE7HjyQz7uWbhCf7Kva9dGzNMZ7jzVvwemD13vWiMlharaQ2bC
nS+1/ZiIhV0RhTgSNGdfRbEf9kIb7g22P/gsQdiT+8OxKXrudLhyZhqFT/th0sMaIx9+LmPlsF3r
w0VnZW+FQiemBKslxN/1LkE2IZlQ4OGeEXfi6WAVSMzXRZEoDt+sGUYMS7WWCBJLhX8DERj2fjpw
YEpMPysbN6syxWXKyJhJlB3PyguXviN0wNnE2WDE3S8fAG3NrBPuptms8EiWrltpmmSaa3GIyUA/
SdNQCmC+f8CmHbaO93Aw+VNvr6zLd12FGQDYBCJipAOmVPVeecl2STwCQCJ2gfTq4H4R4KItkCgV
O1Z+wN7wMfVu0+d378Rp+KTapXTYDAx9ChongY9wfcYe5QOfkUAR2CraMw2xJ66/GXCAzu9hhZia
6iD6WOAirnugdcGYS112ERNBGIiP1NrLte6oqh4dgpXiNACb1WuB52gT3LGVBLfAmHk1+6Ed97XL
T8tm1vVYxFa9bNVwEshDt3b+t7SU+MNIksxktJr4KfzvLdNhiO3INwut5o4koY8H9Twmxrw78DC+
kOB5CQYIGgxdYtp66WkIOA8WLqpxs67fYEIwHkSEAstGvqQlA6EoHfq48IsJI2XCcbGiMzQwzyfX
zVy8kTosc+DMAhQpIFNtL9gz2cVwsgu7Z1jvJWAs0cR72Nl7m+6VAoPP0/3wuwwBpOrSSRG4eyP2
43PYLDXjChNCITTLu8m3LBwbFWypBVzXGva0yCfbMJv3d2kgY3FOfHn/y18uczdJYXeqSArTMwLN
3UtAXrjyZqFHlsft5Fx0Z4vcYHJHs2s3L5U21XwuJvDdEn/AzHkFfn/Ev6s77AtNml+T1jfp4vsy
6Ip/ot7igRDkNGPS0B7XDP/bOy3dD5rmwqCprBcMUMIfZdevSZtLw3v4hgN8aLR8CLkWNyHn8v9B
AoAeT8BNHw4f/YJtxbLMlS/tPiLLhjv7guyxgyyHKkx7Jqsne84RsSPeHdl0MVaJdmYab5OvxQOl
OEILNjbVPZnauJSM0/0EUtRCxs/OgTUrffWAfIDhNhk7W70QIarOEgQEFQQ0KVxn2X5qcGxhC85b
cjxTxBIUKo90CBrf8MpWOZ44AAus/xpf7PIWP7/NuK746M9zVN4zeETlO3Ai3loJ7Rue/DignsO9
9Hk8CfLF5somiah3eoOkIsNrr9w1YdmR/BDZq/KT+Fmkhx5trXE0ebF7BdYP94N2xkX+P2ZJCfV2
S2n2qUIl51lld80hFbywlcLBsmx9YlxlE2iSPty/Q7W54GQVF/BezPKK0yu3BWfELxlB+RwxXo2w
7k+1FgDxRml9+JPJIyTO9fg4Z34LPlC+sGAZZ56sEnMKAmyFT1krmvkZBZ4+3ukg6LQHRnb591Vz
THVpbrfpY8yFf5W1vBw9QBgiap5URdYoCTGjOa76WNPe1eJmlojiWydcgBMlhjib1vx9QRVlcRri
f1aP9rKv87NCt0ujfNBapbpFxDnBMNtnhRTLX2XwBK7kJ575E20W/+m7L6EHOb4jT94EAdbkATN3
jSMaWNNLzjqPiwHGs1czFHI9HA/nWE98yk1KJHUmqUgJlnrwLDVvMBkZavmiq2ZqG3sxMqrsu8Xm
KfSzhqHQss//BRepKhZTB0X6azKdPcdwh/nPk0CIQm9+bGnIpcNIP3HcLXhtKKWXhgo2oJ3Gd+tI
+gkaJ6sROK8jilhNdaQt2OfcMsMjBYCpWMiv+97qYU3KNDuk2ZMs2HnJm/k4pJzwqeKqZ+ykT2M7
Wr6fUKsdbh3kAEUzdiGtCdVRRLc8s1/5UayAoR25knniHJdZFTVO8kHsBZzD/JrEkPMYlTNtgO47
i9ayqfEoYJ0Wz2A525LqH9XqKPFz79OKO4LeuK6B3Kwv+9pVeFSMbKEiVQvDULVSQpwHeKDEZhQI
oWqBs4dvvrKfnM/K3oK3pzRkbCH1g30DlfEs/0Ur5fNXqYFaU1eeRasaI26jxmY2POzZFwhh3InU
9+4uNFyaUo/viUNIh/xruWMKu108sqkMWTX8weHaF5d8IYZvtftH2zPPDJB4SgyJwWk8EQycpIqw
TwlNY+1nFgxhIkIkvFWbMx79ruPE4XZIN55dtpZQ5YtTyzG5pQ51FROOSS+NcfWwoays7+9emXdO
btCWX0RT6vTFkxZuZswmbzgR6P3efIuOKGQAoFVGdt0edwB6kFTxFE8ODmzDjA69iqdBXqHB9BJa
p+UXcco1SShPwi6r8X2mFPrhjZf8dwJTxl55EQeqR9CykkKk+vKtG0TU0rNhAirYsvkyCYhUphwy
eIKPiZthCyC1Yck9s4yHRrJo0+DFgoluEeDn35CTWKvXfmtmWaOf04WjHDNIzw+/yPjaA4n6trAa
sBwpV1JAeuDB4y4hicXorp+hZ5XIgFxtbH3Ah9YCNOX3TeVETUU/ejMWVEM7iadtmW5EHrXAlwbJ
vJuolPZ6gOF5XNND0gk2v4vdzJUtvc2uvXhGj1jHCHtFZma7Rhb+LqWaPppj4ANQoHmffOsBkYuJ
92tam09vaV6jPYjP+RUGr/JMeujpled+iLjWlQUpFvZ8lr22k0ZhhPpXfCKhv0EXxC43AE7Z8a/4
Khv4KHPW9V00Um4BQw/7vGMdtV6VXRr1YVqSU13myAHRBoMpCYTNf+tt94k0Nx90Y6TAChr0GhKE
AHuuL+lPEl8lpGg5Ch0rfUm+MtLcBKULsM404HI0yqYo6DL7JZgpVYbKMx7yAD/lNYtQTG9MC/qp
SKjLXKdn587MiHW+Nt5Y820n53e+J//L7Q1+3fu64bDsoAxdLAkrngX0PbAggcroFSOpbifPjXAb
wt1DPz0HdMIkU/wl9VzhtbHkfbw8iHaqiRDfM2Dsbn1tjyHm2+iHEoxzrYUJY3efJsBEq8+HADwu
DvW2dnMhEeRrlTWbwcLwaxc8SaEDPxBiFAifDF9L5pDrlzUG4YX4lQTF1AO2cBvOeGfXY8SoFCQ0
oOsXu0OeK8S7BNpvo5oRhSQbbCSh7IkGIqRHaqmvv+pd4IJUP8M3LiVnLt/a2SUCges7dvVJYqe9
mSpQ7DjefZwqbhWcJuX0ZunKPAOFKC4t9uLuQSZYq5X7+yWmFVxtVfJ2mvtptvayog4W0R2rK3bX
iOGQpnZFCgM9WBgObBLkJS3F7em7OSXwZsI3n9Gy5Vq51FzCrcX26rCvbmfcXVfjdKGTPT+9SnH0
rVROVn9ccBAWFYTLVfhrmJgzbMpixabTQ6FVZQ7F9F3gIc/QszozJ7bequVLkxfNHsZQVUZSD5tE
+VPnPXSAD68Blijsir2OcxR51vGbp2baCLBvi6VX/7iReOTT103TN6Yxj0NxF8Wfw+ILpxowh24E
XqJpfVz0PXFS+LwFL7CxaqvdyKeCtBK85aB1XgJH9LUVNSOVLtwnuvn/nLK8g1zlu6mz/W0Rb3St
aivo3vxRvw6rxx2OWV9YdKFRoTODoVSZWZKhTH4NI3vZjfbGUeY5v+tWZTIUux+KprSyecRaN4bM
Cx+NZ4DsJR1IcQ9ls6v/Z06KgXxO6pg/iOGhgUwnDYCwN9tvntyPW5Tv+ymlbS9g/rAtGUpNRpZs
jNpb9gNTAOGsR1ZyoioLhzTbB3fs09VTPbyBN60LR8NCCLA99C3uAUDvEPPOcSQPyxLpNuEy1jr3
MiZ9pEHxPFHdQPvV6aEqmsBuUHRP9AaNbEM/kv5MkUH+3YTG3fZ9BikhhvbpqrI/r+v8P4kj2oRe
DiXH/U9zDSxXWFplIRhf+Dgfuf3MTrxk81aATPYSWWI2mocFUuJ5R7V2lJKYJE4R0C018t5jDPKo
B2bY6KFcOEa6WHpwH3d1PM4MLj5+UFOFHcDNqvUQpBtGpVu3sA0TlD8VisAb6yyuy/HUMVoQIgyW
n/juTkZidophB85PThOcn8/WBg8+3P8YQ6k4tM78PgRsgcZHoId3o3+9oFl0wwb9i5FCiL4VHs0n
4Ah4/AVb+JGQlMQPEVN3+KCt2EniPWv8IK3QwsTVnL8QDYrkEB2YBweRg49tUCkU552FrozzJ6PH
/05fem5Ir8urG2NBbcO+hwyD99e6+Tzt+ljrBQvFSR0DxbIvtxI7jY5mUvBjpCrGIsHudffFv5ue
IT4/CG4YzjuWCoQIeN529YDW8JDGm74fu6u6qvw5BSqFRoxF/vX4fjUd+MDsezVvJjeZUgFyXFyV
E47OiE7kSWY5mcF8WwL7lKAp310qwECBM6RzasgRQGREslAPx6v6AvfRZrXzJ4HI8eh9uXeVGPkO
4bQ1b07+MfTC+LtB4eAUvFTO8Y1K0cjWYw7hkwRgEB4qJw1mwIHRPOT8Vl9XvTHBH3isWWj0PSVX
qAwEMoObXS3bgeQCiRKMjCgMdQc7qiiJNjedxvfxqBMtbvDe0ZGyBX24JJJwCUwEV1f4Qh5YrRuS
y/VIaqO38FsjzDI7Z047L4eJ26eI58ZfhBCdHbqyYt+pLNDpjdjXzM7+LqGO/V2yHRTaR0aQgIAv
rZeu6TND19B0vFff3UYmvmAGcnDAzTj6hbIc7JL6PevKD8fUJZ2KIFwl1x5Onu+/s7HZO3fA3AUc
H3PM9MHdE6To37acJO1mM8vjP9h9Ajv1dH0mvXmLraLBepMGfZSqBbtVsk/1C24OrxnLs0kuar0j
yqssRSE8mXyQLqQcDznJAES+6/5PYgdHUI4IOiztDu0hRnj2PJccZeE9YosodA2ou2aDIc38N8yY
xcff2P5zf9zkx9fZ2TCxJwQU/gz9PH5EhF4net9prHsGpYJI254Rd8lPPAW6hPhIahTTPpF3EVHM
D364Dp+1q1jizCTKDqtgvywtGqVyEjdAQxKbiCZ1sjlQomczJ6owQVTcBOzIrxDKvtC7rj1E04zA
vtp1EovLch1SunAk+xucvg7LnOv2xOjgE5Ar4KeMWQ05FiXIPZ7P2g+X90+u9vDszkFjnIxm3lBa
jpf674DrT5j4RYkJ1CdZ4k57fXsBlC1WfZx8ozHsIqzD/3SgLrsEwNpJw4ht6JyX+QdTE4pvgd+V
qDROjZEj+00lXuqmwUWT66Nse/V8g/KVbjZr4NSyAvPEg0n81X89Yvfby4xJOhG4B+5wlUGa/Buc
uuvclc3XC5GcyMiYRSbqcNeLhTTujO8CsK9+OixHXLgctJXX+7fqwJVjevlUsVuPJX8K6Ff6P7ui
6DqtNcpyIPPTEy1Rr6h7mOqiMr2N8udfvpNB4r79L67Q2Zz9jz4cXJCgpg3pwr937XvnN5pQ1pjR
CVVXGFEZ/aXnRCoxHMGU+/jHSd068owlyyclaCNMTbFpSQD21LkvS+sLXzsLEttIaUcHBAqjoIKd
Y808EvqsAlCOTmtSQ7P8gZV9TBxaDir3kuzXC9MAfD25WDJQzXIIyavgT8Q2ZTg5WFHgV0XQQ3JO
kVPUPXX6H5kbVcwHMC58DU4l7K9MceCjCtsYwoPr/tbmNQhKeiCHt6537ng2XX8YVz+4ISqRNR/M
OeKe7R1TF6gBc5jHGF74ELA4cEwE5zZiMvLrSuXzbdumfRfvTr5B5bJggsXJqColmeWp5rcPaEIS
mv3g8p3LKCI1mrKIdwNg5mp7QSGRWBgtnqfLzm/jRjF8lhIph8llBvnBUcyoq1Y0b1yg2WFBAguS
9kxKqV0qc6etYUdR7XD5jEzksvpZLV24k+WhskzVBT/0LfNpKh9hDp0vTxUG0moU782NfC/iusqw
8O9jQb7hUWovWtj/gj4sOm6U9lyKnNX7PGwt7Q8BgXOjPbJWhbYOg2WkLdjP47R0pxZkBroy6cPF
P8Shz7O2sD4uvfWGP1hv6ayF03cP/cCGUBXcxZjZgX16dnDT5ibaXYM3HjXpPOfUMDC+qz3UwVeS
1hKQ8/HYGplTzXlT+97lyFGg8AOu5/4ItYoMj96OQr2M1cLZIJG0wihpw4Tgl5CZSYlTYYxpE1wX
f9LyoG6/DvHWeP8a3zeMRBlf59g5avSgn9tplDuimt9IbFGIQKw+l4NyVuSe/kb3cn4tUbn2cUXO
rDsSDwv3WmLx7JmupMpz+aw/QMDmmJBBvGxD8zCOfC3b3WZEOJXX73v3PiZSCTSTwXOdbEFr3dlR
0SLbtmK6D5o6SDQfsziuBShzCI3Mx+W8uDjH0mTRFjR5ylbGpWDEDIaNmNrqryZAgoxkDDXq5hE0
JF6mmT3epkOS88a6RIFia1wp5eFIdCHOszQFxG/o+dMWqpgWwcRXIVcQpcJVSjxhTVC4eLL8DVh/
+lzMdRaS/iXEStsr/2qj+fCDqs2fCiaiFbvHXjya0pGLmnrw+aiZq+7c+zBFfm+vsWysIBj67KRH
tmctXpTjFaecZ6RsbO1vTIdXPQzeJLpUHHLNJu5dUfxy641OTzwhsoIKRlsKPg659OFj+khF9fU6
+7f8uUvZBUqUISFN6InQYFghxBrF4gf0nv5cubE8EWWAJuErOCKzMTDEne4jiNus4JH4y0OOHz7P
pFdtLUpHWpEIPKb/+fhFzt5tfM4VWyQ82vAYQ9C0a7uoPMWV3WHnJswetNQZl3CeH1EnmUJFS9Iy
7dSo5MRcRoccz2SGceNBz6ECrjb3Knn28bhL4gYloWZ1zY927aZ2A7Nk8/zrLeakayAXEOM5nDQZ
cPlzzjrfLXv2aEg4irYjfmt2Op/weFOl63q/oSMeOd4JjRZzdve+ek08Als0AvpuVY1h1HcoB8Tp
BqZnVHlVmHwUnOBG7LzKHqvbyqswLGVfA8Hu1WdkmtnnnhzZIEYCJaUnAychGPHB42L9+QKjySDj
J3+N8wx4rlHYFuBrRTg/CazUW0CuWpfUuUzmGkevJPYrZmT+arUE4GX/NEkkzEXQpwoiotvf46YE
qy3Eq3HLhGjSE53Fju/+T+HdbQRdwsJRYaw7trPAlxe6bzsEABsicOYjGHdvQdbvY/BQ3xyIcyLC
wse/uJMwdljGaD7OZt24oVsPMf9nsvv/jxjPFu49KfwrA0kQjo30nFRBlohxv0zhrQeUUqSepzVU
fKmiCpS0UIZR02K3MTSw8ZV2T+yrsSE2/aApOUw0eGuBWRjEVgfygpWosqe12mkxRPOmHj8fMwaR
QBxQAYkjVOi1F6goLJ1BT5jAZDbuvvtnpMlqXQLweYkN4V6yZ9imfAm2nT/W08o0wOVWGRNnWRw6
4lYpKg5keBx+z6xHBxOR/skOwYwdn7qe7lJ9yrOptmDCmyR1IUq4vTRCfkn9qD8sy9YnwEnvduN2
iRipVh9EPNap1b03GXq8T2AW6EzzU8KqNNXniEglWXMQWYEDTmSAU8E80eEq8Pdc1EG7oz6asAwL
sjnfn8zguFrXyow7J6d2Ccq1KllUD+K4lTldgqSdvclpQp5eOWK6SE/jGXnYr2rzhusiLar74L52
Tq6hp9A6g0WSliT+gLrVchKHLOa1UWGVe58l98Sa7SOh+EPh8MOfdMOAV3brf5MbnXMCkzE83kia
QLDj9hWuekYHy498e7R+RqSu6NKstH4yGm4pxekohKi/bI1PwDVRHjSQQBE8b4FHTSFKI/XAIrBy
gYrUaPAOKNRF/aIbegOLEnTLaMohlnPcNRfg3uGz4e6U9B6dXu1q06Qb4F2+/rL11qJzP/iLfubY
uCsrYr7CpJuJmOaV45qey8FpazGbKsSbcg36n7FCppO3Tmyj7llon+tkZeh1N+FLzSXFKwrtOZNB
BsnlJNBuUPanYWyKqVuR7p4bapqZEWgM+3wGHd/AmkayL8KNZC9WGrj3KpNtcMn59Yy2DY5N9XuZ
5NlCWoY8TIDKbWaTiozkJenapZB1gKr4KJyLYISBEFosaKwkiS34RaX0/MqKVxTe+OB4YxsDUIOJ
J6jBaCeUVqgGe/XINYgrv2Kfyk7XEaR2NQmSE/n6s2C6yG8EpnKMwqz8Xv3LyGhwliHthwFQQZmf
1n0XqXC2/EdUaXr4OfljMh6ir31aXQLTYMwzLPlsGrH4Mv4SrDuSI2hDkB6ZIHWkOxhOPl7g/iKR
1XxTfg9k52F0WXMA6BPJuM0tV+K/PGNiAVNand0OzuuftQU5MkIXMg/fkHLEsT0tsCy/IDAe5uXy
xxm9OOrYppkIssr4OilfisjrLoE9Q/wVXdOuGIsojuw5hZHwcwLn6/pCjbTbmdstsQcbRo+U6T7J
KSnoVi3SlCnmWbet2wBAdpFBsKvKWp1InnqnY7aIRzn6qb3Yrcuj1PXWAuUmf55RAPIymZWBeQRk
fkh6+Tfelre/4G/qrEqydp6MCB1QkYeqpZjWc0nn456q1jIn8wu7diHZ85cDqnrsvtNW+0CW86Ps
s6VATW8cNyTICC86YLT5ADi3aNP1Z7EF9sLZztDkOXgiLPQ+wHdnVK24Ru1FQBfgxBcVi/Iu/afk
HcD7Ml6TL/Rc9CONdRUy28OPuHCrVB+b7WwcQj3fl11NmHrjb++D8yX6o5vjIwquHo9vUtKtF0F9
3oY0h8HcB86aXMh5uzyA8F5+sBltRZETveQr0ZFmpunaabebvx8vZWR3nrlr4URRVH2H8UoPzsdy
PeqBK8TElikbzOUAznhYOPRBywu+CLrY/8j6slu1v1EKiRPWU/syUKFevQ3gH07jBlDTUl5qjrCK
NJD9jOErAEObc/eTHdAc9vTPEn9dxLIzAf+br0lQo31Rv32eRp2O603wjnAuZB8OJuC3y5WJ8z1b
ftzY5/npfan4HfpHklpuSZrFtLGRVbpzenoDLKvTsw7d7enmWdigKPigDECeSukl3+x0k5FtxjSc
0liQJe5LH/OF1Mg4JD1v/75ntmtlrSSoH30kdIkGZJTADc96pkwGRJH2l47aZdY6mW3SbnjsyM0Z
lG002BEHZD3E7VRpAqP7pDjmm3ElGQ2HaFSmNMkxAEjDjUa7C67kle04eJpkz80j9sKG68X2ZIM/
it5ZB+m8yEbfjY9ASz3asgyvuX1pIIvhouSqWkS3je5LOaZj9p4PYk7a3u/LnFMuUCB124AahWsv
Dc0ktukz5Y3riaPdcvt2PBFGxWzPUYBZdWfTlV15OXxnCQYiirJagpwAoPpwZW9g0d5OqaJwkYpG
Id+J6TXn3zGKY/IGye1Ms90K4R4CPvFKFPe86urdddML56BQyUgcH/Vuc8PTiM6Ll/TjnrQa5qH0
rijD6fyX6p+rZOY8EH0kkVeAYy50AscXxNbFLemwazTv+mnqVH8/6+940yM4EZcozja6LDvApIAp
zvqyujz1cVirWaDEiqiyGuJJsGBYevoSuUpzr2OIsSarHl3HTQQp1+0TPLBU+aG7+EUQgEsNhTrA
ME1J5T7kVNR/B8R2fNQVSsnQ/jAC6yrX/BcaW99vjBPFzqOM6sMAKrGOp6mI8sPvhK3vwNHguatK
Vo6GiTzAF1NTXbNQYp0cm3wZSlHMY5v8T37kGLiRE/OXw5sEVPY+9yOBKTep5lWaAYv0WPGgFLQI
rNL6JAMix9abe30cKfeyBP6GYtB6zXSsP6oonaEKZ0Js+sDFs649FbwuOInDpClM2G8Nozh76GXt
3ZX0Hh5BygybNQSq7q7vhaxoWCaxrb3TvBDdqi8w8ozQkiof3wL8a/Dh180Q10iiYTyPj4Y88dAP
4nsszSMCzP+k75sjKWL6JCwsW5yMaKfo3bzVQiq+OwcR/q3r+v/zzqvJ9H/r/1e/sbJz3suUQCY/
LvYsT/EEMbek+mkyIkp0yPMd7HQwd/PNFhlczuFxCGSdD4hJpgVN9X3zl5InNNncJR2PP1HKAq2V
sMDZS0+ZwZP8iDz8L4MqElcNwfv5GbOHDrdw2KjnYG+1PRH9f5ei5R/4vSMKhlVl//sXwf8DivXD
eGyIgpoZe4gTdyl9fpadoAt59YctDDiyYHTyOYcZs41XnPg97BM8bRfRziNikk4wu9aRs49gv0/X
o5aYyMktjhx1NlTL9AxyGUYiGRRSgOff6Qr6M00NWohzluyBSetoL7PQBR1o0C7Le4GcRnkXOPWU
1XJw1zqGQTLWKtOXWyv8mRNC9crAqx9Q/YLRoJzFAqlOpb0n5n0rMHjdu1EakSePvULT8zAT1i7Y
4Jqyb0zFbbJpGtOo2juF4jkOq9GWT5BBDBVDZvwzahmw5akInXSNcbUXD3R6ApF+Zlg0bBic25cg
HgbeFx45k6rFiOdjqdmg4i3y0Yz40+KV2gG8GQnyt3VRUNkOp1X1xxj0DNdeu1t9Cd/gy5XFdO/K
X9R6RY8I3A8E8XOWqHzljbIfwvHzkiosDAFBIVaayULJkGVJHpe6/H8qakCWWVItK5aoCwKCTs/2
Xzpah+7GnX6lGWw14JM0lsiAZyLqj8vbfUmllyruHqPuS4i0Tc+Q7V6bhnBnx/bzZnLB7r9ISsfQ
/wgr8272M0gu2tBzYDiCuAObzMBWkciciruruQ8hbfIstAGWMK2sOgpCL9JJcNNKpF0UqSgKFA+w
Cet8yhOniIf+YSJt+zKpnvLvq2a+/ldOQ+bMcrTaWbk7ZadpUOctmGX8/bPQtkdI2lXXenXiCgIJ
0YKNtKnklYctVqp8wLhZ4jKfkD3sS6YicTK3SVVMmAhwBjGLW4snQwnUuxgJmkvAZk2wEjZwe0cK
kcLHScpQa2+uKQouptHt3g8AA+eKUXR+597rApCZHUmelx1XjrI1BEST+4Q+GA6fobhWLNGcA6gD
RdBL+qzNO4RRugAZ6pecAGSSjMqLLlWzNziiTeGXmnGUX9HwHPLu4Up8t3Qj2RiVYdyXc2cTwlvR
8ylTghWgEdx8wjvoOGWHXMs+Ch60X6p7p6coHsx3uZTKUrlA3nAELLKd3tIKBOVp7ZIfnV1SKhsq
IE9tc72yZ+9bxBAUC3vYMh7cQYIXFurD2LxfOp1OET+6ylOaP1MSTjfYz6pTN0sE9qmfPzyGciHN
XXlvsINAjrGI5RaJcwRZOTHkBsV2JXlBSe92526BZ4hWtM9C/mSAcnQiXDtKA97+MMU0u6aWHJFm
oWRU/cFtALskLMQyBRJChPPviscHb8azbs/qC9v3YoJct+qdL4/fd5hfGCQ4fLidQSqXLEmrqnIx
H8xMM5K3Ub4lahio1eEzIpZE+ya/XrroPoq/78lQ9AXd2sh4eJO3/AkHvGsC5eZV2l+e/E1v8jGb
hVBh8XEZmvvtkmfRJTNkMCaLebDsOd+aA0yTf/9QVlGE82DpZAyyO7+VB7FwsNISHOGGyj1eGjFn
yQYvNOdi2XCg07utWeSJiq5xUStSwuLLODnbGt5xOFPb1o3849yJ6WlniNypzup7sX2lfBd9Ls9I
IE+7yO+gMWLA+d4nku0oYxRdco/NmVuvdVjTrG4RkeDYwKDK4RjIRtsFpAoGIeapS/tvBbiuL11A
uoG6/K4PY7eFrY7IG+qgj8qxl4XeGxNkdGPdNsiCid1ZRFngAnXk5w8OBHPIGI3Nh+21ORgKSWdM
wjSwfJ/mLdDwEtxLtNP5YPiJm113JpW8bzl6eK28dtFih/EUyXVkwhFtHPQoMxidXSdjwVyOP6gI
Fs5FXQ0URf5oBEfuNnoDB4UW+r7MpOOWL0l9ComCBmy4xXEe0eknShMWNLB2F69rT/iQx274RVGf
YLHmjNwdCEykWqPebPh/0v9HCfBVQiNFccDWwF8k8sXXLq1Di8t6xBjMQV5EGB9UeDSWdt4A0DCA
pqr4E2szAtTqInqy4NRFX34jUO5ffFukkEQQJHqSC9hQ56WlX7pZKkojbI5tQg+7/S7unHO/Aqb/
GA0mIHdlhHzrKoPIJsfYwEl5lWII17jt76ix+Wk0Gmy3/2PRyJlszWBHqi+AiMO73cPqRdHuK4og
mn5/Ml1RoURY5ers2IC2hYPGpiq3W47ZTnjvhTVCtt7ltuOik0oleUJfVoyJxnaoXBgxxahm/g9F
tETKBLbo/LdBUD+YlmX4sBAsXY4vz05YdK7+Uz+jo2ZJLJ5r94/1xzsZzdJfJAgyvgS7Phx9Vjjc
ckwp/ilMI8UaRRQWlLPOZMl/70zrLyG6TDW4ID8X9hGF0uW5m3dAclSWz2mAb4FikvDDpfwJoi2Q
bFNfiCBd0tsG/O0pwUXPdpXXtGa+XUd5xZIBtS+gYX230fr8uPF5LjTCbuKRcE8Osh/k4WM8YutF
QRFhBvRkPeHA2S7s6fXZb0EkJQTBLK5KCAm2DrohYlxfP6z1DFNpxSzPBLxZutfld4N7IP980Etw
oPBF+uNVkFFmxh3rGVTrhkt1kD8NjenoiJcJ1EdPRMilAEMLQw3X8EB6aTd5hfjqgGaQJ4uaTMS5
T2BQQeJ1A0ty1M4USpimzFgPyS8cx88SVcaiqcV+aN5nPUZzvx2BpE9P+9aIAjmViGrKjO6jz1Dz
8cYXb+5MSyw4RS+180UEKfACvVlRr9bCgrB2T7Euxoy62kzjI+m9SyAbGsxTtUfIBFnefBPpGtzW
02RpF/zckwY8IqQrmccOVEUv4OWbTeoHkmb0ieXHIIvS0chcgTonl8kyAX9c1+ZsfLB8fMwl3S4N
0o4OsggaLOClkeGr9BzkddATxVkeNf9b6u/D7J5ozd7J6dsnioxk3dEX2k96KEleLoY19+ZUQEOr
kuloL+3nJ5Yyl0gQEt9bGwicuoJGXvTQK7wyOctPbm2kaAujVGHMfERKi7tXhHso8A57Csl0842D
lI59xjUZWEYEGFHcS0JRWD+/aabjWXLt9niSg8W3YWw2eVpxKF+Cp4GLfY69T/GHvfZFl+uoyz7Y
5nEOwQdEe37p5jcRdon6AxUTSE2L3z+PFp5xwiQD6CmJ6jsRIhn1OXFuwudmFLEeVOD/vIdi+uf4
Wb74530GPGac4SXy8MtG1iQPlcr6YIk9ie2PNzo69du0Cs+L++xVu2i1+haQStI5MRzkNK+lXIge
7xHhBNemqoazeA/023jGRgUow1wTHxcLk3BZoeUN1SD78r33ZbXS9pvQiT03ErsvgO0GwaCP90YH
mqb6JtCxmCeI2mcbpBP9kIc6Ade2iaB1hAM7gDGYbkS3JkA01Fn6aJMzAhXhYb3+xcrfFfFVsRPN
CrM9F219Cia9yqSRMw6JI9Fyy7ThRd8n8OdJq0pkLvLQ8mdK4Ja5fJdlgtgRzx3nJqBZsAEKAvqu
br7+HH2MF/4itqifgyDpr0yMR+e7HelNy6KFCXfkJg0TNV8acn+JFvH9OAVTXPGsTk+JA2cLBMxb
Mjxxm6qD4YKZC5aGvBNmCyoqOWtC5VN6efgn1SESoQsUO/QfhRPEiCdTh/YHyeak4y+jPDkwURLI
vhhaZymoDFK0gCZTSSN1B+Vy6V0t3zbv5m55mbovQQhmNF6I9r88iOtOTkOkeQ269Rv5GShNkfAN
TKEqLqCiJW/CaNvZ6Xf/CV4L/wyBhuSGZdWy19LMWBGeIEBJtcVoSExGBLy2+9vWw77xo3/OJvxx
Y3tU8N/+ccBTMz1iy2JfDvq0njKE774Xu4l4M7xogRUz8kB1sb8/bUF3c7a9KrGG6ZGMyH7Xi/Sq
Jzzc2SOIL7mHl/pLEF7inXcnF3nURa4kvCYaGC2cG6CawL4P0gacKlhEY1GAIWOPFJ9LeIZnzEtZ
KjFVMl0Owtt+ZSoqRWKkjyNDk5X5sB6YCCCZHJNUATh7j8RiVUtE/wWjQ9kFB2SoxC8qYS0wT2sE
uLjT2OlZwjg/bamqUxvJq0ZqGUrCvrpDxptFoQp8R8DA3fJee9H2NArDIlJHv6wURE7NJpMq42iB
2IgrtZOhJ+n27ET5tV4sOyXfnODURWCrvrzY7Cg3BxUBDmDHOBgpqt967YfX4QMDGDMPyvRdEFGr
8ikXxUj9014emElQ4r3cec34x+EXd750QqY29D8+RhQkt0x2JiB668UE/zEURvBBVH4PlcGfTlDX
zCbsq3PJj5xg5r1UCmvovOSG9aMlFlGRXUqBDpxSXnTBOO5d/WXYABouNSih1GK5O+4PyA1BEqcs
Z3u+IswfVuG/QYUfPt1JK0ys82p+lxl4qRQ2R9jhtrINkHWBrJ9vtsQ4gNfuWoo9exL1PUUQLa+C
rNzV0ZHokdnw7prLkqWWWqnBdDEEU+5oSPyq6fOX5NWzTPTwbyfhN96WUYuUmQ57UvwaSMCYvcTt
sO99Z0aHgM2LVJJNkYNPEMjw0nlIbKyC9xOj2/gA4QePMtEmyN9JL7Uu3oSC4ZHa6PW+5JAvtVYI
Vu5VC8hzleViodXMmw5gDvm0MtEZLqHarukJfqlLewewbArIAyZtE7TGMcNu83i6A0Cyyb/tlNZS
5pjVnR0rxcB0/dm3jeDSYKJxcKPF8yVDpaT5SET+tqBCMJiz/v5lc0P0CKrBn3lNEVzqEJuDb6or
XZfQDGG1eNAKjbChopnWA1qL44+oe12lNeiRq48XUlt+6OtfiNPaG5uc8JXOkDwdHclKJL2JOruL
rhb3VkjJYf2ymSEaPb+0PIX2t2bHvnLs5rCbWmhJRUpcV3JYZrM4vlCeFrwwxC6QPofQrB5SlJBn
brwJl4mWNVhdpnrRYFrag/R6rZOgNmtxesq9kRnCFFFleTNP3PMXQPeofhSN1bm/jtwdUe585Y/B
hy762xJ/m/4yCOTp76drP93WAJyEayWsxutjjE3XC+B+omi+CtDewCACCy8Cs6phxZ8SgJ4FqsdV
km5i1B1cM2U+iU6qiaHdEuh8btLDIQ0seqGBq7jRQqSu7Z9wOQjxpIDDXAVn/LkjAV0S9YtA5rQ+
gUsxUKDBWSvBQDyUAZ+ZOj6y6YlAHHZr1qlbBRD/0cUfUWS0Q0CAcaJNxmyumMSFPT17DU6YRIIv
T+nMeTQJZFkGaGoe1fQTg4xrZ4ibjlEGI9cC/P+x5dZCNrT+dHT0M8EZMSh+CCQ0cRo2gWLLG97v
gCL32iSJ6fI9byiEavWRC/YxwCkA7ELwsT0lS/dFiL3vsVbuCSBIGkOeWR9I+eF7aCwDgCVh3jMW
d5PW3q+TXFvNp5p+6lsnngE+r3JdKrPUO2XQzhe69h95mYxodWHrUPBd1WBCxmtC+YQi49PEr4fT
kLM9KGz6Pgc0/5kFR7NvpAHINkzXDWvZ8SV3oBLFFxox1JUv+fTFQHpCmmRvn80/HEBY8xmG9ZeW
YlWFwJXzUJWuGXn0Hcxm2yuVvTnbWFzRpleWBSIdxCxDb5d0Q7GipmEdrwm4U/sPP25UBi95dN9X
cUK2ipvkU0WloNdnJQk/JgjWB+dWdUelIh9QeGuMHHwEd6e0d4tJ6XHZeLOFC6nRrZ/1/d2Yb6t8
117STToXX4IEJKM4ZJdBSjEHbUYn1Qeoj2SUX1SbxwDAvtKMCiu2gqXkqs+Vg27pkJMcS+QNrThT
rG5p1ZYBj6SKzgSu3JgKKI3B7JZiqn5A/EpVAmTZsShU/aA1ygKa9kTj8Oi/tlPPfuAa17Icjejo
SAx7rrvqVzNaqI8NVvQ6j8Ib7aolQGRt9RzFEwP31DrjuBXiyz6sRQmzb4i2sH2WkJIpjso1/ciN
QYyJ+FUjYrpPsbnOuUgS22fq4/SNuf+p0Ahx91HKkfp6zU/wrbbHHb5gouujUpiBfJxA5Ex3i2B4
j2NbpBM8DyENzuUFcm3dD903zuefByn6u0+wQngAMLaczxirBgRArgpkLgb0WcjOdTnZL28+DeXW
QDXJmiD1y5YNv04GapVexzTrT8kGSCSqi2xL9MrV3vULBxpkp6EAr2cx+M+nQmBZ698ohv3f1py1
yoa3rT87+ZRnT0XCmwhQBpzSqWNuEuDOmr9ARwxUwhDgyjgmcOqX6ZkQddNVNlgwrc8QohS+9607
EtAx6V6Es5AgA9eXDNWrhDo5DCLDZBFb0U191S8Cty0vwnY2+aKK45IGRdCsnsAOFASGOfhX18hi
+KmjIF4MYvLkeNR0vH4WT61blXfVkEAuZ+qbrPjrLSjOnP1bYgMxwlUlS/uzuS2kBl1vSrswMANq
0p/Q3oSV2Z2YszCj4sT7iq3zHuPHtmGgYeQt+lA/PPojBSaCArT2sXfzLUtx7mNTfF/7mmz1I9z5
ysf0L2PEhzPmxngkocJqQP1UKLFg6X+ZBxhQJn4bD7h+RW1KBMF3IRMbPkZtChYuq/aQX56LRAIL
F98Vi8t0qKJ3eJJeCg9LmBUzEuN29uq7Ak5sagekEefccVy4CLCFHb5n/UXCBFDlxKuK89rBZje/
P7sca4luNdCkDWWkUS6H7w0W9P9yNjD9dib+0zmRaFb6tBCf3Cg96KGYyJpIBiBcctGwEnkid+g6
13Je6SBGlXV/jer0lC8g+lBUxmHMhKLlTZDp8vyvktYS9V+lV0mPeaqz+5nRZctNeNCy2bkD5xP8
mxNAIo5IAqnJO9TaprwB3RBaTB5E5LNNZoi9JgB98DKsjAhXHRLHW2OzBX5uVFq4/QUqQ2H8ho4S
4w03S2NuoleboGTasphYbeltS60+xoa1l2cDA7ti2huI5tFyRcsIdRpFLd/4ts4rZrpS8zHaG254
lTf36ZvELiuCrvf0CYXXiaotbCufrChMZVzRC3u7zwJprLLdFLfuna0mF66cHrhKm5I+WSjUIhvu
xHrYg9rByxVD0/CZyesbBeJsh996TVnCBeGxnZ9RyNIf9Eu8dzl6mx8e/HLk1/BH0vGCNqVeEM06
p+ioCHPD/5/ajR+t0PK68bOoAFS+DWbJg34K+VyJ3HGn0vTMLFRmETV3SA/r6BoiQxCGOEb+p+kM
CUIJbbRgmfy+/Mwr1rIxHC8FqGDn/XuD/OA0xRHCQ6gKaF1Gca3tDZjNR2fXJ+gbNAaAyNYW4w3J
6B/fgnDJfyHqXuWEAKuKJbGg8rYD+9PNLo9fsRJYicsyqAXIwOHgAQc4lUphcJPyCmX2fT1L7XSh
y2sPNPPhJhRoMHwH7KIfKbYD7HGNBZRYOISKFvJDnX9dpCRQj67xzqxMY15Huo3Gs7nWlwKeUH4y
kXazTxwUZbtB5AveM9TJP0yElpuh5BXbRluW7urUnQZ3nphrimeV9j/ggSzZVtaXeWd07iluxFpM
sREsxlpPFilCg0JvlQE/8H2rhfFnX9kdEPfz3/2c4b+78pEqchqMh4p0Lp5Ta+v3JqIuPHBFaYLS
ldNM2fMBeheDauIxBwYoeM79mPu5nqcX7wpSHJQQgHj5rlPhh9+JU87R6zRYY4awTspuSlJNTHY7
vJAOTwqqIzPJEz7KRYVG6rAGYx3T5FKBOFF6I9AOkkc+11iBRVrq/K5AfxCpIavu74xBV//ibBg1
2Xun8ylqghmTq9AGKBYSroJg9xOtRrnhagnQSVtKI2ndI9VTeqjVbQuFO/NRtqP1P5cLg3ja/Y86
I5xEWdT5nOQOw37v8Sh0n37tfGk/SsW+reZJw/r683c90GUa/Cgg9xgZvcw+CVfcno/TrngQxWbF
qMtUg608dLKFPIEPuwSci4KYwrwi21XiZLYPkvdWYYfZOPhgJs17i0IrQ/0SQT2TAt+zw4CwvoJR
Ur/RjmjbjMppB37Wr4zmBK6FvwGR3iqmLHk8OwNps0DfwNoGarcjdOPeLn2hatTMGxe4COyF9DdU
BjCKioZpdqT74dE2SobPqvo0jx5Mue3HkNPzWEIuckm/9ZLrMWgmPz157b7G4wdAzVPU3ctEmqYB
Dd2nswGWWFbKD09yixvILImeYxcscEdp52dogqkoesvpVP71zafqV1SVIZoHV9DwM0R5+jANjQjg
hwH9jAGCVB9IRQ2sqy2KpkHeiOPHs4mAngD4Uo0lN4vzOBPDOS31NDeQA7L5dkf7mzNSM9VbhyRU
GIgZZdc++UUS8bWICwsAy9jWpAXGxVhBTaK/xUPGTQFtPMDMQ0NRBpy1DdPz4E9dMNBl+cnMtF9X
IbuKYpHv2uTShVmb7kwILN+UFXzGPG63mOkBVurqQ79ZQSitHnoMn+ewXRPMLLEFzpEe89vfjLaE
lrdAanK1GgMCboij7CUBd2GGsfdZSDYcun9hEugIiwkatFH6fOFACq5GLI1FxqDx74Yn3asIx3D0
u0DZk5IJOD1/FO5NYqQKX9O39MvGhpdkpcEJ7FOmaQPDdQgZ2MQd7HCfKLTtX4cGSXLuQtfczBQ9
FEDrB0gmMPhR7dYu0VRJHyc9cRlc/17UBdqzmIKwszrV4RB5vGiRcahnZIHHN/4Fm6YE59BEsFms
OlwZnrRNB8etUCSsqopg9WAygQeLfhDOEUsbKYjpA+rxDPMQHVJTRJtH/w/3O02CKNuvc4UNfWJx
mI/wxsWKMKas6oy+xGvnuCZ9Pz1zYUhtuXYLYIg0s0VQU6Pqx+eRJ+jO0skYLXa/o1vGgf6kXLhJ
nu0FwkOLKidyXn5S/L/8yiZI1wK4avRqVOhz3RJEpOF8JZhZDbYIexvFuXRh+P96S+jogaIkblb8
gd22yXYx+4cYNFLFMIWOXqwgd4rSfV0SGTUViOaa9yLqhdVWNGN+SJWpS7FOlp57Y6cnaQlZSGNa
PErI0/VU010AyTDKizVDtwpqduIN0MqaJE6WhXBY7JYcF7qEx2BR3duL/LXNhxVfqdTyD14xGE6o
X7VjhddOCfNrmOYNIB3wI1/Z14GKFk7iml1ZOUt2SaxaU6PW6d1BW/OpHheb8/VnEwUa0w+qeFUs
fwMvT9uzoQgW5djHi+haRlzV5UiW7rXxmCFiM+c+dUORdCbGOt1ygjqLdapplQeOnL5QXIZIbtWo
PlForrPl5kXuhCmvk6n3WjC/7F7dxG/WysBucf2v88ugyNRfi26LDpivYk+vy1LK7LkhIakMclfm
qIB0wl4tMW/Q79QR6MyZG9kRZCfna2IVthyElebAoa6hnG6S6RJEuDDcEneIYFftxuMgIgJuvS9s
fIYfIligVfjrX4Y9kQSi1ejKpCDHbqhz2Jkyzo/4XSE+JC2Krk0O5RXdGlbEq+3Wlmu1+AMD0mhv
6bDctWS5prncrdoo5ObV78s1rFRSPwG0r31gqjlhRj8CY+plLvpceCat9Zen7zysAmAT6XJAtGzQ
PkSDSnmUQIP0K01KLtl1ebbmDkM7/wqTfkeBHV6bGhhBFpbPZTjoN01lSxe+XsSzZhkUWgh+GoYg
BgQRHgpfLXAWqvnnkZQ7BzvDA1WmET2AUvrkzTlfBoTjN8Ww0YHqUO4I9DREuao5lAXkeimqCrh7
PqMq7GhIQYzTBPCFEWSh3v5sH1GW/gshjYDK0pzi2qJWLaK3SRGVDNCF5zp9+s4Fjh+jTL12Tv/9
sTeNJNp4edZQqQZNTg/44DTknCx6uWD1eNWZSUVFazlj/n62L3YDBo3Z07hMasaR5tjMzsNhEZ2W
qBPJV4MzmfGlZRCgAyoDZY+7YEcGiM3wEMxEzJuvh+Z9rzncT/ExS0z+eT10+VViVmzTck4R/u5c
B4PehAkiwGC56Ztk5v87cClx6O+pt/gIHPSuODFWy5kHetRxeSCs70LKRkKgjrY1K6Xe0HRPOU2b
uLYot9YQ9pGtVbGDoeFdvFj6bN48HIwAWoqDp9t+OrvUUBkFzT1WPjWFwr4INOc1ODWbaYivBF3p
QKQjnym4viRLOrNxomX+XOCXc5wtR60uKNEjxDHERXwcjCjcDOK6+6rQVJv0jWqiSyTq4yAP46Kg
itdEGl45JcCwqArPjYZh7ElnbbYIlMnqJjyBi0hCM+GXNbVf3FLPIGsnLVzsrOSo64aq6Y5MH0fC
/EslhuHjh1ZYW+VwzZbGhiiHwXmkGIJ54nsPkgbjvAN4YyjmaU8empqGUwQJjT6A+QP7Kse0+jNg
ANXxbl4/ObeRj+V5RfcTe3hdHFyNdYHb7ek50bCP9mVmBlQ1v8pU2qCGTX5pYZJ1WU2JSvD3R07U
9WKVlMYPNngZjed9xzSZne6GbUNanTc4KzQh5JFri3zlOuNngNBVa37eJBT6Dxnur+eXNWSRfiMk
DdPr1u/SbxYnbfFo05bmPnuP2YA1chSX8Ze66btBVImYZ/EzFMBACZ1kFNoBkba0Vllg8zRbaHF7
ZWKmZL4GqPp7fDoadYKo/sM9PUOXYwpuCnSuZVpSk5CH1KUTsIpYN7PUB7TMihSyS5+ApuzU3Hxe
tJrvG8V+u1mI3hUfwciDsTki8mKx/PwAq9gx6eL1eYp7VGFBaDQIalz3yjhIz30bVAjlg+Lyod48
rfU89t0KmcWs2tY4f0FMk3M6GMnvm48j3yUM/aVS5Nrua502fiKoFyseKI2Dy//5rAkkI+TPD5DH
+f/klLdUTO14MaPsEodpY5nZa7B1jCZW9XvlnMIEmLRF7jQurEgNNxBGFvVIH9Nn4BPJB0BVEyAg
Al2339XrojNj/S/jBtW4lhbTi+NlUgrV1Fowo030WnAw8XypBvDMHmL1sn6vNduioLgakcuXBLRG
slWtKImgju9MjLXadgXIKKi0jcwvxbP9encPOJFZHu679veqp8pu4k+vJBJAh27VsMfpnPB1c8io
SOAbminra87pWy83HMNZeQ/0WqoBuf3fWrwNw8tAeRFxIouNPLptAy9NqsSpm8wNVM339B+hir62
MKVauX5IpXNXNAiHtRkhlU7WNB4dWsAOoF5BPl3xa0cheFB9Fu0n6n+r/n4Ge4gCIYKda970Y/F7
vLe2OcCDthuERxuAZmwrdD/V6Oc0eqvTKlt6MUwd7GROO8tuYzIHDOqVzwmU+H5r+xS2QhEY17MH
cxp02fI4iQKr0yj34nU5g4wNmybxnsFyzG4vtd6blHHxeCWtO0EH97DA24Kh6c99WYpIxoVOs+EL
Rx0MgaewIUrvuWNoGOM8JDC8Zff92FBsbohXKliO74vgIisS59ZJfma2ey7Dsbt9p8vCYjB7nLrh
4BhbG4U82BqKNJtZmiI30GypfK6oXfoLOkAQzv8xYrrCqWDB4GPsgFQgHA2cg+Q70ut+KtsB2hQ6
uo3eGG06CX453nSAiP1Ex6ZiuAR3lGOWikYmuuOfulxliqF12x67Ee8CIBm61cDHuxowAHfbKgeW
lquZMcdhZsuIc45pqhbJ4Woi+96Knf1kcS9r37644SJcR0QdpUNv/eXE7OMr5vEOnaWqh3FOTUVx
attedgBE7DydLGpgUDZcd2p5ZyjvP5DybYkFYEb7vMmW5CHw5E/6uNg430AaA8u5IeP4wj7cLXN3
wR5dVbYFbhPuZYz58+43BvrNNNBFeeoHDYH3DgWkA6aRM5STwUPlHQBTxOhEwQ7SuOO3Mmc9vd57
hmSqJ296YHzuDhqPbIUBEihwGMsNqCK+1i48fiONxTKhYDjkdVtfPDJXNy5yECJGLVVcfUD0myl3
OJc1YzSIvRI59cCQlPRbP6/d/8uDcb4Kb/TcnWmgfGft4xF9dI//VwPG0BGrJUjOxzfeHODkOsY0
uT5TCJ5KvvTF9zkVKlD72bGjlop5CqIx31R1P4Ba0Gk+U5kHGeQL1bYkA+7dBSCC1BOspb4zXtEw
9TeLCDOpy2NeWCpebcbvV0i9Iz8kntXRX0ZkqXRD4X7dlXXG9aUVvfzpNesJN9ThYgh8LE3EJM8X
857hWHPNj7C5xn4Jf0zD7Z1AWF94jHCXXbehpz/pr9P8qcK8tuzrqjT/2zGTQEDj5HFZpOmfJ36a
tzSYcP/VA3l1mXPAUjXe1UU5PTqU99tApkAQoxMWgsbdL1IQNvXbCdinoaU1Q3xcYzJv3gN2fRCw
WNFvNGsm+5sWb0hsDi4RhQHWtCYjArPWwUlzcO+xzzFG74Z5zq2sP9MAUfjyOr4tO82xwpaZ6iuv
jfofUyiu8PkoT4zYFMBkFF/y39I1LYbSG7ddwuTjzMSWmDDz62Zvk6DwSS3/BJ/w19G/E1zmw/va
rSgbcH0BDAZRHN2yIoaGbX+sGig5DBcrUp2sy1YUgsbKUIiL1sYynBBQm3Gi4R4RWNJNeRc4V2K5
yE5TD3beEzbwSPNJ0C5s0slQkV9uLQrX0cmW9/BNQ3qZ1xJL22JY9PxanrWdNEGhpQkYzCOjVW/R
e+JqLa3B+Yd1rBbYMYSbTlVc25Y03bagViq8iJLHf8ztahIHEdT9tHrCkfnzKIbOpzWNNRCraxv8
oNKB2Q8nmAPZ27js3BidsqpLx4bbu3+szBKWsUVziGEjdEEKgrJ7HjBaRQQBrmd4scJKAJc47D3P
WsOXuYXg5nNaLxBQ7QZtmLLYVjOJhKctuQy9AH7ZhEr6XDiNVHDETH6pMk/LUEet6rkgui1gsC54
ogrs78N2vRpifzMKl9ddjvRUAdHFg6BgH5aE9AtwX5sY9geUw/3FSr7cbP7HKaRDfrcEqeuLlVQy
K+dCBYnt1jOnwiLCQI4BM3ka86YfPHZI1Z0Yf/NL6Pv9s3bJYcdDDf6ushlpHO/cT6QeQec5iOf8
UWY+qm7Ru1uubQGK9tWzq1G0xvDKyqtDcUcN/93qTdys3Fka7TDtDGjuTmoEsbukczOLGsg+xD1W
D0MH2PvRUULBVl74S6YTifRuYRrXXtpCx/WKEcN8rv1aiL1K88g+IIJeXBviIddSDM7kdndca9Xo
mAbR0IbXA4bnKUkfmQN/vo+swKBJmrPIyPOx2g58PufDccJHhHrHeGy9iu+s3lTDERMDchUa1+ba
VBA39iPunQ2Jc/0aqpZq08IvC6pBaERfYxYkX8M4ELWWC7sHA2E4Ly07PO3PNuFO38WdlayXeBdK
yQjgxXlKcf/6PvSK8JZKvOcINO6quRbgK3t0RWhSnGSEDrrBfdZ8EiF6VTOW5q2szhO/gA/XwkWx
0jnEb7TJPH9ZZrvlKYpP2f+ughq9W4F/CUOZAegyZZv/6Jl4AkEaY645E41vZ3K/KrbSq/7tImgQ
hibdEfyKEuNsM0v69tjN+afko2/53pqS2DhlGuEyIFR/hUxEVadw/M/YD83xrg5tZxdxFjaVBvzl
D1Gxo142Yr7y4SR1XSh7KZIomnYudrXoU13dMhLH2C7WwIl2xEM3L6brrFO7TWnJiSN1+RTH9t02
OHHOgpI/k7QYr+WiCoaXpO2O9RUzmSCErszAwlXO9R/QyrWpejLTMahQKLsSsW3+jHvp5IM5IoPo
siNU32htxis8IuFOgYB1cVhmww3Ra5UsCzqURxH2YrVwDJIOXq1dIKWpr6qJBmH6d+uRcVOWg6Eq
z2B2hmni9U93B7NTMLijulEZgRONQnHGs0y3n8GN1y8yDHAgxoMCff9DvFp4JUhJ02yOOmdOvpGU
nITrijKv4K7Ew2rVWTUmKYTxbBCd5NIcxpUB7UDs1WMyxDe0uSLYk5NcrIeQQqXBJpjQlQHfd2WM
CUqJ3uiVvXhdUyk7ttCIty3ak0UyBGsconzACHjUuZb2gz3yM6ZsJEkbPKksq/pLMrgSku6sTph2
0M+KxUKUBGcQBPsMzVfSsdQyvSKFb5gIMJpFewDokYMDB6fFwnV7QLS5xPjrQALQ/aUpS05dlglr
qnCLqohs3hshzVm+ysw6SVy/kZgkQbjhDB2CVNmhrG28LNf+0vVouo4DZjB1SLPuQwYyE2hcV166
eJozyWPUQKEOQYninftsuiMNWltz+Cw6JbuhdHunMwoP5JUgCsxVpeB/W82yKnwxR0Kwu91HS4rg
eKeRLAGroLahosqmnPb6lXK1n/kK2fgsdxrQymLEA8eopbogdO1ZdFNn/wbkLiDY0nZVmcOSay80
hxBpgTP++vQ8fvIzDPD3/sFKRQKjrXs4OuKyD2WFM8FHGt4gqW5L69HTJpasfNbOPk9OckPMgNca
4YADAh44lLK8HxiV94zqdxhsRbcFGnlgEEOANFIHuynT6txxDibS80W1VFb7CaG+QUd5bDxc4Q48
fW3M0agugtMQWEkD5A7KmgHxt9I53bm7k5AUtHzA5A/hoBPvZ60h1xGLSXYixjh9YGaG+Srip9cH
8rYc9UUoh+VjQHCtWnO+SKOasl3/so8fqoRSKgBWfTZOnTOQmDbPBwvjcaXGFzDEcpvynUNa+D7N
zFJpN3h+0xkHZl7jU+D+x+vaiG/8zUUWLb8JTwY3SeHTZhnmjuYOBTxFP1bYEvwI0dtS11EJiNEu
luDVM0vWStlbEj/q4k2jSUJkJTI7nl1ScZH8ObSUu/xoh9oS9KQZESQerMHCtE1FKElpft73FJl+
H+FeEWsz8vtPZfyrmf5u4BbkDVI1uKomfNgGCLXXvovkEtRQWvkcO/xE81DofyIgpM0l5LEc91Se
illyK3hLYT0tPapn7+vrPjCVbAjp6rOHrCZbBdyzyEnsIr3hUwAnhmxPEpNogUA66J1rvpt9Jlb3
XD3rrruRO1pue627NfrgEwYHp6PGdgqoBJ1PZTI46Lxon9kvVZ0/oTGryN8PMzbEIPI7cEYdkeV9
R+3Q5LkpIsKhHCsJtzihKONZi3fMNRzO8eO1YTDVksMM9Abk1EMLkHcMmZq8iVNQ69p/SCCG5wFj
r1R4Qc/MdkR/yisPp1QA3+VB86zJJelShHi6IkP9OGE4j835W7ZGenZHVu1gjW4MA1XbQENCbqke
+DAMv63anDqJaOST3gl7ap3pXuUTSoY23Dmx6UJEf04uhRYfVRHRY8t9nTzAGu55RZzF2pJ/Fsq9
mvA2Oo6r5+nRjKXFndgp1/DSXwSxDN6Etia3Oi8aqgwx3lQMcOFedfwPfnetlMRbLrirQe1uJsAE
NKQuGlYhBno8eOg5eHCQq/yBMd2av0YEtlu9c6DQX7m8GnobWt6ZLfinxU9QWwfkwtD/UrGFMcfv
X4xDEqszB/KqCWUh2phg37J5TUzgnuSWHideeaeGELgJeThsrshfUJ7UzqWwUOyolZukJGjZYs36
CO6D1zKFw1xi+PNaND7Ai0DMK/HndNzeAXr+bpAH288nE22gTJSgWEoYoCSLQNUwpQNFq/uH8gqd
rOaR20ZvUyhpTeFqdVyTrt9s75w2PYC7EOIiL2t9slxKAbExVOmooGysPlXKzPT9nAbzM0A+68x/
omcNyNwwqkjP0hTiKiLwwxQuCb2zJNs592c09dtbskQXGIhFm4OJ6rUrpz0nOcmy7LwOO1eTPENh
b+H6L+8Fa2+UHsOQrowJo2PcNKMj9g7963jgK4oeHPFyEI42tseUcLayA4slYxu9nWr0jRFmwNjR
zq2C3uLBQ1Skti5/bdWzUvZ38B/aDY64za2ZMXOn24qFTXMP8UJhVC+xG5f41/+Z5xwWHeZZESz0
BbD7zKTvWmvihJeL4OogOQsudZyTAV1fiudmwu2/DmF4c9tUxDQVqQP3tqZjl+SqH6Hy8n5sykrk
GCKavOyQYeeEU3foaMY1/q82wbHWtu4TgZuq6g5Pe4CZaWcs6L9ILNHfBjqW3zo80qIQ3Qtt8jxz
/Jrc+w1g8ZvLUNzXSQq1yk5J+L1Lb5atUhBty6TMzPv3hYpE1bp0vQxpu+8/fyEmNF3K2PdoDj/I
D4N0MDUcmz09usG8SeNhd3s7J7r4IlhB/j6bEt3gK8P+7MMr+OBn93hHRV5PUs3MNW/yg+5fVxif
4zKueE+KvqXqfcLyVOYrz5e80BCm3rZg+WAz9WrWXfk+xJnvgRauncnG6Ifng+n3zX+xpWlkzM2u
Z//Of9PUWU9QPVDHdS96u3HF6xnJpAbNGEJp8T7G4u+qQkBzU+YP9lBZSY0/RaVP9Hymh32zpgU/
5boLbG2/a5Ph92yN8s8cl/AifeoJMp/+Y6jUs8Qyzm1v/A/zO+U5em/ZggYLwhfH8eaY1uCiajqw
5PWuA/+ASdPxa6HzEHJPjfaRYoV5NWuR5rjka4w7A1F+0HWqHa5GZC+U0WT54FEjaM+AzZVxnBtR
tu4kPwMaAxL1WtAUn5QLzA64lq35z15pnZWBWIlHGOG7VjXtjpTS5UsvaTbX3qkeY8/ysTz7uMlH
mqBI/A8choVSkhlptgflzwDjiGeIlnaafI2/CnafKF/q35VDF8/zvRlWcU/Phpiwb7OpHzoIqByc
ZFqF9WHvt8uN1WOlWz2XTPWu8BCDBS8+WF+u5sAqd7AKWklr0RISTMTTq7idpLwlXb4bQIs28H+a
bRZ/R1lyKh9NB6x8OlpTHp9MbVz+UiFByoPtq7zqStZJ7UnDGrjkb/EZcXRY9Jb2qumThr0sX5kD
tJf2JmUKpOATNZP6ZqHI26UKNbh3wtM1ZMeOZE9NfzHaz1101PvZcG52bn1AR9+c1zayhM/YRlne
hqNjaQ4kGzF7m9axEHnqo9MgguQgk/k61BDYX+wD/+a2MBMSzqUSsAaQxoZxHMgz9afEDsSwBWaf
9y+4TQyC6NtLD/C+GAPw1J8H3drk8BxKpy5e7ckYl1MFgnT/cY52Z7SW/YdQuQ5dt/U6HHlZiwpd
fa85SGaSOZTv8VbveSZjJT2EF08lmWka2m5ezG+hMCjxBc50X1mPff8R4+12mGkeN9GA/rCGulyx
2R3iq1+xzDEfr3/P+bi54mq1CLnE2KXywXkyd1dir7ih2C+JDID5ArfRt9WXnxVN2uyR4Y5mLJgP
R2EpG2iKH2zlcf6aG7yUNoa9zQE3esGS8tO62NFJoKiuUQhMUHPjtQkhVB5d3DNcHBVaTxsQVMe1
3Vu8/GM32JXs+sYepEgyc2rCv/YiaXoDl9DweoyIxh02bYZZLyZJCXT7A2/pT4S/1oZFft6QQb6p
Ez/W2QX8GZBMG6SME49X0l3w1t3TKpZ1jra4Fe5dbPuk82ys6XUAPgvmp4pR685HPA/4H4TcFPbd
cJwupmqMrhqPX3uiPEU1XvegvfEnVBWdE8S8e0ONoIKWqiGJY/tqsGuHRjScVzPjjkHYncLML7Ac
JEPyqKtrCZfwyz4cCm3lQLDhoqb9yHjJdc/KxpmNJCBxoIgmyqkWAcmOVOckE7Teg5IFsrJcnAah
pBMg3QnYaYqL8hC120e9S+4mu5JzEJQ2P0w7vRxs5mfMPeq0syxeo+PoqM5GFKh5cQ3NnmODL6iB
+nmvwmMS6lHpEM+C82lPPBJ0Eh2/k/fabCuvayVewTTMZuIJdJBqKYROG6QXi/VBy4IEU1XNKaYl
fSa/MLzwq/ujOQJRknE6HlAqQ2KdnkvKb9pyCyqMMY59PUEqFwtiRFiZoojpx9aDgowrgiJBoqRd
2o2TPzyuqpmw3udRSiTgIQghbxT67a5s/jVyA4j63OuPQhtNhX0nJJ7V/w6BhiajwoXYZwpeMC6S
MnmsfsBKW2B+BX5TvTmqGYARcpkv4CF9+HxWjHJ58iPx9Lly4QN8IQ/fN0eZwXlUl7CenarwGUyu
VhVHSR633B9EYQz0oXGCWgABzNJ44zOtmkKyUzp8zf0DjLd76I1WBe35E0xu5bv2an30wGVMMW65
66lVBO4+qrEWR/rceIy7XidKVvXghxzagGj5uIod25MEOtC6tuONILhQOXS8bD+g8F79GnawnKhG
wNuQVasysJ3xcriXFJ4b9ZMpEhQk/dns1SQjMvnTj9sq4NPpIYY7ayLlpQf1DfvC+ZTEAJ0rXEBa
4QuiVQGvU3Qmlym5xXP9Xe0Mn+BCCATj1Dugi42cCQLfMd9We+hexMIXzNzcFSiWcjjZQevtlQBd
yMUrA7eQI2qUCLMSQRyA/S2ViaP395n22dBN96J6bgtg0IENmvlFE3T93wZxn3rnkwfr/+0LL03/
q9Bjw6g8JcI3XElkqmVPterlHxwmUS+QQA8GJZRTziRDqxMo2+2DJ4O8vH6b3d6np9JgE6GamPRr
3RMWXdD9FnS6HgEl/eNlXwjqUAceiMwHPUdjrMcMBgFHT+iLtHb9eGeSuA3z7+sqgRfuJAetzyUh
XAtOQwZ+GpgDnLxI+juuqvrdDGQ3iyDYTa+nubJd2iykM+CiXnEz8qc5HVeD4ar3ctdQiXiGWk8x
+VvwxqwGSJ4DsWMvFej0QjO2VAdE6RA7PI4jTqDiTZbHkexom7IIdRwW0jBr9Mgfs7OcJVBxyJPP
jIQRu/jZ8ZA3ZGaDDm918JB/y/Jo21oo4elJhaLyAx/rrlAom+lsDIaQnfJzmu1N5RnYX2FJPWnT
Jia9fEFDojlukGn8CfgNhchRluyW2Yn9R1RTPGvajMXYsPU32Bs0CtvvgF87S7E3NFrUPGH3mbpc
ZkEyzFRZMO7o6GE6ZNxl/JOD3R8xzWPz8jpNt0nqSMBH1qmarYA41OgCshf/PeTp/ZKToIl4OfjH
C5CkM40gj9y7+vFO/0iKe8aMlc1axwA2QkE4HrUrfLAiUFar2RG8W/IeDs0ZiRbzuxEI4xAZdFkE
HErhOldSov1xhO0pnyyriyjGntM1FQkoCcU0X0DSZZUW6Xx4dVoJ+2JJGr6aslBfzuPTT1AbGGPt
qnd9uumKy4VONWINAQclWFftj75jCFwbshA5jm911b6VQDjrKvW71WKd3d/Nxy481kjkcSOMNQ6M
m1as/QXOSDgYNSQsxIv4vlnmQk3xquOBQKGtAwI53skMgciX2eZwR2uEp5BRUf+p1Rm7ku9w3fjG
rI40u7/4BAvnGFolMs5wyL9FGiOntQo3LCCQZjLKTVCtTB+zqKQ3IzHkgyy4grFe8agqG2CD3+sM
jZxCVaODRVJjvT4JGnKoLedTHbHB9ZEfwrTkRaHMqM+fjhjubDjR4Xl/KKtofCKy9sV2/GzVK81p
MmN0cnj/iXsipO7vWH9+t52yh8PefUNha+Y0hsK9EzJofP5vI0JSmvc37pI+fRHam6zCkcBETppD
VZejDBK97ap1w4s7JRYiI/hxV0xrcGFwsTTQLKA8jEXd0r2/k5h/lLQ7gnStyuGA9kpGwge4Ew1B
K7ymjwuQFdh+qOp21CcN1ZNQOvR3Aj1sbbyPKVMb6RRv/5ZJ0XMjv0VLdIx4r0IKror2zJBkhNCN
8AaTfrPWT3cZnwjb5Cm/PJSQVNQsy3SqNHNHfO3kkZ3PJozLFcAWk/kuHvcjm8iNUo66cEKO5AJW
5eaLOiK61lwWEIOJpgCY51rC15ufQGYlz/xx9X4IuLH+HTaR19xvfObicgCGIlgom/oVIfGvedzj
oECgRC7qHNstpExHgy5sMQ5LCfx4QTKuBWh1zPS5RsfZMc4uRYIXaHWNliedLcGkLZWQDS1zXMq5
hQh3TJBxFsq3nRoFTCJdEbsalwVMTHaVdlJ32mfnzqocuGr59mBUDTEzCV1aAue5EH/0pw05jSYc
bPhCQNHmIz3JN0gZG6LA53ccc+m3uyBLz+OP7pwVsAme+dMKnMa8kFrcOs8zZxi+mL4X5vkuTWC4
n8zsFVP0YkpHqpEQ9ahg+LjIPN/GI7r1JVbBGPH38avG8coLj8JbHWPmRuPLwKdris81jpAzdGZg
Y5gr8cwZ7eoVUTayRM27iR96MFumXJal+gFrfO3iNck47TT1ivHN1ue49JNEVwXZ3HWnt3tJAz4I
Ytc9off/mr3ZC4xyx+ttL9xAxCCSHZXrGEXJzQiHRKyn9IdtX9QcIwtrdHkEHAdTElG1xCMcy9qd
TZbIIqn8O0JobBHpNisCkvoRvdEERVu2cmr6RcIpFNKbup6KC0TEwSxa2kUoYFwvM24C+hWPm60l
dX+/AJBTrz61XSVcPFN3btYOblNAAFv7y+4Ax44yixf5X3i8444FF3m19ZdsFDK2vYUZ0Gdk008c
DrMX/I0fzeeczW5Lj2uLn67lCvDhY8Zvagz47nhAtNtSRbqTljqNeeyk4GZ3lob90qk362H3mlug
ahFkvQuGmlNeJRF5/aupKiEkK6sotJElqvQzZH1EJnpHCkOX4czibwtLMxpFeEYH1hUWv/Egdtnm
cPF+adVJWNPjpLLMun0PiEvV/DX2fzuHYKC66zyr2cwZKgoBcIRb3t9YssoycTNbrzutPReWAEC/
x6TIcxk1poe4FO2TDCorCJJNF7crKR6yIWgyJEdoj6lGjP/8jvNGg+dg9mO3gZUoA9/OMBlz8SDw
rBCgifnBpOf1+MSfhIQ3+skvDE7ZNuDWG91+Lz/HpcAR5nAq12VZVjHAt7Zs5bPmF9dO3cTjSma2
i3qHwZYvKFNGZ2CtGaDATZytzpHKUMpwOleEw2wxaxwjwj1e7qLK0EccIKSG63yCCt2NTcQTh/vR
bIU4qbe+e/xZKzP4nMKiOBCYCl/Me2w03cM7QaUXIyzmrtO3usAg5j2U7gweQl4iFuEU0oc2vJEw
xegMn7xUaiRBakemeR5899iGMZNb4T6eyMD4SpQwzo9gCqg3xyvQQBx48H5fnfmYhY2WbbV8Iln6
rQ38Ec0iXkVIOC7+CO901DpQPHAj8hn1+xrOX/VOqkB0rnPNe4Pe8B49f6ft7V7DXm/RNfr3f3lN
yja+zGBPZ571vjA3NPEzoqGfFXxIuW/h0Kk71T8lFXBk3eRzmsV8c29qFtzlpfrk7emUHJWZYyQC
T2LQ7QgE+G88sQ0E+/9s+QceDUo7I6LplqToMCsgirlyxDBkCAu6uh2c3LiO7K1rh7hvZ5dLWgjz
eVpiQTVOAD+tNK10e0aG2VrdAvt+UTE/3VvCnKEgm5eOpkeJt2mZUPviKNDyvQNnrOf20z3dFj7s
YBtPE4NWjaww9+tWbyBssG5SKFt1G158ji3cEPRXjRn8Qlq1nVCmFvpw+nCd6OkSlLOcEJzlg50Z
rosxkjdatmCr4SSKpVvhTThTgROoD9zr7UFMhaq2bsCDSP8qOhMthXpyIEYL2mib4TOxJM+Ksqtw
h1qHlcgdAaDSoUH8TKA9GRkxzF7qN9edNQfeHADd3Cza3u6wcdNFb9RZ6Zhg318IP2UN8pqkT4Z0
3VEHR9eO8edr3Y1+na77mAbZNrV1i+LHDI/qNypaChnVDCAen95Ipr2I5QDYQ0vFvVJL+ib4ZMs5
hDx2ManM8X5+1OoNCxVVnGJYowv3KnjsKInZVc6tFeJ7bpfopfDbn5XYfVOhAG/Kon5fq4ThRQWi
Bv4EygYZ1VHiIsHzf9z54MDii3qxuKEZo0+93AAzgQCAqrIM6L9HzkQfdFW2woAfdU9sE6FXN7n0
mo8GkHevLvDS8CieVp5Jz8mvP7CDPKYKxKwZVYB19yu5FWHOYlm1aGCSeZcY7ILTDMtGTazG0ap8
Dh87tSDzh98JUDJlHpVmzdmfM2QKkbq4hMA8JyypzaZX9+LtSJ3j1EdPytQa5HO8n5Uu7HuEtIB3
RfX8RVYdo0a4wHxUCs8qv3dluVkqmlvTW7mIbsxZt1JB/MXGQ1iqFaZfuzsi2wuFp7PATUEHYQ+d
gHypa+J1CYh/LhNLbdb7g9CPW1V5up+fjdj22+5H35QVlqQKMcbhwrTUWsgETg5ErIu18Dstwq0K
GyDkLrSD2h16m57QOBqK+QybiXkqcGTP2SlRDojHYxVn3wGH5mRCg4xk/1ALRtSWjUZlbsaDqQuT
EJQwQG+jJZ7Q2/wkVKSvSPr7WjO+tugXIP1/95Mu5iQkJxhOe66LGMbVWcKdTULWeT5G8oWCc4p8
SplMsua7eVSWkKSK6BxCceAFcrSGAwcKdLG3u+OhQzIVE7Yun/HVp11UonKS1QLwX1qctLtvTknC
mlIOd+2FOvnXHHaKR4OhU32Iz2dGOZ7z3UCHr7snWFuvV2kQ3aSXXGjtCSWeWLnr8Zyq0ymhES7L
44na/VJQdjuFG1cOCJWaLXfLffqaqCuJw3awCHKXL8wWft5gMsAWJrRw4WZuWi3uAYVSm+4XYhWJ
NkiI+o6vOz0QercnSvfqqlE/7+6HSXTSh4nOyJ+1RifkbltaSrOZReqBysez/umXcXjsU7ejxLy8
OmFEVzMUVvtt1NqThpcppfTvrm0kBWfLxH3oH2Zoo3MXl/26e4qeWF6CEmZW2KQRVaBVc4VQqog3
JYyliiqlAnvskqlPT97ASvi2ljrB3SX51wgSJLLegUTaOaeGxhkTHBbeJ5W/o2bXcEgjbL3Yo3u7
MQDEY0cXgnAZYqu8xCsvWzf1XHDZd2of95kAbzqTgx8l65dTh/XUnQ92DwUyI+UyBD/ugO+irV9s
Sq1unte0ZcY9sNiHzmBjxdlieDvtd738YmGViiZJpmFL9FWhoJ8cKTpbkzi5ADnoRRbxnDyi+g6t
EByFbbIlseJ3bgXETduPRyNSrhyjQoQ3RpwfwaGinKpQb0bmVOFm8oTecIElqKVltyM1GNyLLBxb
RNWukRiAG43kEtgVsDCR1lTywi08Vmv4HfVzWVbWe3NGVs/h+bN/NzO6SsbTf/CFmNOqiyO6wh/R
X1k56tAomXUq3jPIPnj3SG2qQ8QDY5Q/CQCpaxzAW/xaiVFOcXR7+pOHtJAvjMiYo+Vbx/Whlg4P
Z0GtZQH2QahPU11kxHPQmePlczfAux8erDI4wdKjU3LJNGlobFH3w00wMA/dSUZifMxgzvITCGp7
xxs7OAekxSn3/iHSJvb2ciCSVKdn4/+Ykm7TN+G3EhBZQJPivcGTqcbPKkHxejktB2v+YSyeaVr+
z4/f3pn/PUkitTMx0TOOODthAB1ks7YaMgJDvPu/7DjU1koG5Qj3TlawQkjJa6xq8DUIePKN+ksm
s7l0Ciw/XOLgl66UDNbQ8wR8fQZM81jp7oLubtH0Ua5xau359StpEIBwRVONzVQpe/4BdBUvC0N3
EAy1snHgRouMZZbRHe9+0yosPwD9/wyPTt7m8BrH3qs8MuZYaZJSwGXnD1sNjVR+GQKvg5B0fqva
67VLeItLbdadgikD+jfIuQ8Fg4UMjTFz4bvwxx7Um4/2wW0Cn7qIfQhkUcj71DHIJ3dgZxF0IUVW
hW5wu2p9RO6VcGYMqIPUUarWwV/Cu4oAz+LqB+vqOr9PSchR9HktvH8pe5h57hjCw34iAzRPVyCJ
hsXYH/YE1zC5a72H36q78iLlAowuqXZ94xBj3koSufEslf4e90Fxe0fYrHTM/zb1QiYb1dW6sGAx
yrZ+0NXCB8r2grOIiGbR/dRS5jCZ9+wqp4uo+agiwNFFegB0yI+6MkvJx5SnDu2xBn/St+OQwL11
DBcdD2hMP6oUKnb2E35wfjJ6dCg/NnKhW++xXLaHiilR8yEIn374cMp0kIZWBgRwJJhvBObPeDJg
kdyLf10fVzZobPxg45+8vEgjq6FlC5Esps7PX9v5xOEP32wBaM/2l5FstFhWVx0EuGzFISuCqFC1
WNVB3V7Kr8ObjFSekT4ulSpkQZ8QhaUmnNsNM/wLmR4KkfL92jM0QxSekU6+URQrLaxImmD8ryJq
srQdRcJtgQjazlsFa4kcAJHnaL/l9dYlErWpzwCPFHRf1JeKJ/lOR77LjOJKv/Jdp2hM/xMVBOXg
coScjdmXRxvtS/DbQwP6ZhtU2ck7KIsWUJxF82y+md0zFOnzPbZG8S5g9HZPnS7rzDH6W+STBqQt
8dkJ8bOEDQzT7yyoxRb0UFz8qgSuJzjjb1jTxcGMYgx63WivTHN1yzFAqtUkJRBLOUZ6RE1eojsf
aEZzfC6hIFNYFFl805Kif6gPOai0Wq691+QjvIkU/niO7Rytf9ilwHJGJ5N3YZm/81POY8ZPRLE7
E1WaxnFvLMLDsSyWUqteu5wERMGfzx5gWI/Ul73EyqocO4DA8y1b43WN0VsBnIxEXzMLcOdN6zNL
E+RWLbkRxwxcgxagHyODVbWv7oj9KujwctB6YyQkz+mtM7Rt3dS8TyPlwa7YxxY2WWg5F5CDI9f0
jLnCRooKg1wPQhxRWUjenjj06P9v+MuWY2V7NbKv5wYOurqzH+vmdvex0Sm0W4Lmt+9e9NO8QfnP
fih9WQHRYrZyBxsK2X4/oNOECPq0GfAY0o503S9/0TBK8nXKIIKfrzUdtltVSR0i4S9DVVUqmAI5
TF22pfPy2TIzm2G5sCD6DfiiLbmOfMlqoyfx5cTzGJw43jueStyVfVCOBLNelRcyTDwJMuin7JSD
FYZiAKIt3JwIUhVwuAd+hM+lyqj/S6gmNH1tNL6+trv9bUryvkWtorLdaEsRn2nteGOBTeQ4cjQD
RHdbowfuFbN17kWDse9SiJn5bP8TA9n0nVluXPJ4GVhyTrcN5DpltyOiKRYX2JM5Aj/pgyGLa9nm
SZKFbwNRentcnLXEVtwYw70RQne/8ejDPCmqCFW4kdsd7/f8WI2tyV61YpiP+0+90sBcPA65RFLh
GXSbVuVZ84T5paJxkWVZAeJS07dCGZMVxa13VVVD3QpC4BwlMwk4Tw3xQ4Kl6LDc1ACXFtTB2NRa
HBDKe9oPIFa5U4dLCgVnfm7qzz58NmJse+F+6qWzirX5yy+E1kmYldt5X3+C7U83NjRCb2BK8uHH
uE+fCnwbIsQfAaOBd9veQsv/3CJU4eZKqYXWn/StzqZIbPV1XV+VuaY4uSgFVFJXQIeJu1pZL7CK
wTj0gcO8aHAz5sCWSaIJku7wbl+5Ti8zdKTdvbGzv7EYRXvyYgFKJgKXAX3av4ZuwBuTRq9mJdqu
eVVQyCF3Jp1dKExWADXzEIybJ+Jl7RWuycQpxMPBHCI5BT67L2d0cNAsELgLWLhMyv9I2FsjfOsq
PvHaByRtdL0NjmvmoS5pwguHNJKbV5+DnH7WQqpi3/EhVYzl1lWy9+X53ryDTxqpWEMtz+U+yTgI
oE31LPs/o19giXFOW84zLFb+vQ05IgtId1h5NjofGLpUwRkxIILKkPbIt91EN46reChFW5UuQ51c
okkpI5fqvgkEYY1EdzFNXvSEADz6sJiCkwturE5KTToYo/vqK04K8Fq4JKcFa0SDpdqYq2fvBC5n
J2Z1b0Qc/rE+GnPDJDmda/d41cJb57G28g1xld0ArATcrL279tYmcUTo4On7U6zxGfQ7owi10r9R
5sEZTmE2N1xV/MyM7iPICiRAR0Dg+G0mxTlgKdVYlMiuwA6+xm+1XuYFz1zL2FBuk/am4DRfO23o
v92LSv9nncaRCzAUlFThBD9nrsIdUhEhatWTdy/UDrz9iD8+0uowwlXKCRNrzlZJTvraautEbNu/
vKwxvz9lwUite9D8b0BQDe+Wa1lrbHN6Qu7TbwVUtJWZEopjggKn+q2RTOnztukJoytHzmrO129J
f63jVPkSd0JINYR2W2vSbbjLShFwfXU0/ZNAc1R9agTYmH6MxkGHPnGUT2Ap7LHvK9FOr9dn7nQM
bXIrt4Y0p32CJLkJ95BJ+G+TzTSNWoUjLrJT8OI5LqstVGkaX5L/0DdewxpXUpSUfWab+Nn1bmqN
3176ZC6efuvjQEpnD97kzKl+QnNP2yxUBmlL8w9Ndu+VIUmbQvp8tEMjUywakBUk1bfGDta4lM0s
DxKPPEG2TEaNPNyAjrYw5252DXNka0iSFoMlVyELIfgawC3s+coVQyAS6PE1LXP37jngB044ch7d
fcaWJRfgZKNupIF3QWQx0evHFfgP4mB/X0A4OSnHGddGAkJ6tIhc5Z20gQs3bl3nnsrc3X2qv+Ia
j+dWHyjJIMqBw8eY8nn3FegxJ1Zqmx4+CLJZ0813P6MY6fZuxurj2WAmE7+KLZUsyFv+J5enuCIT
X6jCM6PHZihswBMeduQJJrdhW2DG/yr9aQROqGt/CEc706Tc4qQkYImbHbokKsOaX7shDCcTeEx0
Xpl8TOyOvzLXMl6eLEKk0slGQFnmdfCyX/6HZRWm8KOgfTsZWyK12KQTd1MSGk2iKGRSWcnkux1n
2ddFuFk1Zceinbq/C0Ea6WaLuiPYqnWWdTfYmoQmn6DcsYhApuTevFyDixA2ebaO+2AAXAP25V37
1Czg9Xbtteap3fFJVdIt/NmESPCi3AYGmROh/BFAB89AC65b5790+Nv5rqCcINXIA3K9QMrwrUIl
9YkvbSrj41BlzoM7Q6KS+6PUtV1ZNN5m69FlKwEdxQNl5fy1+Er8ZdwASXCxi+FXZ8XXRki9CuOq
zDuellJM7EjaYN49WnpZesSVqNux2fb6mCPmfjgEEYuWRrCYVS46UBSxz8ZvG01QOzL2vadDkUrR
1/razbK+FShtTgp6PryDXDUNkwnYqnl4EhsT9cbUE3RXsYQlcNLorzNALbOvcZD4G17Eg4mjn4NJ
YptNLyhsM468wXRhLLPH8l1Bundq2Z4ehAuAaQL/LCYFiIMucYSlydlNpKD4EU9nMCLNOT32FqqC
+RAbT0OqfDwfGrhvhz4EcT/pGocNnAOK/EM+4BmZk1E4YpN6RP0gX5tz5aKQshVPZc/pIoiVn4oE
ad7VcDm5+a6aeM8soRX0/PugOh6GulXCpDQW4BecJn1PUOtrCASzuQ8wzuNjLrafToK5ZLmiiT6W
EqQqYH0/pw79Iwx73WA0DELGGvUNSVKA1xbNh23luZll+CZjOP2kiK1zwHSZ17dgqYFgUyWeYkDK
+rrY+RnBO4GAGesfaYgxCjFwJANuzFWO58gMcsGugH/TOCTBiyVLQHl69P7Aet6q9Rwu1t3/rZjX
ptb+LTAJ2227XLUhAGI4Cuo1d4oIwTJX/oywFG/B0OzD5mW06v0AjtwfmFudVScLsiMgAFzbyOdm
YpVGSWqeUntMLERy60CGZ2JRT2r65j611/qm0OqIqtru1XIQZ7XYEDDEKUESrcVv7xxZRRXPqo2o
PPx3uTsIp303zSGmfmihHnRbYLbvXjCTrjEYQkPN8g7qq1M9iIR+dcggH6BV3skTfldT5ZxCHh4k
FtCbp9OZzNdXzG18tUkiCrm5DpmfnnOmu1lQ8tbRXJM2bXi7lTQ2ZvX22GYAVpDX1/Hd7jQ00AAH
dD+faNx49FbexMOu8eeVkeK6C30tIsSaT6OC0+iy8jDgTAcyydKQs7iWe1ItL/hE+HdEyGrWmBto
nsOoipDEOOW9gXAGedsH8ntztTOWHP9ROh4l88XXpX1Itfc17LxV+86/hWsxlEv56EgOZMtybU85
6H+GIDlYE7c0N5sjZreu5jg6axadOKY5v8XetlFt8rwbWGHwynuesJqMf7M/vXqmcXLqzUpk9ZkG
y9e95a3erC+sLf157WfH8EAB/jxeeku1kT/oAP0thKaJ3WQYqzTaWfSOhFWiS4QmAvof2FoAj9Jf
Rlf5/x7UKM56mK/BkR2T0vuKi1ElSY/+cXcUdeTHZwO0Wv9kctcH7mq2TgJDfAel4DK4nIZyX5T+
u9WAEIZ4xCGd0wNEN80ICtnmjFxnO54pdoTf4k6A9G7xv62gVGt1IVrXYCYoEMgLIbN2Qk8LtuyV
N9i+wmKZBhTuXW6flbn0jWnulw8ElEswXh6k01b5sj2iPUjkzyoD08mW5V6BL2VZvDZBq3LgDcoo
iV1eHb1OmudUQZCfx9oI9qIRbCXR45/vw8K6saE4h4YJF3IbMuzZnI52mEz9w0qvDBqoak2KZ3hQ
GsRT/yEw3fY5P7D7/3ITPyXqmoPp5CLpZAwApxMBhOY/D+xm3BDGR+fYl9GqFGohz2pPqFyU+xsY
kJJq3NSWIW3J5G5b+5Ck3x+922UB9+IGQgfJ02CQUfIqvU8CXPSRg/iezAzaNesZOBwuQhxcer0+
S9dBBdLidyUG5ONQkfTLcrEBX130fU4i+dzH5iyKA5wt9rvST/YvM0xkhXDTVFy5gso9xzF7HWbS
WOZuXJRb2t0DyLj3UjDQUxggG6Bxz8JgQ+hVkgORJMgKQJh6/n1pmLHTlhm3+9KlRkXsuNpvMfPr
iOkWkHB8im72AvfZfOTjvUOe2SJg1q1GXfIW1ysEsPewPHIVJVIgU7RV/UB3MUMEpkbYYhiLlzQq
8GqQ6Bo3/ITz0eOcgYZwAIWEEh7gMb5ifiWVXOIDhBRZMI1zjR5WgwASKDjNr9Uyn8tZiZdrDK5u
/SHnQye8zPZuLhE6QSNQBH1D+EkRyaGuHRC/AyUjNGHf+AZSj8t+1eJWm/wTwwkzZO92hRRrxABf
APq3ozUy9IEoDz/r8pGrU+k10MGG91KrWUz7jk1tIQV8UAQgfxTeHNUVmCT9Bzca3H7EoGvPs/4S
601XrbnEIlB5KesjItsgpz/GNwAJPL8Qg+iMEjiIjBoxWxZIy/v7Q+E7clvG9Fl26GSj1z4ph28t
HqXOQfBhSy/evLib4hwL6W95E00dFYdkPX6TIDSswNd12+h6M1Y2Zx6JM8rS8d9b/Kvfx362ofcx
3l9a3m2uQc2apE/nSXOYdCSfetMEePuB3BEfVtgXw1VsUsR/2mrRbDDNmxUFYRQHFasNWWbgG0zO
Smo4EAQJnTz8U+XzJfbxfNKmHgF/MnZgdBR6Oo/f/5sps/W0QzhHfjCUCRex9ttL2Iw4ROYKvcgy
G4zZ1EsEIOp0MeLxjpswlqm28FN4XdQQ6RmAd0EeTvUVd7VpFtY+WglHO+41xuXLEO4La7MtbDRL
DR25fFW1PEjpOMKFocV194HXa/E2SQKy009aLz/cT2y4cmVIh85q5yxtp1pHRkR4iLi06fkFbBqs
BQcjBf/mhI0Pp/GKSlzNLzLkk+I3pOJFp0UdoG2lHVVim1CmWW3BhljjfXFFn0FRB4Z+EF6QC0PB
zncnpK+HnKLbVS8eKHGo71upLyiFJwvAXa/ea8j7WprAbBodCdrgW9W4NLBF+X0mXndnDNPZP18Q
yeCpfYlupGKME7IY2+Av0wXtwkx5fQGXR4EKCcnpeYB7P+U4Ca8J2ocKCI11wx99pL7vyavd07Y/
BVX3k9WQGhsZHcpL66Yr+IE+3if+BJcTZcStTB24Uylastq9h388Rd9ImzW7H/y6IfS6ZVP+zRXD
p+/CdAFPCTTt/zsKEXhfUmIBBXgr1/k0ktar/BSrfo2g1D3TpkfctYtrU742ZoKOqcRfn2JNAuSS
vf7zgdn9d42kippea7o+48ZOYcXXJjpDzsSbp7+XyYaANYqH64lzShW5qkwCcMfw6ItdhEF7vbdf
KeR358ZzCvmPuR2gppeHF64gWpDub09xL0AxczF/TlibJTgquPSWoN5kP2LAsPuQfU98v4RWDK9/
FuwakITFLB+vctvmnjWUJReRv0yJbp0W2FoX8si31/JNtFgi2ytdTdkqYBao5diwYEVvyraQGMqG
Q/sJ3mQ3sShMhhwl5aOIyD91waDY8cU9OAXKcoPY2frAwJLJ186NAsUVrWTaqcmh04NOsnvRtccb
PrbwSSCFQkYj/IhPQSi3wqs9rYd2+14SzNapPudqiEgtjS8OmYWwVdmgkjQ/tF7pa5TeJEWtpx/7
G8MsRhVVpWRcU5dt9y/X88TsP/c9Dy+sIk7I0M4feNyAMomIImc7FKaNKngO7sQbC1BFNqtfDmdt
OyTBSBUP4RXydUBeliPI3LwQUoYB00JJ6vE5ThL9TWmtGlOQQJpccv8QGhyc2fTicGYhS2zfPoY0
NFMbkWh9SeHquY9X1ncJ4HkuMPhxdMLhc3WqOq02trPDF3UA+HQjmWvSUSkev17uU0bPfqyfuXT0
VRsyFIz0nPNM3vSJEWSIoQuRnxZ1ojwHiQ9+eHW/60+qCPfd6uqSQKCnaGdTMMBBkWfPiPqZKO1v
jd2EPAYfsRvRpVhm1x7rMhTM7/GbInIn7DFtKCJVUds1zDt9FWfyMZ3HR+Ivwx+bOVNo1RnfDUjb
CZGLmzO4s/c8MQYm7yRKRcuK0v7ci9cYEyndrXBk8EpKhyPmOepfGMtFx1d4iYUcSEFJK4piZ6hW
xZNCKAae693ulxpmq7XsITAeiQdfpNrOkGtaItUlg+EPOIynPmSEIR8jz3T8zGV6K2+4vyMqPdrX
7iyHnZ9q/cqnupwQZ97AP56amoszpbhwhhYANZVvDHOzl+8a6BAPr+KM1ZK0maY7SXMNk+qPs543
AXmDTrozmUm15Beyw3K+QC3miJpON/LjfAdYP9y03i7frW6kFMOzNwgWwkMxzvg4ek0kaC8xjbqC
W0UE/T7XvfelgEG5OcN5vqGOfgqT42lNP4tgCo4xGBvEKf8c1LsPv5HfFrik7NA+9kP6fp6hiCih
b9CzEoRdKVhYkVuNt+vkzxCy3H8gccaHh8GIzs0zRuGWb9JnXcwooi7hmUWCiQ4RJ8RWY0qd1Q2S
Gdj9EyU4VU5scqfYd4Fzwfrg/y9zZ8LBdPP8z7hZqLNJJjFT7F87GHToFgDXbB8zhYTocrr9Hesj
NNcB+5gazW/tsUVakGV0ojCR3ZhYOMe8HKq9BoUiczOumADIOyzOxaLUGMMpdFTM6k7EQpQeZRUi
VoAAlofGEusgC9wOMNSyjvbEBpYToR0kVMP3oMewzsARptMsRM7O32d21o+jF60pFYuKGiwYlNzP
J4itgtdUHqkaw0Td76gnWtou4uEpBIr+IwUUmb0Ao1pUqjGRTCi2Yw3xkJIF/QdhXAnpKGnVxrfS
z2cJujO6rfMJ/wDhLo4HRHA66q5tdfDu0lbmwPDnRAaQql6Kvy9dcBzuqDUboQS5bp0h91Hsd2Tb
d41BRoOVlg+vPTD9tG6ytMVVDt74RhOAVZDYfjsiPy5RLc25SF8Kqu/H1BdefnO9ai+zAHjLzRfS
lQd+8+ytfBI0/HKAy49VQrQdx1pQBOga15yVUoXOmleVskd5ENzT6clbgM0WpP35JplYIW/ys68W
P1UdzVk1o/+tm4t4GAIzsoPNXxIyWLTGHA6oxUOWZ4ZDF0eh1SVAgTUL7docDXmiE1lFj8iL6Z8h
W8nBf4BBQCtj8T2i4xrjP7hC/qIa5zO+Kfsx+/CQn6j5G5l/Ibg5Zplvt8jjSZGxmN50C43q1odX
PYBn8q1rwIKNC2eg3wsPN1KB/R9FJISRUDUfzDsQzJhI0yePy6ZNvry40ECH89PTlj2b9XbHVsZA
Tx1yUil+380d8yvLD6N1Mb8TPM8wPDzpWfLSkhsEHm+IKFfyJc6ByRfcam4pevE2onUK4wc/gzXb
0xuSyUqbZ92UCdWx2CdPISYDUmPjPXcqqFbWkp2jaBUuXlbg5Xr1Eje+DAoU2HwXnAG8oQJzQ8TW
h0uNgYlojIF5uVl0BQTOEdszKZhFoUjPSqS0/qwrry0K8sZlykHUxUpGPJg/xbeZ0/ODu3sLoyM7
4zS/N4X4lrZoDM8KtpMlbEC0Bp6K646FfoReTpWqDhYig7k3LRLWGLlZPgH/iKJUouKAFDBqqM2W
9SoF9uuWiH7hP6SITyBedfx1lB3rxAVOKaIMNJuuyPXm5Rteghnb14R28JqGYBShYOZlqJ/gSoz1
4fnybLjHcwpiw2ETcUL55V5G3Seg8VqHVSPigLoRgZHRue6EQjdIUXS06/tIe1D3Ydn1JfEBQzkI
+eaDID8UmwVWTueHW4BZ6qvk3+bLrUjmF5sGJLAiQj4CyJRhLQZikEOqGKVClIIGtRh8bwiB+Lx/
TjEAwSjsjh4sfIMJR/iBnhbjAn1wqrBe1rvpGWyx3UteyxtruyS1Xe8UBckh3LAE8wXWFhG6kbsy
e5nclSdboamx43fHNmHwyD9mWslq/afFIQFI6QQMpH10UPECbZgdYnn9fqsUXBw95mjrGjRp3H6p
C778tRAPAYVaq9xn+3EkUbN2sUwluVpEw9fDLVbHXfuuflvigLDIE2Ju2gqZZUJkIxjjcFCRCrI7
utb5xP0Jvo8Pr7DQh8QFE8KVLMSm8zIdvBQVqTeqpIOqKvQS9mNc78FEb9fUWDmOeIqcxaxfrYxM
vFq6DdbV37j9O9R1lJRaDbFmjTCqfxyGz2jWFHY2fMONIKhOuC3W+3T4JjPCM1UoiplXjOYSs/Zn
CLISthuSQ35ADNk2KZDgGiy1n6+RsazQ0OJp/cAQDhyUX0p1Lo0HDqXO3BdHFrqfYgZZq8Fa2Mp2
2drDWi3TI5QCXvd5GHvAz7kbVPo8AUQpsl+qgFhpyUvuJpzTggDfy0dUE44nuPzhY442WNxtIDDC
YR0cNpcDOLMqCU63luWgwXkQNHpXeFpdidTbfrcODEWlHGVsd29Z/BJXH+TjgBVS1AZlbXD7N9wZ
yloIHStyATQI90/+QjT1gddXulabrzpATFLD0WddryH0PM2f8hyWmrP8Z3NY+c9YeMwk/twSDK+C
jhkOU8b4u1ZTMqcUUF1FSZ2pUiBeQWyPKUrXA8BmxGpJBeY+92GJN/hcqhLILoD0Ro/gk7JVTDTU
YblCFj55v1FxGDB99YJ0t9tRuc7vr473QD948AjjH/+sLJFpXc20fLuMnj0PNpW+20GLDdOvv+K6
oLfjYJIs8uI7gPMxNtnZ9LmTCukTHCJDrON2N7a0meVg84ITchHmZm2NIeahRbNMruHw6y6IhnS6
h1bBmOUxtl0Q18Y9OeH0m1WFOk/EzIdi+tB2sZBXGxH/97TvQGHKqFc/3ngMIrBaAz35ia0w/INb
yiyVYfV+z3+9Z0789ryvzG3l5I+WKe8keiF0YHABltLnUQjAJVfb0VIPU6UtoDhaRn4QuvkZaQh/
tYMdZtlDEbWpwaQR2MBNuqoDmi661O5KbxmmVYFi+f+6kKavJc311ndv3yG8qiIT5Mes8VM8x7fM
dG01hLGJbR0rBSpVI3C0NW3FoiEdW5K3SXVx3Dl1DsAsdNh3u/1P+s8KyHCneLHle3VOL38keoqk
ip+f7LTJlcIVrJ55wAHRGO3xk7YXve2NSrN4+FZ8dFaCKQx6UFcqrwGoEozYqySWPmSBrYGut6I7
lHOxNs++wSH0EtnnH6RpYcpj7F8O/hD/kZEHecuRDgflfzTlc7YnPIAaUhCEUizzbg55UoBaNX1/
MkYJ7i0//3S5jdXkFDWcf7c/RVg1EhRLl8RDL93wzmHzMR0v9T/fKR00LUrX+XNmEcUkPjt3wX1E
mbHUmQa1pb/qL3SbqGRcWsV+ICbsAmD1NzSEg1z0AU5ar4BbHuTIT6H7zjta4c0Z9dzUlCW3DE/r
5wkA6Z+gtEOWcMQFD7RMK1mtzVqzaBMu4gzeCGVC+EEseffl3cg9GwUKlhEvdGvjqIzjWf/pei7c
uMs/x9YJVm3QBB0cT3X9MLkQ1oF5fzOPaGl2a/j8/zgX2myU3KM7bwzk+HKjy3Bq0zVao4UH57lz
TE4J6slF7wCrF9/XWWtAJgbdrOXe2vsQPV+sK4hMDGhYwRghK/w8NtJGS/hfsyNs1azqWLhRAEVp
tzVbsVN6vVWYsdDKwpiayNBHP51MDiR7mPGh5hHMGcr7mL4IHeB4zdrH3Luc27CoUxad6Q31JjZM
q2BD1jZCJCuFyyriz5L7F2cEJNNlgKduJfUmHmL+xeXGGGE7y88frPmxnF9Hqj0g1sm8omPJX44y
cmKllFkN4D4Ijgzmeloa8422Kb4ZWp5GPCr01/LbzuHYs8/OP12tpfFfBvkRETI4IB03ZBMsnwDu
7/AECPxOPWDE7a/dZo0UaRrEBrjwfGWXOWcIv647cH8YhtqniYAQHxA/KGuzWMXMLWPzwGSDrDqU
ms12fjl/voygR+j/yt9xXeoI/xq1igjf+Bz9kx5updl8CAQJuUiU/Q4I3vZA3yoKvBk8uNZ9vPgS
oJ4PKV5HKEzH4OO9dJs8+gHsxDJNQHzul7zGzP/A8qWQb/+oYkqOwwDSb0RQuKftYzl6wUzio7As
Egi/kDvGRVuLWYYajNBxi1VIL4SNGwMjPuJ5Ruj/HTqdxjkh3FxkrlQGz8peT6hKYYXjibkpSPk9
PFP1mSzCYtv1nCIDjjoz89U7Ete+S6L3bI2fAo75nSFD0j7B9aheDxAh14RZmTGKTCAnbgUnm2Xz
xYIxj6IBDkOGKShxRisx0D5gCFvWpkF/LllTeKZdyTlipM2G9vxZJuLSveE2NHLG2CG3GrbgLoPV
guH3vHnP+Di82hRrnyaVAhdDfwuT42ZWgepsv/uEUOzYsJMVWRFSaEza8ZV1W6+1w1DhOdzqqZhq
aWobHxRhiRfGGX4oXCSuYcqz1nkExr5f4hba1UHiTG5f4Uez/qRHYfDdBIYXLu9PFfp5MNknWNE6
KSmv37/aSOgbQ1xKRYuxXTbCXbvLfSn/TwL9L3qosPZRaB65cY3U80PTp63pmkaqpPRqRYgejKMe
/ylmHPCl3AyZ+2Mj/wItZhuyw+qlIdQ8c25kq0jz3zQBOdDOJxYqAyDDq1PZUU6AFQqxadWgDY1B
ODr4izmUOfttkyDQxoIhxUSLyuZuTGBdKi7PPmu9DbbDh1W+V3Gy7LN+5s3FBWZwashl2YdpiG98
TOAq748Yg3P5Q4dDl++GhiL8A9Z+PmeXczVXpuujkJdatu1qWJGXS0zBPfRtGcEUDFYQBRIaKFj4
+Yar1rOem95oax/BEBujICLrA5vn+VGOgAi22SlspJFPMEZMugVHZ0lj8P/dOdMdUDdWvEHonqLS
RozoJRZIpEYsacraMN78D2/5fy8b8XVPIV8Xg2askn4cv9qUdAFj1G6vSmXdqemWh/6gSK/wHnE6
A6+lpt//+wkV58httWSwny06uqjVnmjPYfFlAyeCxkm2rbx542wgHTs6n5EDHWXrsWn0wwrifGXS
i5aIjmmckc/XqCZ+HfTXkn7TIH1LPLK9ffo/kgBwGhxtHwG3CM2WVGlslEIt7Z8EfMYZnDQUZAC1
yCRwAWneeKvtdRQNA+BNyR7RCIg4HNEO5V5joePHhsTo8HHaaTkLE3bIVb/Xb9ZAH61nBUJMvIcI
oPE9g++PuMknZKDZDcnIegqlLFsOjUgdkgJxd+yE+mx/sIG4FtbxxTyHO60Yi5iayH3poU2EzMfl
Tk/L2bNPJ+sfhTqr3KTDXddy7cMiE67iSiWMkc25P4AQUku9ktfQ8soOo6oVeVEi8J4TlvOPg7zM
K97FhR9/kN3PnigskzH0SD7RVJKTbfvyaKnWbWSzi3O2mnooyLiXMpVWgIhf/LF/r4zPIALTLdVc
IOmUeYxpUUj43uc+dhvCgjcLKQFqeXTjcsSweTlCWbSzDTGVdkFLtCiJvTqnZhHeXVkz89QZnMqb
tc1757qD+7MP11ZU7KmBDKF0Lhhy3cPkeLLAi09qBWZXPPySeuZygcahuyRG+j0wlwSXrD2NiWhR
jhi7cW9UAEzDsXB56SADVYN/t9h+B53TnLcph3mymIHEjv2FNmGUlSmtnmRTiIWeCltL6DDrZkpi
kF13DpjmW5TOuFEugZgmooUwgBNPy+0Sn1hZFJKaYUo9BccFIFaJKa8vEgZjEARiZg5wY5nQGec+
nPrCcmMV//AJk14kV76oNpvNbhdF9amVC/ii4HfCZcCwdzo5kLNiOAzNK6yuR+XA7Ulte9OVuuA2
mxPQ3RfkblnjkH1g+ciE/P6B5TsgoGrmzkUjmb5+kOE6cMocngvqQtjwolqYjBhqwnyL/uOmwCkr
qALbliOh6BHHTv9Q9T9NCTxfqmn1GM29FV33WE/2XmZWbl3tX9mq7am3WrD7JU0itpQ8VbdTf/mJ
TEIxd3z2LmHwdH4sQtiTkZZBZX3CQuQuiv4AwmcDMbmHRhZfQcZQYc7wSCQBPZtIQz/WhKBGda9+
u4kcom3xbBogysGV5Z9/3dlyRGPyCqoDT4y9QPN6+HsE73Fr53Gu+shXgdnYFy21XwD05hMyegGm
DtfhXL+rTuDvCr+HIE3nRJ1zFTK85tqCf8zlcRzs5ZT1Ni3okeOcxDS30smT9XviOr2HKDNZwvyF
RJvLg2xtUGK2/n4z2qbkRDhUK6siTDfW79QJfIjKA36ejcyw+v9rB0mjV8gd6NQfl5FGUhvWT752
Txd0n3NppTOirgGOoOlSz7WKrMraQsUhzlmgC65SdYepw1Z9OE4T2kzCVNdUGHlxxLdfkTRHRSUI
Zl3AtAvt/EocL3co+woeAsrLa/OkBZI3+MeUYSCnf4JW48LW+dLOLJ5oO9KWlf3iUzPDTYPK0Yo4
xu3RJ2wNIA12LmfhrlYHvTBDt6gBbkKUj//tcjNSAT7Jqziwkm894hXafa/BvjdgTIYvoq9ct5st
kx/5b8u7T7TwEYjZfc00MZjGGGM2kpUyd6/lSDDhaWHXYK1popVBDZK7dTAXv8s5X1LXLlk84fz3
HGir0cWXnzhx4CHs14razCdFsTbuslN7lD8fM6au72RWBwNWY3SvPc7Dn/PiH4K0Amz42y1iP5Ji
QYvz5GTurhYbPYLEKPPLbgKOe4ryY50vuTnz3VtFGU3/AeOAEcN0CqzpSJR08Q2VYFfZ2R5MLC5K
AlED9PZSjWKzvvqj+EGt9JRA1ayg0runIjSb/94qxWbENypabprjlPJAfm5Adxv++TQMSdzetCyL
PvhTGnEPnjI8Tkk94qvqMVy9et9PtK5uH6Vxtr76b6VtG+BJR8ocGUVCcBZRuSjHtR+7Gy21Rzsl
i79lfGnRi11BMPd9R6MbPgv2fqzo4gSwmnmmW1knitcQdKmbX2XIFSWXGjwHxXhXm+n1TulaBIwz
LLLKTX0O/6jhK4IX+ZUL5CfoepkZlCLGu6FIodnHkfY3x7FzAcqvVci/A0RLGUMSj8HC2NHWv+Gt
Z9UalbbE9IqhXmS3RpO+EA/ZDo2ODzQZmSgFiyqH2mcptVLZaUco8xp4MkjWY1zP6CfaINfO/hli
wjkkxsg8UFWOAAbETy3WSEIc3lA5k4Lu+l/J9SKSZ+BwlzBb6AfBM5pNAJksE5GSVnyAEI4Kr04R
EFqfZvx+uzEyfYFM6i/sEBBCDj/KoaFMc/Ud5dU3hcCAkrVmH9J+irOtCVBFrjgG2Tofxx8vJ4Bp
CoA4BBkS85uYq/bInvvNR9GzrwfRVuWwVpCFaYvvX6gfZgkEA++R1MD+uDnnyqpZXv7fXmZyNNYa
usrEqt0HE3nSFaWac8fPgCA8AUD2y+TesMBmGk28Ixs+nmeUQp4U8Aolxc48HPIgjssn5BaTXIwB
RdJRdtaTc0hCEgZbp0VpH2hOlhxlWHWZaOsspnAqFnJSxNrLPfbBgbqeZ6jAL158nUlBPR50mnrW
Z6PXBJtptXrN48fQ7R8VeSzbwJPZdt0zYf0eeu7rYdYQ070i72cJBchR3sqzx7pcNd+yPWMZJ5Ba
fKdhtDqNZjq4XObNBRZRZ/pKoVX02CJjfbWiojTtcRne/m6fHArjsc8K6GEIEO/iKskZiKeOqep0
GrPL1gasusUp14pTRKQ5fJCmqmEFVFLOpAVp35EiKDd7hvQ2WWA1O1zkifrajXeN6vXzyZIg7Qtl
eC3T+nzjn1kHTUfT/XEvRW9RG9v2K0pc5jaTmciI4L0p162L+nGHMFTuydTrZ8a+SaxGHem5MtqS
FCvK0UM/jtzHUeC18xJJ/3dKnSjKd9HwKypIRk3E1FKR6tIefdGfo/l5r6ExjwRMpnJNy0ReK8La
IkjJXIpu3IPC3XnctLytRWWiPLsg1mFRBJJRgq41dM4cOlhGE4V53avRwsbhzjs5B/5ZOerNdXNx
BMHqJQd0Adole/WIj1kW3s2f+QYpDiUmMJPse25fZB9PQjR0aMHJ07adhclayfHTtXNZ+Bxv9J5R
qvkCZaJ5pCdp19pjmfIv/Ik9sghynYmLPt5TgBs3fx+wbJ5XVJlyqZEUBrcnVG5300fmwxndaitv
zmnHJmDOkGMFDrdFUAwh0wmjWyNoxgSDIBay2naCUgFSmMavSw8BSDVtGfgerlwakNw/HwF6WPy4
iFoBs+P88XQ24jUPiBcNBIwv1daLR/gFQ+v+bP2L7F91yo6qwUWXG1laB5vT8RIsNRmHdfIGBT54
7f6uO0r+66T/klc9zgq1EqMbHMtFHUjD6UEcuF5h13+sWKD5BLF7TbXixjmehYFnm9EgaD3Yi+Z1
OG900i8i5d7ZWn5fnz+MOu7AURQvSCegpcxTaFmxq/o8+EvAjXFRfdeIAcdUGuML/b4JZtwlpxob
9TzZ+cQX5JHr9yjnbldf8Cj8Dodg8i9LSOwPIV8XYs6vH5F+mtB3at9xj+VEISNgSKz7IzI3IntE
CLnzp/igDN3gMT6SAoGi2wVSdIk72x0tkUnqMk89iPlQn+2FcoXOR2RktVNrDPS2zyZ4iK0AtPw1
qe6kZ7ty18DVbawJrADZToPtI4PLSV/15BznbNkqluxcBicI6kZ8lLnX07GqBzr9FvYSVX3ZFnml
0nIu4Ha2vnp8Zy8w1wb5BVp2fyKZ7cgTG83dEvQ6WyPui0KBdEyq9SppHN5DsjGzvjcDaSNCVmcj
gLZl63Kc1IbmKYl8IUFMitIg6+BzFW8mJU/F7c+siFwJwLvF297FiyhccEuUkS696Zw0pndhHa0R
Ya79z4sCAHP9KKM0tkxMZqnfnLW189BdfFW9lFS3WXF1L+andi5a/2wT9agtkZ/OwaxfvSkFk6cW
Qmy8zV/faB1nyd2k2LNuEAt/AoIUx3cofuraik2q98cQZuqtrJQ0Ecn2l1eSJTSJ/88OyenbmH3Y
lcqCl9OYT4P/CCoCNk2bK524nKU8uiGW86zMy2r3lkMdTYcBM3iMXn+Vv1Sat+toMEEBsbXwj8Cb
MKZqyFSXebO8g7psLkiJWAO1Eg+i3hUiBTa7qgyX9H4sym5JPtqEDn7ON8mTpZDLiwgu8V5M7K70
exh/C3cXEzF3DclmRc20FOlPZzJ9LHTJ1xNGrX/eYH1Jq7KuksykWwUnwwRTsPgY9ViW2P6jQ6oW
5pkPt5L8E2lWzLPRhyChUcZgiYNBDMOIPRfmFfzM6ettbq1emyHP7HDKkdzBKRlA4OjBTNwBq3G4
/vJNAPs3MZyb2JWY4WDXh8JMYlF+7CEym4d18B5eNLkJcqqrFHyIwZsun3Tzr5lfvTmY4PRD+sTy
NToUSIXyCeofcQylueIWOzr7nP+MiL65hJ3n29YhHW3d+A03VYsg9Wn9aHH78+pB2vmU/UPzpnoK
yWNXCOGLobjbfT7XGGrCAg+IQ5CdiIc23/bR0QcIK7r471CwvxtbECVNyHnxgKTISbeyYb/GUhOF
SSX3/6cYjHwnO8+24uDvkNkKliPaRjRCRbhlnjIUHZb4Xsz3IfbzrIQECkhuZtybmpo8rHGxsz2R
LG8az3ezwHMEh5G+HwPk5/0Rp84OGJPXycyYX7xKxAG2T9/rfxYEBEAjcddcwBifIqlFCYamG7Lx
Bz77As9aMzLFYWaVrmJK1E7uFlhvJvSfxlY4GB9BrqJrnwpvsGh4QW46YcnHLMf+U3tNPXsm2LeF
ypXRPzwKcpQsgm6ZGvKy8FIKPo1oCyJXAUOAG7NJ7HmLORDpCFPfI9/70SfayB4247D6AHzCU2ra
CPXhDk4SWQjT+lAJBeABBSRVYFHENQzzr0afA2+kn6po309WOOU7NWIWBMVguKdd21eirEKsAQd+
rWtzihHMai29W8WmptTTzKWRbdA88XXEnFiB/7jmnXZcYzTYQYDtrfcOYqtyQMRFGTKj1FkU9ewp
A8Ep/E4wzy6bDz2/jf9GVhSg7xboJlY96Ab21FOAPsadWnX44XV5U5+olZUOHynM92ShDqUusPwf
U85NWvXkNKMXcISaD/CKDUTp/jLi3sLoKgsLKNYYrq89UBl2j/JDyBcRnOBYZCrshOHa/XS82bg0
2INz4+eY9+8hJruJJVlnimq9sgdPeTpm6D57t65d1mFUCs+a4wT01LBu+b/K58IizGFUFfYhQP93
I5KtIXDNGlJFv2H3rEEHAxLvd2VjAboaGQ3kbUoz+3hBUIc4E4xW39fcF/iGVJ6BD9VxT7qOGdRg
D2kdZxvpH+hY8ozMLA7h64B81agNkw8l5ptM7OMj70xIgEbiivT5GTVmoOHyAX4fl69QRSKT8xL9
Yp0o68sdSSX5d5veEOgkPjkaU+BgyhhUlPvuH1XplF6cL+cj+BuN7dScNgqzcTs/+KiF7UTllV3v
qH9vmpSo1E+uBPY/mPoKD/CXrb0KqcdExzMUPn4a4MmbyGbGywh5NQeVdz17vBuFLfJVtRUoE6HC
7TGvMy+Y/mQpY3dmylBmyZv3yZ822h27N4Dv/Atb++EV+69vdpD+r3PAfugqma59TL5uGe9tTcg/
I/I4myxy2sZ47yi+Zbt5cOCYqe8kvgeTxsNWkJpBjr7vIeFAr6109zIOf+6YqNT/W4c7JNejTBDC
t7zIzA7TNUq+r03NFo5HdAEI2bCObJWYODChkBLEjzF1jheBo6TaordRS/FMRMpsw1jp7leljdki
Hr5WQtJvG2AR5hWIgcFbZhXno/UPUrxpA+dQqXuUFkmHkX0SR14dldEbO8rxiTIcSg2ga0vuMV/q
0Gr2+Xv/0KBj+IwCddkW7TDI+vXJGc4TYCclTYL3JPblEiFp/Nx1xKCKpE6U7YYMjDuuarv9NZuH
629w2iRNvIiAosBdpMgANPRnLirnSvHHU4J2rN/tv+drbsls/gu/b+mEXfeQciw5VUT2tA29xnko
rPn6H2KmIPgEAqV+nqHg6uXTG0br36EozZKTwm+z5LydzzWRMiabAIIiul86yNYCUQa4jqGhm333
SA4fRS0Am/Bc0mj4rT6ZvdDaZduPfH1wG3IIIHIeFFrdQ2vT8GfN9Hzkfj41pm5EgF6Tt81D5BJc
g75otlMlPstsDPKZs705brjI4adgzrKl3weOAEjLEaZBKG7pw+OCnTe4CmtmglChge39GBtl2QNH
vN+iGcqbRvQhwehe2zNaa1m7veI/bY2RBEFvPuNpzL5RhnE1U4LqLeSuLVevpaY1KNnlnUVVp55B
hS1FS3jFmyJiw0lP9NtHb6BBGK6jVZP4T65tmiR8OSg61Y49ajJaHYFIhj8C9yO26m0KAgOpIVqm
EN2BGNYfDEO3qb5+E9g3vSuHbnR+DAxp8bf/A3gCM9/zesxb3pb1sOzOM5UbZgWJl+MuEx0/htOf
mOqTkTr/cGY6Sw4+d0Beiq2Q/cN2GcQS0QKJAfD+R6CF6NdJiOWb05SNTlh96aIVhvpsSBVeFlN4
IY/KeiuoGR5L0z01tYR0AFtLz0l5cLRpR5m3wi7mSLXkLSwdwuhkZVZF4ZlLHtbjFddsbIQUTTfP
mFYjzTQFRes7zHn8HFimdQFCRXAtDGH7nV0efrwsskKoWfMwIfHtfyuIPkVEv08ItPLvS/Sm2w7I
jtf5s3yaKvyYFxt30t7ma2guldXjEWfNht6/wLoVO0Q+YMtH/wpB8oIRY4Z7GcIwmJMrf0Tq2n1A
8RyTcwCQlctO1Fn72v8wdl3AjEQnsXjwnznG2HWge9XhWJrIci8v87e7TFgVUoo8jX034ROjfo9d
xsXYioeoAxYqhim6DJ/IX4cCbC6ETdrgomO9y1BJI5AjqfVU5W+zWVQR3klQ2+Crz6ZOotAUcIg1
YlUqjibNJmmxCuk/HAR/yZBjjXLUU8xivbTAdzBl7uJvQpcrP+Ye/WOJyp9zD+j2rO+tvrH3kJjz
Qlu76wnOublXhnDiJv4RwXRl9nDiPaE1R3e6c9PokXDN7SQKqgwjCMhCFP9m2/j0SrbHqET1ujfb
ayoERVlEm7bZDS8FQn/4TZJDzpjIopVcXgwzipH3i7jPVHpX0g95miF07okddfQVMOB0oIaT0Sk7
K+NrLJQhzgtuR7RQm0xJ7jU5yj5+WJ5ZLVoHNgmLFMhuGR+RPgfzocX6MhawBSH9NXZybGxIgEhH
JiQXrwV1uQaj8B60xBWE7P8QTvxzpPFJdyyA+LtYaSdUSsQsuLEGBOwmBXHETt/oOXf5tFekvspQ
jmbegkuxVj8/9tsz8T0qhkF3Df8xUmSt6gSIVQxy5H6gNLnS/5DSfWaURkDA6Ju+hFFbjsitR2yy
KOCYuBD6Dyeb2gObpcP1np6tQjw0VH48uOI2JcdVJ9+DkqMvZzIFjV5CLrcZmeeYz7+3BGeYe3vD
4WI9LyYfXj9MaAVE77ptEwNUGIuG31A21J/cbpcJinVdzU4KHXELU0gDHx0X8A7KhAvDl3sg8FVQ
/emB6luu6dPu3O/eKYVGATrOTmaUCVDbw/qouD1iQ/KktJviPArbR4A3HNlwJjiVpor9kYdNWMFo
T9vtB3YG9nucf1Boo5qwW1fuEhuDTGLQUdws4O2oQfC8S40IGRqUbsYTwfxxX9akO95lcaJ8MqPt
vm6AB/nDbvH/8PuHdtkSbR2bGevLhqTlOwFTddouUv/Wy/U32ydsvNdj1pOKm1EAUfklFdhRp6Hp
ur1Wep8cWaKMdjLR72WgzDoa1u/GJTgwcfUDlUhoBcxmPT+OLHe00J0nK3ZOM5nVy5PpqzJPy4DK
vOlgO751WhjZnubyoBTuuFAfZr9kpnIDKT3E+2b5v9uPL0LxQtyA1Jw8rdUcXaHPh+1kZkBKacwa
rOt2ocJbWIAZBHs8pCUg9d03dyEFwuZPOKPZv9GredVBHm1J0cMBaVzNCHThMYdskBnkWnupBa+P
XE+gfUhzj8qHhvL75L/2HKDw6JlOGE+gabyXou8JCwA8ILesDKGE+MORNIb1heIefJizwtgz64Fm
RJBRFfkeam6hlmUDBMUJ5o+beNbaS2fKwVbViTsoWNbNxI8CKC/bYnKhnfi1ZoYMCS7OnJzowwuQ
WphFQzbezOx5qEvuMgUFETW/lAlIIzPiC1OrZxJcgmK1nynM9+dHZbH/V2YBdQaie8cS5tsO2KA+
a84wHLGXQ9TvhD0+kBv5QvRznVrqKITw0zBqLc9RINUqb8I77JNC8Et6UIHuTio2ePMMHRWuoNh5
iZ8Vgw3TrhdBA0ofTklYAj1iAcFWV9CqFRVl/DdBgKHO9+pvPsSHwz5eq1ZIkhBBJ3v4wK6rDsUA
/TNBPwgfpD2CMZ3dj6t5P+3trMxbhz3Y3/ygmmAm//ufu3+wgVeHkzl8+SLxjbyk7mp2Kf2DkyDM
GFyL0Z1W4ZoDM+P1aVEgT8/hnxegkBhJP2L5YkXup6m0XjxRymEXCQf/F7fFGqv9CqUBrm5Fph6N
/I9jIS+tQY8aanxz0j63wSgeQBTfoFXx/H9rSaOG/B4VZ62NVG83GVYybKfeg6v79qboM+plG6WG
S9NivA0T1D89GlkPv+FU9HjREHxug+H9uLvA434bXoID45aISdWNicFFqXCAdGg4hOlHc8uI+Dq9
ldYFyH0W60lkV5B9XfsT7soUjzwbg+ljWxAr2EYx0UAudJz4X65JtpD4DK1rl1wE4i+RZB/Kjble
SzYfEJLlqaib5qDdwF2a/+pWwd9slQdfwRY2s3+JQpRVN58wjN7/jOMmUJxujciAQ4XGYSSJ0IUO
Yxk3Bm1l4yH7ESr246XPFozEF2L43Pn5IDBt6fGzB6N+7FDIu10hmroKS6J9tadMX4T7mO7eC0jC
T7at62WXX4vwmiC4wjDjeZ09fazBN5P5O4dq4Dql70WfN/pVOv4M5MCiVe73fJY+4pRrFSsju2CQ
aDvUKQ66vEJmsF2vTZiZ45JWra+khAEQu8+N/P6irUaaFQSnVRzHDQDhMMx07MB2vC+zXHzlpu0S
Tqxwb8kyA0G0/p1MpsW6QGc5hURHZ5vYPVmXZi65K5G4hwd58j4FlristMwviMuhdvtQAQPUjUV5
6kopXICg0+ESAi55KmHsGpoSHGVkriY56yvsaZupWeeI2UHmqBCKwl07OnrAMly15sqyucRJH+Pf
U5aXM5QKdGRM7mT537OzTg6XTEvC9vK4FuWDb2ujDJZ/LvtsYjOR2dvq6RZx/hxOkB2/fs+goL0J
+G4y11ACS3hl1NlaERVeW6xX2tm27N20ice0HqL0VYY42YW3oBWH1u/dKmd0A3kECroKuGQcmOs2
XDMSHZXpu6fGv2DqA7OUNUVPKcoFPUnzQQkR+Eyv+sIl10bKyqSjm2t326g7CeBd2eY6kSNmWXDQ
d3NsXfrByRl9igTi+A1r41TUROEkA/iH8kGDDuJRVCKAQPPU5EspFkOx27ZBA2RcZ7kMzG9ASF/C
zA2e6ThKRxAD/LxilKnKGJDX76V7EzZRRWeC10GOnbI6XH/CmZsHGb+cgsiXrRVmHm0Zmu1U0c9B
m+z5cLKo6//7L+Sq6OzJ7vPYhn+OXopKfEB5r8bevhVPVhQ2nvr869VF2ZOvHVjMSM3HYvuiUd40
OUbJRq1z2/sG8l7s5sqQuLUKpQQ7FQJDRM8nhRZWzvl1PVDQprSRwgZFj7Unogu5jgp71ARqbtuB
tjD0Dzji9omV6dW4SpYRCDOEIdDSESgQKxAHC+gPa/7fsCpGCv8SLfLPgTDZeBWdmAG/meKooULS
x6SPO0b95Oipe/lM/f9Sm0Ep007sNZhl5XKsANAZvb0nMeof943N84f2gCNfYhCtw81vtXOG4IVM
7PTKFparKqkfsk0WVwpmhb+gbU/KKdpPdtrztQa80Le6R2NKeIvoiato50F/Xmp//GEHwNnNo+Qs
GflvWJvP7RblFSierVhzXUi9H96xzMuNxkSDwuasjME4JTb9cfHH62KijWz4jQrcnTvlLogsX3wA
XPC96Tu14JbH7+Q+ywXQ/skul8L/yBS/W8javccrBF9Hq0FvfwvjMKXbftuouhjCiw4x4PLwwi2V
JeWGMBfi34LdaIOD4J+eksROKmTvRNlG7lGDBr/9oJiMSSJVI1UdRjSM4YTLmx+ARrRU5T5wOVR0
P9SH3mk0pETKdkUbS5HZg26o0pp5gkUcH02D5M/ihI86ogoCTXY11Uy5SDYOR+9G2/4kLdC+BH4z
p7nTPKpmEtgHRaejzLTJrEUOaB3m9S9MMIqKAKKX193t5DqLZia4jf2WVJGSwih+SldDqMwXk0Lc
/nzSyYKlue27uH5j2ybP8ruv7PV9TiEXvNVyPCdGQ4OG3FM7lkoScqmFyBcswrO9jfKhOphlhMZM
TuaWadH4ADYWHCrM6G+u4z49N5Fwt4PunpyMq5VoM7nFVRd++8Dw0f0LhT23jnSf0ApiKLVWp87z
NcgPuCjwuZM5OQyvL4i07ZNksZW/Bs917txjecNNFRh6jo0RoLtEIknTrPLispnAFJ5obBUBBPdW
tWFAh5reSkEzAehDiWz+V+1x1MwiDzZXo82LSkY88BMYiVTHYzoqavCuMs13NbV+rgRyx9doRr2n
rxkZ1kV8nlRgALwCT1aUutoH97WHeP+FV0865vL9y6vpXs0QKL7wa/0WQPd+q/BtCqZzEzB8t09r
zkpjRQrmBWQpVaxEK1C5QDXnrzm9ItnKR2Y3uvwKXKuudjhWsIlNQCByVGAZGx6cANL0SkLTchLY
Xr3iuthv0KY6lfot86Kt5dlclk/Lg/u42wRWuT9QK7iLNv0nBR2W4gUtz0MabgglSDAy4w8CzV/q
GvgUs9hHKj0HZ3d+i7M69C0xOVUNfqkSOE1zYeYP0pQ3tLKhr9X4ZyPLyFxbYiAp9sczr4BNtsHh
ZhfijYlA2gCpcTxoPuzkKgx92qzZxGuyAyVPF1AAVHkY2QuGRR/LdGLX/iHoEwClhyNmctXDAySK
txVXx6Lzv/rJWvakTt3UaYDMKzpMXLtJIfE+f30a7OYf3E2iZ1p6FMA1V8CdtnhDIMrAsLiCBuhA
TRpvl6Athu4qmTVUT3ZrJ9megGURTPUp+lpGGzYafhljZYgmOnK1VsHW8umyrlGmIp7t25uw+tTN
Sy9DKK4ZzLUA946ggV22LuRD/kK8YCUhYTscimxrk+K+0tc/hgsyjyMT8c+6MJNMuxQWIzjbZ3z/
rY6C3y5X8fhoJbDOOexCw6La8bRpHYt3gAVRExJB3dB3EKXwWbJ0t8VO5/RLhaVo391EsodZACSQ
Tk8h5mH6ZJMG87Ol8ZluntCWGcUqJ6g+vAwgUleCSNjc6ecH6fg1HUcjqx3++YV/l9W6d/wgupHH
9ypgNAcnyNKTzE73fn343CttifOwHHdOPj5Fe5l/lQfyOR2TDBDO6wPJVInnJgtP7j8gtQoXOaag
wSZAWvZi4We1endczjS6Ib1uYILeVPXxpCZU+UWlNsc0hPu3DFT0u/eeiFjHaGMGLu9/j1HFfsqS
G3v7kjuLroO+l3ZdZR705QpSyC36iqAeh4CJyFSJl84MJzHxvDy8SWiOyu41vpzW2NeOeC7m4tuS
1+vpIIIYj+25DB4LvESj8ZXDNRff75X+v9RElitdz5nGqfl3jdY7QK+Qg6yNUy/SWZNYHxXQd49q
Qq7y0yz7Zo8o2UiRC31/n90DHyI3NN0E8BhkNJ5vP7ZH2/NhIB/5ynT2jLgbRLt0W7FMY+MMOUgn
EGLFw5ahOybxCZXJY/vAKhDBQa7h8kHcONjpgPvtaFhLbTziOl7FwXGOWsUpapd9tFB4VSej/9g/
HetHQyLVmUjHBe5rt6P4VoE4bwjQqpqMvlYu43SqRBazTsJHGZN0kY/xKI4fJuK++NjaNzm5OZbS
NjnwvhbIu+sCRzbH+wwAjerM/KuOGmfzVWv0yyTfxZBE6CoYms9xocRDC766w5gxt0KTOt5nxjA8
78TwJUo/eedNYhg/bTjmpt0wRAJae3cojWkzd8mhnSBJWT1fmO8r7TsmMq/dSAqYv21PevowthmW
Wxc6Xput0+N0/xGZ6oN2IfiKE82RWOb3QONnvFpGVhSkmfSNhFcDDG1PbyaZHfQNuUMELFPfGTPG
CFGf/41wG1dnLndyvDOTWSm6CguogJo/BsINRBNu4oVfP+VuXg8Ud4lcz3Q7ZwJDXd8rbqE21C4l
cesKGEyDkmDpZNlMCcrNAgM55FptH8A4inFf/pvtDbLJMEqzWEskLYKGvRvE7a2Efx2eAJVYZBZD
FCO8sf2zIwA7jjxrxfGA+Wo9e02GL0ZGo4zdKaLJDk782q4m7RR9CXshZGkRKXU/9CwU025LB9AW
eQ4KQlNta2P28PrgvxBskKtBxabtsyJvxoMOZuBClPqL8hu4h+MnsSefEMCssy/6QkKiqF4nzFYO
2QqLOgTuEkaNRPNcVEl0XZ9GQp79cGkircl3EJHa5AMPLE/dUVPX8eS0Fx7K0NNQ8ShwbitP+7oh
He5sg4ogfY5i2uRnz+xjCv+24MpRI8PB5F53kL4MVb1xsXyY2wSYhOn4POaZaM42vMEz1zN9h3Pl
GrEhRjDIcC3OdTTzdCtuV09529ufC8Gr5rXjBm+IoQgJDVf3FLRgeGKwq8z5ZhBM+QHmVE40h//M
3+shEqOBr5Nslj57tmINmJmxZChJZr3jlgEYf8aN+vbCLR43q7UIbpoGeRn3xd5BpdizUMvpMQV0
6oP3M7Jc7OoWsV3bjLBoWQLNEeTYLQn9JDYihnfUzUQmeC979x7OU743nZHLEbs+JoiGvH8Y6wUK
3BvzfwKvz7qR3kFLKP2ye5EXT2axFH3Ouopft8B7MITCKBSvJsNaF51njdXjltuOGxkfWJJ10MbP
x0gYHYfxXEnu/8NowKalT+o7g4dCR3MbTjuUi6gF5qw/2WaXpYOl01UY4353chSxkBSG/QUCpPam
XvonUplye3CSZn2v0tXUd+Ue556Z4Cl9fa2VeeC7IQz7n8qoaNWe+5n5Zs/tzzzIB3jNOsInfLaK
yHnYiX9exNsU6FII1EJ4bJRVm9FmPB7PghWpBpWX7twaHhBjXJLqKTv5Qc1bsJV/bFZc6kNf9Fa7
PzOpz3dOfPq1ClnBDCQGnu8rpyvyxMcn5t9PQ43uaPKlzyCz2hhutZ/EDhWYYPzCjKFSxctsckye
M6f9EtG5s3rrTW+DbWJI9B71zrNlKTOT2HRu+L9ASIyCRIwXsg453lB7Uh2vbxIAz46WPIuiFlFz
iA+9xtltxBWmxIX5obaTKzyBX1V5I+Z3AOqeFfgieuqROGl5l0aVfM6Vlex1JdeEdJ9RPEqcHIa7
muOT8ZJhfgzdKVwCAJhurXHEece9s/l1bsZKSBD9eVyrE9dv+X4JcxQCBbezy+teFciU5n/FEDfM
xH0cicLMWHAKLjH6aDoFfVZbPMYE95Dro2sZQVprFsEdiIyJoobxF3HfbaKdR/fqtii8N2NpEj92
ymEh40v9O+QJZHyVLcTcP94CKP/p9iO2iudqguBOtivJjqvb76ZNSAF2qrC8CSMKiwxCt9s1G7x+
+LetgJLL+ppyNEOZPf0I/KGx78xSYwKb5RCIDbrAnSzu53ARsnA/cd3VBSuSbjRXogSrHzg4ViAV
rfH5SOyNmtoVftC2g+V9pBRr0RAqGV7NWet+Kd4vTgg6gHNFwOh3KqtTiU47WKjWX7AovXfbUCCa
i0wgZ9UFTiArzzZtQGfxS9GQ4E3oLjcPD6hif3FS3prb90rXl/K1NR8S9HaHaDQPvJGcDmvZLUt9
yPvXmSqanBtSRt5yAt2wMhTkY7F3uydsUSB9WnBFYDDd+URYkrNaWcInW8ZdGa705Y9WJszFyQPm
sFoE+4088V9HtYjTIMwbV7jfoMHY49Cy39iqoAbsWmbhV5OH30di5GI2528SnFxcKLTvaeiczDIX
fLgiZNuQH9s1LSdgWGS0jo6CyKAv6WeuQxW4lpPrboSSJYwQPJ8+SgXR7Vd9iLxlPVY8jiUQop+Z
BsCOls7DBv7evSZs5erlY65Tm9XzjbmZOTcISNNrNnxY0bZIeLRDPPutJSiqhplpEKZRDBDNoz85
UZ+GSRvQ9UiVYFWxf2gN2pKsg0lNgmNwUSrrkZiW5RFUlCM6A4iyRC9FRyBkup1VBnPxIW/gwZ6V
r/31ebbWkAigbDs/QSFvG9w2X4TUnpHZ4WIEpTH71xL8aEi58MEeTLNVvuD6TarXo+7ldziOoLvf
e4BXv2UPrI4kn0iPdWJ3sxag+5s6HGcsq9kRVF8kVcJpsxO4cJR1gUZE+Dvi5JWKi6hpkj9VSl23
ZZWgjr4x1COF8ina1Le2N4UFJjxGayjFTAiqRuubgiDoLoP23/T9kheu1rddZLyoX9csvi+8hBmM
9XeNs6vTG2W9TlnyMj2QYnpbq8UB9w/F2BXzMqCc23UBmGMdBj4fLHozBFSWFRA7Ilda2svYXnFW
ByTeVdhGS6mpkSAWoDMvfPg0H14cQhJgr30TEl617v5nw19FjeStbWJXOEFuZokNJ/hFAOsDqyEr
V3wyOCV3S9ZhgYhfwJgVwDO5oP9jkiP4JfRZd0YJEEsp9ZMFEru6ZSyyBps/FABSzvnTNX9V8ZOt
y2CLiBXoHgPT+Q93tA9WCuDwAnD8K9+6s5l67evdO4n43q0S1zA1gBLLIS5GvVJNvF2jTBBG58TA
9r1NuLN7r/w9meETgwdO1x8+2AYRdmhfH1UVEZ72un0BR7hVn9SGEyi9oBE4IKsYHcqmXJLZuesm
GUR7Pn98PHXFOWnlm/06UiDFzQUdAgKqldloYqKLyJhMnkIcefxvD/odD1FxbeSES+8O0+Q52GhJ
D2vqY6qWg8zR+ClEeoXB6aonQDJoSP1CxZMfNobJK0C6i18X2T78HvNZ1FKm2zPbExIiG+JSuMSN
NsSET7N/Hu8mRLZbi28kKpKefI0jySNQHd3sFUbgU9gKmEgODUEcHhXgLqcoiJNHjpABtRMnTcTJ
rco8Ns9AbLkDCCY4nBAQmnNz8UG+pmS7z5RCPxUnwoeSx/Ef1HNP3gxtDHw4lyXy26OjxBcP4Gig
M4byvQCHrtqD2X0Dd4FS+1IQ04JEsKfx4EpWTWFcDzfCpmmqXKkAn1KvwxeOLMrAe+mB/X8JkLk8
ct4mAiCQRxoW5W8eXtOsBnCWrPsFEzbJMXiKHbAkxgVi4EDeWKFb9hw3hlYnXDAvWdMxgfbrZ9RN
79odbLdpaydv0p2LDSzSrHxoVNJCsKHgvlNFdwAfc6T7ctfDNeDh0RW1sHD0CooMYSs5UquYt8M6
vqcf9umYkvCUVZjdoiU1WinWTJ6D98aS+kBE+Nyspwy9v2lxQLsMq2CXxgJATk7cafNIqLYHncdj
fWf9y4Souw8f8g7J9BH/a28yi52wjpsDg1xJKzLqTwftQavCq/DvdV6ks0YlCsFC4v1N+/2QHQgH
XUoOHV41jPp0SYUhvofbIeLp9bqjzQ4SankclXK43ScXjkEzbZ1vDRmrnEk4hQo1MoOYXv+8Mj9z
GWY+MOA/eHX4FUcPZ7sCmt8ZfSJ//DMCjK9uJd/Zg+KFDIophKNeDk2xfUzK8qKNIGG1ooGGsSIb
OSJVTIijnkHY5OGxKPqktx70xVMXxrFPn76CGdRtdACCbgs56voY9o/rEVYNGjlSfvRV5MXSnNRe
Ifu8IW4VoDrU/+YJDaOOlJ5hwhc6DraCLDITuGPZF+S6OcarAE+iM1ukCIrTEXtfMhZ2mKcwjbAm
hIdMGDtI6oRKc3RI6U13/EjcupD3L6bTmkVpb96Il3HQsvtPsJ3r4NL7owfTbERy0vx2v5pviKjn
mzb50Iou+Wyqey8Z8LiiqC4Q8xNhVPGhujlvsq8d8i6UzJfdmEMmqAMcbuxFhRuuZ1jZhzxhl6EG
/X0wpceNSJUHAS+fTbWShWRQiIaETlKf5UMy+bPctcxLQ3CAcGE7yN5NglnbLSxHDKlcCyxPo8la
oDH+9ErI4AvX2WHyYqNHNIrXLh95EBQf375Pi3dTwuLDu7l3AVW/M7Mx+ENZ0WJKi6LgJJ/3ymW7
BcDVeaHdFIlXjx84IXmiHw7w4Uw/sMnDx+a5JG6d0fvFFC9USb3SwqLGxPP1lVCvrCLiTuOfLmh9
ROhnK6qh6ph6+SCP896h5a6tUErA4UEgVLn564VMIjri2QpokOfbzdOL5uf+v+rnXHNaZmpTo0aW
3i/hcGd/eeINKkbXtS5Ze8XW9SFfqG0x9KU/T8FZ73lOVoCoLUzCYEs31t+9qI/HHCjO+LgqNrFn
CdMwxoxw37h87pRmlF3qRPU441pYWi4IEgbGMltwlEHrBEhgnhzDki98W5qHBvFCEoieiTr7qrNP
o0DadwcojG0gHap0D8OjoU58BccMpMPDCMPrl92IOQ3rlZIpHQ4IZFatcX5D7277hNxxG1hd6oPI
q1X/T3s0yB7OF9nQgf77HrKfdPEZFCQHlKjQAyUYcpl8dQE+gdAUs/aubdHC1FypDXw9mFILiuF/
w/B5UkpHijGzgJs2smFr30KEJNfANcrLz5OW9bXSj1u5DvmJXlIP0tms7SHh9e0oyaIIQvZL4KHl
z4NWwTSjPkmRugwr2lp1VvQI1D6MQzILz8EVdAKI0Kg73qdyGK5Fvper7B3h8J0mIKqFa8lkdjcR
MA410XOCAujNDeMV7PEzjJsBnhn4GW6TuaEYC0V0bTrDyeIWDhcX9X2KKF0KZr8oQ770mUibW/N/
WHvmpIsMPri457y3JJzyZ2t0MJnqw5VNPr/sd3OZlVKZjUdFDmeu+B0J8TL9Jlu3VTUt1+X0F8Yo
gU0fX68VnlZvLs+Z7nOvZDu3qaFTNrqL+5BA8zoI6K3L4VgWvFs2af3Hu+rkL8aaNfgWaJLNFdxo
cXeB17/vH9Q0Gy+7O7i7H5ZOcjOg6/pVWefq1CGhunXszVEyj0/IN5OrL6bqgu5Tim3RL9Hj4Z7Z
yGJDaVOTlm021aPt5q7hV1zW18NwInw2cj2l67NEfs6RPXblyQpTiXbKGSF+JDGV6ETvAi5maEKt
DG/cO2buClkI10IzBOA9/QeZdFo3HH2VTQXhd2JU/dqwOyRmnySSAJx1nGg9QUtA+X872lhQDwoP
UeveYrtNJ/c/HqmRgctGZ9ypn+/QH/47KSmt5KRLFBnADDso20kXySnSwy4a99ktIrT41WWzL5z4
JdgVZsIZO/twRIO3tZdOznHZMnoJW1jwebAsC0gwVEH0z0QdfNYKrw+QolYOpHb0iHMGFQvP2hPK
jGhG8caepfB53TTTSFRad6FuoDjcyQM112YTMReUMz1cnBrGnJZ8Mz1jFu6RzXDNXRD0EhoIrDm1
uBrZ1qt/ZiZYtqRQpHcsrQe0FMwN4+5vYazSFUUTzqFiDyW3g90KFT/CbCCZDsKLWgVqWHzKbcRQ
E4Ady4fQTkkEtBoZ/IT7iYUf3McZUh6jeZuwEsg7iT2ChbT77V8pU+NE11EOLnnzevl6GZsK8WQI
o3oCxt5XuHbJxcxIxrfanqWwWgKESX8/f1GQLadELNVNwNMfHRViijW9Y+WiUYwSg9eDBo85CXiQ
HuSYjbdHDtyI683nwMQ+YZDw+dRlMzgxiRSAUhShSVIf7/O35V3lP20DKUcXTjSbOgNKBZeE+jCz
wFYLqRJ4EjUqdYP/tDx+xDu5J3R9HTYiLkPWwOc01Txv7mL3tcBD4mh3Ib0k1XcuQdVP+MLnHP5Q
UrbYvui1gzBKBxLfjaQ5jy8xpPC0bllxz6mnbQ+w82oL4DrXUyJ1UwOsOI7T1lxDJeHs3vFlfcpl
7+ipV/flIVavZEAAA/1mQU7WJcJEyV4flyMkCpV4GN8H/a5ITvSURzdWl+ye4QlLMdfaTvlWdO2d
PfIJuktA3pk8q9WIquX6+CyEQ9FSb4Dt5biLZUSnah+s7gffgTBXhsYceLyqQ1IWk6nti+J6wCn+
6oYPokoHqytZja8RW59XK4P0scKTPhQWT/KOJ4o+3JQt1qy4Oxqsdwa29fhr14CHPy3a/Q93ynux
AaOlkibQgMzuKNZ8VjD0+hcscCFJh931kksAJn1m7+OglmkHVttyqV+EDIX47L8wW1+ZiO/lOwlu
4u7+NBTVHNXSNeh9KcBg9WTasbI6GrwnmeFhPAYH0GsQewIa9NVYYmOzem5S9yDdbMlbRzgEm6cR
/kneMI3HjZbd6SCe/cm0snFj9zf135cEbyTJhyVBb/scnyME8o6rgsjmaAtLENU4tPM5NoBgU+sA
UWy1q7jBfz++1DEGXxljSuLkeLNYnqZSim/FC9sCI7wrWsNPPqUg6/Mp1Cxd1jeT/EgGTOCGgFop
16KQTjQ3EbVq1WMj+NI5/VOelgWh8hwtp6azKppd3kd3ae5iAO05RA8oC+opzbMJBdM8Kcfzn/Oe
HnffjfYmPcEOm9+zJrf9EWT4m+aucHtap5FofvN+tcK+4ZmI7KDgqdo9jC2VX7A14zmJkTWuQKcZ
X4e7cVwd9btytwqCQZ25qZtUa+7VKSNqbFYgHIDF0tUiKntY/FuvKQmpB/fwsVLcX0eIWpp1nuwi
Yap+zfRUcBnDr8wdlAZ++veT0s83xHfXMUl/irHPmkceTiljPGmlaqQ26oxhxWj5LW9rQM3CkL0O
zMF+f9dTEnYms3tU1zl4W2FuOO8uIk6WGeokRtNRWT5cs4zrZWBkqb+uiZiZpEu4FQ+1tATCHI6E
owCmOUf7+TIq4O5cgklYWyMcs4K/0jFYJ4tFtHomWGAtJeiO0/ki7/VIkLUrGu5XcuRPH4+4F8Zv
AI9yL8vrPi7a7zLmYg+KYvLJOJNAFJhSvqialKDK10qxBmMBWUCbsCAb6yEX6dzzTHGhseIo7+Jo
rWSrkoRkKaGpYoH29LKHLPrYCLENAI67tTkVmq8kWNSRXCgLicjVSItVFf9eMswXmLYgZkYH0jls
FDpSaSaXDyt6oXfoi0uG0aGECM5VLW4n9tf7qjpP7ZHUqkR445dOAWmzP0/q30ydnNorQTADnWpC
8WZ2TyBkanHSlhnS9x0xe9qx8bpyy+oNMUYbPriyE4AU2qJjzp7bpmgBVPCTDg1G8+Lmgb8qSU4X
TCD5ZXvQ2zIufib2HXR7EoI4NbIf1Y3mq4pe9vw8Zu20Zz1OzHVqzmTDNS4/rP+De25Fzh3Nv+OZ
GCVdbffyWF9Gcab4bhBRaVm7ql64/sZhHxp89eT0MQsuuogQyelC5bQTMko9l0WRJPLD67yt8J3Y
vodvhYuCECniQq0xWf5L/ulYBycscMrULv3afoW7KFXAdrpbNiUFuU5+Mi6JGwwtnpulPGwsTRDw
ClShGvejdxogSRNibN4xtmSBo3UlpROqljqy5y92I8Um11hPJ2zvpGe7SqE2HSCSVJ8MSG5JbNUQ
7QDA+XtqCtCQwK0Qb1y7ftfE2aKEoDDEKug93bFRIBX4cvPtEa9QEkedQGB+PBojs78Cm+MJD6lG
v9F7nfg3J/mxxJPayHX8ME0BOt+HcQIFpAo1tn5KNiwiC23RD2OLf52MVuz0Z3nJsw8MASSHSE8M
DVgIjAMQ62pTmE35qoamS45VIyRvfPuy6RyNle1yw6PXtse68R7sTSXEgMdVrNtndSnzAvnT4IW/
Lr/gsAmFkTgZtc1VXus1KwU3eX17AsapEh7DFWA3WXixv0A2kBG1+XA/7mg83oyAsuxRSp6rvyBj
IsprNx6OzN35coeRlg3GSm5YAIUrkyeKREy3nVTT4HtufsorzBVg9Aw8xNIhWMVgFDOau2DyPy0T
WVccM+OiKpheeorsqwV3Oix2MUVDtJyUvx0S6OdRApaarT5KVQ4lswn97dcIRg1Vi3ATwQp3t8c1
hXBRYKU2pS2xAtWYdbq4hMvetOjZPD7u4yh/f2V4X2j88sB0jGr1r/GC5bbdqsGuKMmBgu4Cb6Ph
9aVecNDd/TbaRDfR6iRKGGwlbJ3tkKmTJSgmPtJ7zmir2R+RSpkNIE4qo89PGXtlAMuJNZuMy9Xu
EyPQffIuAo8p1AXI0nM8PvYVo9VcYG6gc2b5BSuux2t0Rzdf32VhG7vLmvJ+MJEdIWs9vbArwDab
KRoEV1nQX4w7OQQ09oqRJPVSJh6WOuZm6MfaTGTNkagh3BAA/dpmDMSDOeYI6+D7zJNtQEUTirjL
SepX3uBM/HR2/Z9dpjb98rytJ+TvQgRSY/XdspTEk5eazr53EQ+moEqbXN8RS4dkMr2byz2Zgk+u
a9erFdB/uMbpzYJWzXRLp8Exxs+94hxVt648os6ACV6IE8dWYe0+TuJS4lsBumHQf0JHmP3t/KpV
pvpthr27MWaSEuo8Hi7flUfdT/sb/X2WzH0y42kXR/GGZID9GgLsg/5vl54dG+tDBM2ngvBASZpV
O+Mc1jyp0C4Svau9Gjr9DLcZb+g2YP7mru/Y05+m9OjnIBZ06evLVo+M6SFjlkMxdo8/NDAC/ecI
gzKOUUWKzhme2q5iIPOnmflrx+WXUV8hTWhGmDJNm/7I/FBIfqQk9PN242JAMbMxRSXL9A14+m8x
ikd0Gso7SBYXKM2XTvPbAX7uxlh6WjUFvU15IxoOpjfFDdUZ0XM/FbDzlMLurlPcTdj75dYl8Nxt
xmIlFfz72PIhbMwvGfpQ4ky4B1/PlYfONbXk0C7WKB5wcxXKiPTnc+hhTvsP/e33pMYZNGDFBPMR
vk0L6y3FcqmvW1tzHy95Lax+nsUU+R6Bx6axV9cnyRu9sTfGxHlKH4k0qxchAd+HUIOrfPq4V146
AcNkNuQPVUqhtp1FbyvM4MyTZtj7MOiaFbxHaCvW/e0rwmeRLAfzLthAB1lKvyNQ/TsvS/mlEy8d
TDjEJ+YO4p8qIjGZlN3YfxO80yydJkL7jTyqdHt/xcOHlSUbj8ofRr8HZ4Wskp44qmMHY03axz32
T2ncRONUjviuiu9W5Ncf3pLS7rRmQGBk0uVNIWskl7WNqFohP5N/JbbIB0XUWP65j8dO5PI3+MJJ
+ILh78cxLx/lhbQsceih78E/H0cM39abjuG3BFyVPuXkJKAd801tYNbgiUiDV5XjaFlDkHcTnuLE
wBW8Y5jFkdvRvzyU8gK0xlZ2KS6TguezgEl4m5wZZogQHCQKFRImBhnAPAPQxF+IJ8jom+Tx9zQP
tt03/AlVcUYZv/LMRSJ7lL/UJcxNfneV/FIjIDqYTaT2lN156gV//VOVaD/Amk5rhVXpRklF+g9c
PrgPKHLCwn6iXNEJClZVrJOtu++GuPibY4wBjshXhHZukptg2104XobTt66GS2rlW/rGnpbsHB15
0nRO7j17CvTqA36XVWF085cGCH7s5Jln92YkLbfMsqpq62uBz2/3nshOgLVzNr3hSPHI9W1lPpu1
0xONv8FPhO1JJKGkSqXL5boN3VA55jcqSnBjGzQ4cJ5eYWMHnB+qyE3Z9pDWPuZ6QZoSdpPXDJ2/
I8G9x0Kvz2WXNXcGWAZ4Nm0rlZQAMx9cY2BZTG3jCGfNEl8eKgtA/Em1wjf2S1vagE/5ZRyxOXXx
ABwM9svD0f1JW4kYMYCol6NHC9xbgebpRmewpVMyU4tuVuYlq7r5dVy7vsmIgp34J5t1Ouclkw4m
n7O8O+tWxkNuLrw/lezTMqJsF33HlrviCPtvjmbM1ZOQyu6UEsBFp5YYQPxb+YcYl/TIusGCdJRn
/ah3GrMAvuvvDqGvoWuCKQge5eLCIilp76fNhjgF16UhRXpgFxxzRIrepiCqRllJfzNVyiPe/MxI
Fyjy0FHa9ov/7zIcJ5LpHJ07wfK8H1w3s95HLxvoM4/koSP02ZC0M0Tu8xt/pW9FpZwlWXKixoVv
gYwahKGjryhB2RQh0Ax62tqTNzJVaVWJK3ni2ZSoMPhCarkw8lY6HAJU/ko2RYiJaPImnR19+omJ
T41kxNIXs/3g397funKV6AAmGpNMmQv2VznaxqsVx64KzE72NIpg6tZaqEnz930R/7Ba8NXfG6W2
GkvMrUCw7bJfuH3qA1yoQEo2DfTSSA5OWT3WK3KV00JRY4PmRL+67pKr+EZ/cVryy30cx2gIJg7E
21nj65MgnK8a2c4He7qVKD89aQazr7OGnUBkLC0XOI3r3zhf29pZxWucuBsHC5DRDnu849laqsf0
gqjOLQt7of2kRjKJTwng4eTJGwyxxE73K/52PZjpGXJujL8KfT95mCNMRDhjW6BNJ6jxN/vrKiUl
VOXW3NrUtn0eN3Jd1nOxWo44nGfJto5nlpQtL06ErNH1XPfEbLM7vw3wYibOM9EADZZl5VOWnjcQ
sYmN+OqBbcCRCw3PlOEez6Gnk1FC46opbwF29+FIXpn7boFC0ItaVtLmij3Ta9YHrIp6JFFmT99t
ff7MWXSgDfMan0m5+ETpKzgGl+5YWhogq0muUcCeWOwbaazf8I5TRMccG6niFV2sRCDP6+sP4fNB
kF/fBszr7S8Y2AzXfP3ShyxinvPLCqFjcib3uv+lW7nnn+DpI3uQKsCQD+tNaEPqjfpkBe44ObST
/8MTv78EV+9VijmBQ0TY7WXUCSui0z/1xl+3swdNJwW9vv9T5bIVcX821RlRcHzyjPS7/eOUAeCs
GQGTdSUsRdBZN60W407x0Jvl7xrPBYlkfxFg7j86LL6q7xwEv9twsT5FJH3/LO+WkzhlMh7/9x9Q
KUraDr9SvKFh7Dol5xAYwYsSbGRhD9KuHNeU0PWrBLqN0/msPe9B3bI9wNky2d7yzASPG2EZLWiH
tfgOGXl7TbpwumMp514Hi5/Wzt5PXggkfFuqyTEHLWpNo4kfoM0hNdL+P+lrNis20VBCSqCZWDDT
T1/Jmg8/XMGDtxfx4/7iBmVb0oUprkH/GKRYSzAM6Qa1Xbs4Sau4D1skk9GKZu9hwXfh5u74Sjik
h+GaukUmj4PYZuBPJuy7hzoarIFuvFGJmj0SOSoie2lzGDA+NOhfG3hZRBtqkM022Y/jgjc4MAWO
t2WtYSzWmTkpQqZznpH64e0sA1obLv15+wdxX5pN8L7dq7RX9VLcT4oUpFsB8M7TZUR9SE+t3k1i
0pnnjpM2Jv83o7VhAjWzw1cLGYn+sln9IkqX8JjUHuICP4ObPuyFtksm3nHGS0tAHHq0M5aKxMzH
CrbP2FRcFFDHoUORZ5F1S21AVdgH3e41ziahKXx5ZSOzArQXYjZTQJ/+R4qd+JrsPlvDy8U4XvcX
cKFxYP/lKkX9uKhLCOhUzPcDlwqKGBEylvU+4ZqW6r0iH5DVEsZafr7zRqa8KjQrVdEX/27gctNw
dVLmqcFfp67vv/7lw94fb2lUoDY53cC02d933E9eBGC7FVqfkkOiK4FDLtzuKClVWK9ZKcVTOcY6
7jZsORzGAE5QtK+YJ1fYHHarClLDQJvd8BE/oaelAjMITaK38WXU99EhE1eX9l9Lb6w8pSUZXGwn
nqnIDv6wucVLSFrGn4UJd5sKtln7M+/1TY9XrgBjJCJQp/QptSCGobZ7u/Zt+ccoVTHGHymCNC5F
P8dBKqIszTAFKwOKzfw1vuAdHl6WoGIMsorSYcJd++BLTngQsLNtrFnOw3mdyXTsp+3FYdLxxTQu
90jX1mS6onxt/r8TKnItGWMev8/kIch/6PQ9sg+1jCgPUXd+MAC1xkWdK8YWPQou2GkLv2+PhlWG
JwWfHP7U9dDBVcSnEQIJOK0yzaaEtP0+Y55PIP20d8WIQxnrWg3HiZMNiFz+kvVprDPT9PSFXixp
SsEkXnduZ6w+fzNoa2DITKVZcFqusEY0eRB6bFT8YIzuBQ5gkeN+qJF7LEV+IfhypAslssJSi4yo
IRSwYSvXzAZn+EAKl65Ws63qTyxb1uN2fnBUafErm41Ebl3gdTlxkYi3GX7dr2nkkZYFTjazVxJr
yJW1OEudUi1E0mJ/Qc6PVtgHz96v0clEVPCYX6rs35Ie2IwqiL3DZce3s1bzGXWth9KLJASy0dDE
quAkQC6ziZZCbKApTpV7fPbhGrF8YVvx6CSrI9pJCtOXnfVm8mMAvvHcd5jw28u69e1yC8byey7S
Ig/rDu/mWSMeil6/74sO6JJ4mCznDOdDU9SerVuQpf7T7a0QWPJw9CZxFXMivnT5H8JEIpcaRkm5
Hl1xP/uw4JZSq8e3+T7rwgzWB5rM8xmgGTB6AhLbxKB3KSA1HNr4pR2Cc7WQ7bFRadyXUwQSXhqO
CUuLQF6nSnyMynH17wePRefPXCvI2HEMflbwPvWCi3vp4QYh8iOhoeAKlg8Nu2NURFYRo88foo/d
2Aq5qL+EnoScz8tMZr21Ll58Kghgn8W0DNEQw7ZfcAottX8Btb8Vmup4xIrtvZ96lc8KswIUZSqu
6IZthwWFCT6LtKJIZzYc0LFnFkpUeEPzg9Vp9Kgl7lMBo7R+4nEl3WwlxpUKknAHczAl9McgBSWR
ySF1hU5HS4yJHu8Awp+Q/uVSAU33SpyAhbKUVJsrJ5Zp3JbwWorffef/xmbRjkjh38nUf1Lq2OXh
FXixoakGDyZHS8Ss/ifBxro2FTsXBmwgdSPp7sXtggj56RtZYH0BA/HqDy9/3fgO/xqviyTglJh6
wm7GuZT7zTBuvWy1JS2GhKfTlfA6ZSSJRZShZxIVF/tM95MMNpHUSydiIpY6bWePvBF8Wg9eRvDK
XafvQHOWtsTmkYvR3E0gVcW0CBYGHAWakfM7n02SKdlSkwcO6CO1l0n8UglibnyewjMGxy7JtMg4
escT6tswNVwCVzy2+UpGmcctA2VihqhUce6LUTN39R+39t58HMOO/tReATvqqb57BH54xAaj1sfF
MXpYp5tAPT0CQQ7seWLVkfzBYbhBIb+l8EjWOed9PkWlPNJwyyEG/55IzOW724/hzIoBKceVZCvP
gLyUZ1me54v83RfePXuDb1dCcDR74IQGS8OgI4D4EFsEzKmaXyFUiu1oOXUucmtOY/GG10Yr+ofx
ys1V8x2x5ojZkQDgA0sVhzYEClIIlmRBUu8Y/20tATKkLghTVsaBAx2eAUJ4UC4/B/1Y8WaGfQ0q
dVAmqY0PnOeSAEP576s4+jKwIhGoUy/ZhoAs+R+W3t8y9+XM4KuNlxE2rd8DTQE//++Ea+tU41T5
OiCE4jeQj5ykhjBc8z+1Xy+kWD3061DKik3q+BJQ1Jnkdf64l07tai9ewUHIaBBG67A7tEkINeav
z/jwHP4+W3Rsxv8jSTFpAwPV/BHPcC3YXJBgvVU/D6gmEM5DrEeH1wxY9MldX8+SboHPxQHAIzPl
/0KAwFSwEFHVq0rCrqlJUr6wgl2F8KRfhj3/SJcimhM0pj7+aggEYormm+ACp3U0zjmQ3HXk1yVs
JON/WA/recsAxlR2pDCS5dOvJQvzLKOn1nvecfAvh+TMnafnbe8sA+cumWidJ1uka2lJm1jDOX87
qcF/37ZYuGCgRNBOEt5afIxsigHiaNM9C0BYzc2QJ+LZYhY+6uogbbipK1mH//qU7wMstB/cDiM7
56JuSTWaG50j61t9E/q5JFp8E/gyPobsjGfFK1Q26bMf0Q77XNQq8j16eqeNMuCr7/harQEM3vPm
BzEw8GuYJcGF8G2r5sB6dJ/+BlO84VZFb58AO/gYwxvGO6ewKxL5wiNvubs+IJxis5X5MhQHTV9d
G4irl8MZQBppShCUj8wyR4U7x+Y4go/k4zvilzEnsGrmVrEtXiTR5k2NK4/TF/lhkK/8h0obeFV2
FTO11Un5WE0LSgZjCbtZTRaxxZzWW9jwVDkMp7Pt4Xou5Bz+kQBC3RDBvbAvBAI/vUw6xEa5GPc6
O2XZGkOT4lDlPvGtmqIOckT61ampeO5EW7uAQnfPr/NCSgQuB8yf4CQFf7xhISLBc+lm7JhPUK3I
7tmy4gXy9FtD6rtA7LmBxO55vybwB7MKnODeCr5lcpH5xR+NCIvfm/Q2V5EPspj0BL1w82qTQze8
/rPTYTpbNIgCPzgIV3FEBbs1yL0TFNI51mA359F8afgBPVvIs+zuexe5xey/1rWmUQL4RmRTHwwP
8hoj1k7ir1YBXhNpsfybSm616NrGXG4q9yXNUrqgKOrwncc1ynGPDck90b5Bc3bVJ5t7Vx9t4UXS
s3GFHu+8JM0H+f8SEi+cLBE07pdLLfusp7s9lv/FFzPEpFnYJRxj+DTCrzJZ4pbDmcjMki9aG6VO
S1ZBWTzORpT44qgqprH9Piw6KBnbS+ToSfWQ9Br9l0gySzSPiiPraIgC8GdBvEYCE7eCUPaAY5Np
rakOkpNUx8FOctG1OYpPWU7UGLL3xOOn0y+zyLs8RB5YK0/Qs9ctf6WlgxY0ZJ92YlEyPa8daKtP
Gk85LNpQi/lFBklJ71ln6qNnAHaIjLRV4rrzF61qn7xmS3jn13X8NWaHyDEpWmVmxZIANpS78qCC
ZDhDDaKMDyfDkcJPH6SgqT8xdFf1c+eGhjMN8KPifBhM0ACwkEGFJSx/KLh0OQvxEJ7fEZM9NRpA
dBqwSJcyscktmOL91ejGoNpbFkBbCTQcadqNnhM8jT/DDrtMddD9BvfqDeCeuZ4fxeR7rjO5tNz5
RLw56Ii/BbpEkx678KU+l6jkC/NzHpu1mmxhyoGIQ5Wz+BpCjCQ7KPtsOLZYCJfFJY0Tt81WpzXN
aGuC06CLde3hiQp+O+6itneqbWyjSw5J92Ci5lWrFwvMQzZ2/l4LhrAxMXWfUyltAizfKNw5KtIU
2fwAVXuKH97AOdWLUWUlW7rGHpP5vjm3HeG5Eucl0V6dqM9AHQ1PBebJWMak72eiXWcpGH+MCu4M
JUfC5Kezk3YEwVAKFrOKOokVDjVccmTRrLL2EW7DaZZ3eq80bFAZAO5mAjpX/LdGTcG+5sH/F4Mh
Vhy66BWnXTf14wOIOLUptdRKGSODEcD++slpr8FiblbUf4nLPo5ZBsHcdnQ32vIm0gCb9djmD5Xk
L8l0sSPYQNOaC7dTqWIyS+BakpbYTI210xWpgobRS1taTUjNBqgAz2MBTFffDKW18tC5Hq1JKVA1
0m8dED7ucffYO3ya2V061KzQLZPBs9N4G3ct+mV8VMpXvGMenyGjiF/T5RhGNm9l/WzP3186Q3sk
vYDUvWFEWZMdkH+3kXkVMIWJWH+/NfoDycuWMNUIzlkPBeJsldGu2sYwNJ+m+kPO11FGh+StK3ci
jVXtMJhzxWjCEKBoCZkbH2F/t1zyTr9J/5aeY8mLV/ZrAN4vALt36sCzn9PA0qirumPeuUlORjYw
vlcxFdtVxg/HpDtXKkx9dXxwlTcgZOsDYf26E7ivqllUXbVqqHw89IJfeHDTzWj3nZG0echqFjCu
bAa8KiVG+c0xwKazSpaTTyrzJMljSAPIf+h3bq+RgEey4WWQ/5gKkzmpRRkhtXGMpNfOLZBOcWJM
zwnL7l2wh4w1MKr167jVpVVELVfLMdRhh5bse4UWFEi4ziQjtjkPvZhnjNasvstogj5G4cjXbLPG
Od2KxwWEXcKwdWhT+u7h+4AGMLdfpF4d0llRDDyN1F2b0OO60op7CUl2YMLlVis9nAGMYgF31mpC
cbxqz24rSC4p3RQfmQtBl9GwkdV5f7B6tulpD2xyogcSyfbvej1D8lsTxhckYAipRiGDXAZWDY2o
vRczxCJUu1xi7Pim39p6BiVgtyjpGhJEblFSJboSLxfV3sEEjZ6P9uhEkgjhUejsGN6mBl3+1FYc
ihikdiFEX6XgEiQACsdPYpHeaZTfznGBdbOYjcOQQ774emqRnqVKign8Ypqh7pHZ3upLkibUmYiJ
gR/tl1Gu1YPDOFdOf4XI0rxGY6d2FJ16Xmw4di1Aj+shhZWdnogVgZ9vK4O5BkHt1j1kAOOHEEzQ
ORfG27rMjy1LlLNhGAedCzXxYJs53SEKw437JIlbW3Sy9Uh9XAdxNYiwx2gYx0YcjF20UUnJ3n3y
ekyJOIzhF48Fd9FEOtC7ysbZ982+EXFyiJ6vTCVllCYQO1pyH9Wu2RSpGXqYvIDpe7vyzxOlGpSc
tCfB1i2bj4cOV5hh8kwpCGYUNiF0O94sKWxGMlxYJ4V2hEqEbZ/uSVK9oh+tbVNLq5JlJ683kmRk
HyM8V8u8jv0YwEsg6OAQn1l3pFbFvgBRUiNdSWelaAj8qOcT/1vwSwZ59QAhfyLZp3xljOyhBXNL
ONOg/r/r4FxnBUmECSoRzkEWy7l/OucJVsDXGpgT63QQFxDu9yKIqYo1sL1wjZ1M7ZOOQwfx07/r
wLwq0oLoJvEN1o7EEE9bu6FRacvZLa/H1ZbYDnQUk5qk7C4ao0LM4lac2aQts1tI/oRw7bGwhMhU
oEV273pReTghb4gnlIuDuinKouhCWBdFo0yBtg7oSipzbQm5Czt6Bs3s4hL/FGnJhEeMD37w4fOp
9YAUQ5B1QVJOHg4AQrkZN0D3soiho5VLYSlk6/iLhEXiI7HJPtT8ubkbfu1ErekSzjVVxvfMalDj
hhhPeRe4rp+INTexXecw2jXO2545qElNRQtKrvZ6TKsgjiUuvsr4SLPLw423CMlpwd1oOwciNwpk
TkQH2f64BBKl2tAFyVnjv7irC2sYN4oor9KR+l53eKOG8LTa5LWyr/XiejEfcOyhdYrbzsn+odO3
YWNOrAByDK+MZA+JXnUvzaz8tyhPgcMT/kXwfRliAkZdUDRsx5GPR8xuQpSJ4mXiJ6f++FsAIQI8
PpdEabgtuNtrEL0BoYfFTZ1pXoD3qw7jSyQk1+3TnM/P5hy3RlZGeTjyp0mEA8jyQu7nUZx5Av7K
ShZW8FU6jEq5eS5nNeMwI0DYg9u2gYgBcTUWt6ApM9vC7ppgJ/BLlypx/a/Q4FBYW8kbIvfafxha
Wp6YHWdc1dBmGLGuug3aWRCoBGKHPhzYRL6FhcsLcV4e66ngqb4EbvUgauinTx130ZNjYldWqZnM
ffHgC2Lf0RgsBVV6f9M/WTJhl+u3O6CHrsoWMwkqmH3AnTK168ccBf9V2BF/UX2HvZKgnK4ctooq
xPAmIwQ3tQneOPqvHaRVnJfbRUrPCJ2lGEk5aox2ciMhYuTcOrISI3MQa+pU5Tw9pTNJ8+3gGIjU
Cf+xOU6h+hJck2ShGhde17KDZl0AUgaJVycVIWMoMshZNJYbEbWj0wfP072cUQOXrcTyk1Zinua0
+sv4wCErpeMjVJh8ufM35fxtjSOqqi6h3Z70/5YOLCilFprG6ylozL7S7AnZEF9dOlcwao6ZGPVJ
K0/xTw3+PgIs7i9QAbSAgvh40nN0jdKKgwfb04BkdUofLLnG/PHBaP5WmWH19rNL3gpDN00qpAaU
tcvZQsQvkcc7VXoG/HmYdwYzTS+x7hmab/F9Zq8KqFpxIXYFs6DZyxEK0rNbJjAUi8+oRjBaFGi0
XFpXDBdPII/f8HhvaGOyQoPy6Io4lnPfZe1byDcBNdYsFa7kglKf4eI9V2Fab3Tsr+F86jqCQlpK
e5DRZnRRyWhCvseZFpH+VcPUdS00yzxRE9NyS62QbpNfkBvrR7llk87Kvva4sEnLnvFizZBoVdJe
2dc31v5Mm6u1pjY6qnGUrSx2blM3lzUNdKv3Smii9dTLe8x9m8XLzf8RdmckS/i2MIN/rpGrf4wd
6rLx8IQRH+/BlBBAOmlDD6nne5Rfn1V/mWKuU0Nohn2IlRxv7e6ZQ0D7zYRRVcqQJTU2H9EeDnWZ
RbKc2UjHgN4fClborQutWj9dz3EinCU+OSKTMheZtwaF4AWaXO/WeuaDUnTSsRUVrbQ2fFnmBFnG
dViBGDnVz4qy/jkC5RK6dMmMux/VSJWBGs6ncqKpJWUPJp7q15N/cbCZNrBoEQ0m0a71rbmc4ikK
0ghEtbq+Vmm+CZ9dw4b9jnK8jeXUG4oziRNW5Nb+7cjbDbP8GngY/Xjz1JY2SOuYp0s+Afx9/35l
SliDV/smEx2I6zPs476QPZVvb8Vk5PIt1I9mudXfvQ9+73EAH0wcHcbhuIDs3sVNe2DdxzNuPVsB
vpTQPLNxv0EGTzQbNGwDrtP4S2jllofv6fbL8SdmMsA5KOcFhGFgrLDe0zmBU5LUj/Ab+0jrqnnW
BPz3DFGNB+jxk4q3XMqo5qiJIhtH4FH1hpj7vwjLJ7gnWoNIzpxplgtXL0NpzwzuDPcT4BndFhzO
td0edZsnV6UOZwAA5OTgu5c/q3BtQRYQ2IWNYTzyxzfsDXBBDJhERPYkSnfYdVFl6kpDAEXLWFZG
v8B1c5Zgrk+CvXTHUUMW8rBjc77NmuwTv10XRDcWk19ZAoBJKl8oHeukMvG3Lms32zqEOKbq18GX
TVyCsiE2p9M5azPiWwmCDAT0ozoFA63lr3XSm92geTcQZwFrNjsYNRdd8xkeu1ahTmxmny+SUxBn
oMPeOyC1rXukZz+TUMxA61Oe0Fz0/eJ2cImXdH7cDwsIdj3qZjbr0dykCBbJ2oHps7zgKXKHQYiL
an4alKNxyBoH72N1Tqv/zp7NdHdR+Vl9aQgfYusMPYyeA9MEE9e3vunKwQ5OOxnQ+1C1zfypV3Lv
LUygERXk2miRat37mglslFLWOwKPOt5Y20wZk0+C+9kmfHj4r/arMFiII5f6cDFwEi7RBxRJK4Bc
f+8XZLKZQ/9p3RwRsXIqhJCZIkLka3wcGBftpQlsqOPxoWWgjbaBBSyKawDjcfjYVD8uCtP6sria
AhvFi0WGaZ/RKHrvjWURnCVlwl4A+UBqjl7fDhm3yXhn1Q5xdZ9MZDmvBr/84sv5+4kc9mAXgzI/
ZLu7p6HTrejOaX2gPWxR/30dc/pBC0sE04Ykh4CVQnWMAnEA59gaqc/88Kwh9hmi5RL1HL4xfihU
u4ux/9ubF44rWZ0Qb2YHMwCstWTY8Lb9MzlaGPQoqUCibUMs3shqlli3hia/BzJBibq8XXeAZ18J
fAQTnPzp4QZeujJb1xxinjtrWatNZs1ODoVhhUnWDFYW9ayGZDPWYpge0uIoHpntSY7cqvrqdG26
sJmnm1YFK5Z5/PSTEs+4W0oxPv7Zvw+eQCs42z2lFLaUmUv6YVeP9PHF8/jOJ90fFacHPoMpzmg6
5d9wasbrDBbWQXWVxPgry0rEBnoHFbU5kEHLk2AsvYSVmg2pBTWzPWlQmgSB+i/Wd7TFixJeVlx/
YMEgQqcCUxiCeddB/D8gYCnlfwhQ+E4yXN8N5zOBLblh0qNO7dflZWU3pbBk1hE4dqE1ASKXDizh
2O5x1GLNXDundbbpn3+ATMImZ2SfGcGjEWER4p3yIIUG4n3DXPIknJsT6CDwwhOPxrGRdOCRvnNl
pXuamOjhZqqjlBwwuWj46SnEWgDm7figyM8b2FoqpsLk99Fyr1Ip9Us3Ploi+boEMPsxOsZidimA
8861mzaMUwFiUlk7/VbQ1aMMfWNhsYP2J4KPfO1z8j7WoCReDf3n6yn+XFn5grEz524C7U7oyEBd
TvdSjxw1oMJXwdQGMH1uHhO/SBFY/WYjG+rni6xtMFBhssNaMj6QuA93yeGms5I9R7C4EVQRP5aT
FLYovXLqPsRHrGQ8CipovjoR4xr8ipwoPyOYPpYayxDAJ/GdD69WtSx5ckpGZxP3PqWKwy7pKXCP
O1VKn9nFybbAhMnOX6Uvm+VzhZBCNVkGjXAW/UaPBT4V8V9dlZIIvMmkwmeuhEyt7FAdfUz7I7k7
ymFOsARU3gZjZWdKHJMYj71SEJs99uTQKkTwJu306zQZ/rKgDsCy5eYd8EtQOxCcWQRhcREUz9rf
nY7JMcGTht2UBTOLvo/6NaUUZPb2LsbhY8xfj4XKch6tnUMVHMCl09bJZoz3jTxjuHMRLIgT1+Kn
sNv/nupKxk5CRdYurq4OIJHaT5Z4JwlDBoaHF0lPE0QIpZ71eJ6fbLRrSodMlgs62slRFBt+R7wx
U0FKioBB1QSMqjJKWDeYJ9VaHnIoNQARp9Q3caM1rgX0y9fKU+E2E9fAY4G9r689sWukjSz5OOVQ
M6Rzf89et4m7p8Zp4efdPI4Ec67e4HuwaBYuGD5/teWiF5wzyPsZGhAAdMB/RkBBXJaswFEZyHtA
Op7ULu7gYmxzyxhj+qwFRIb1jVfJ4ZY99H+3+Nl3B4q6YzFF+VuQjtwAjohPQQ2IfMDO9BwKrcNI
AmVZQjMmPmnqBFhm5K8ow4reUjpVNOExhfQaauDizUVRe+NHdi3tRpPTG9QcaGe19XYJ1oqLSLS8
zgy3255Xk8PgIzI3wxHUj89KY9bXCG3HjZ5yymw3Okyu45jCv8aQ4zquyiIcOTUFXQaPnYJnQ/6z
WCsEkT+vTJ6AeT3dzH4xjAxc81nQ94uEbZ2XzHhP2O4sC4YN10gylqpjiG3YnzrzxaaqmJIfUPZu
pKev56gu0NGZaSvwm4ExgqewYQQ2R/kpZ/zDa1La0fA00fOiwH8xr9IOW4Oeka4bO5e4kHAFL8Xy
qH5FYVHISVyX9V95ypQ1BC3cHjsXw9oZzWzmkCiGKU4zO/8mLSyaj1bmhk5nybDxEHK8c63V2K5z
tLRXhjXp2+5tLgpDnv/U5mVvBc+X0ZySuOxVnGPDejN3/BKM2cEwoZgpX3YImRwQTZY5zIZ/Z9kz
Thbxgu1qjzVeJzTTWYEJud4OHiANLyLDXQwOI5E9FywFZSxX75igjHIzSLrGrDRk5QmtZLMBJ/pA
hTzOYhjsI1/Hp/vsePPuQiXQRJBrzx41rv+Vx9mnhLSyADYpiwupHJXKKc2mTkPvhDhbYIhQ+fLo
7FPAEhSplQT2RLqZ+Y27uJMNgT/H8QJlgAdkYAwukfNxAPT6BF65IX3dRNFSjXFDUZi9drY3MekO
LNW4xfaMfICuEa5GsXsmLNGmZNHnqzXC/aPmozWF0oJu4FXVKcpfdufSeiBjZAFeYrG1NUCfSmB6
hLyLq7RWYkC2DzTrS7V3c1tNGQI8HPaQkl0QoBHxVlYFEJ0uVjVhCi+erXPJW/Ypc0HDM2tO0fQ4
R/UGabVbqIRpaAVPdP/EDddg9ojB8k3OZByMAOykzaTAlGuAkmsUpxFEUqSbF+RqG6eA8/9dvOcq
DGceVXnBx8Gd94L0ft+BuRdr5JrImKJySC7mOQWu5tLUqxxBxS1xhk/a6RvNuJ7GWj9LD33LJ2Gs
3bBhIFiE9TrbZp2F/MJ6+qcfQMzTlXyexeOsiRElJ7s0ka+EtYARzIyANM1auPbo5aL9ehyni6IM
0/JGZGTylT2nK7llXP6c2FhlryA+ekNxAk20savJaJNboaAkGn3xbApHoVvGvZMtll+KGjAwqTR0
BhWwARQYAvmzZ7VRBkMIEFwaDuu6JN4Y0EgAI6+wAonC3G6WLD4/FbjI7EnN7MbeHk49Y4TbtqPK
+UwN5Oxu0zHSAbYtp6D19TEmrg4uk8tCPE+hFFo7ZoSjhzzEk+we8gbbvI+SNfXapH8nPrv5ck8+
F+1N/DymBYce32GZBxmXV/4m72TqGwbu6TBHvdS5kC0l0tnqW1cg3KLd5i9ezz/qV/Op6272tAeD
rEcwIcbC3z0fxS9iKvHqIPAryCsb3ZyXMw1k77F8axefW/YG8CrDILvpknHvylfTpvlSYp3vcDTy
HCkBmEn6UVMQDIOeBKsHFkyw/AbNnQw5x/CUm2Amsv3Y3YIlEyQnufRHU/gz9Ej5Y3ZkwIwvFrJ6
tlGcoQw0ttRZm+z68Mucz8EpHWkzcRctAd1yw1qeceV3F3HsYLagzWg8CwHKGHcrWFb4SGST702g
1E0WxD4+l0C5wYyEs4kr4eG+MLzT2GKqGis3hWeIYFQNuxQFro/f0iNAvns81qXa38jUBWeKlc8a
ez4yNgpp4FDFBGZ5o8fBoQsrSt+fs6SKVVc20h5lcSDuwg3tqRL9mytC+IaafmzZP8QZW1D1c0vJ
xO6FYD5nLHFTCAO9XNg7A5zuI7HafxLQBt8unFFTqwJdcKR63F38wMIJ+d6BZghwBCWgwwSgGGUB
+opxBfB5lDGajvx6dFn9RjGBtDGsvlBFB0WEcbJA3RnfI+1mSfNZlWe1IWU34KPsCxhTb5y5l5Un
gd+gZHE1rTuh10zkmxwOaLI/KoVo8LzIJt78pioBX4TZj9GZQusFPrUZ3vo0FUOpvTJnxyaiFNmN
rJcr9MVq6UGS+gmNkmETVB0OIF09pywlEIRwfGbzwyna0S6TNlw6yRlseEu0E5fbxlwAxV7G6fXm
YTOK91bzkSTrl0WR20O83rFis6cG2WWzlaSVH9o0PX8FSD9CO85dcvd0d7IR1R01YFt35f+cBdKK
AQk/NslYIMEvx3JA+q3hNFbfKGc83FzDH1cSzKZRSA6EcUm3sJaudL0SL72DXUmJrwqhT7A72Sjt
2EdyCcScXszdxwNHESGXbJpd6ZNqpeb7TKAkLlNUjTxxDFOlOkOSfcsQBEISYedzCd7cfQ4FEsaB
cQ8RnMNR13zcTs1kOwhtLFzwW4AfAknnMNZbyRMCKMR/sSdsDdEae7kqxc5UWMq5XHin6E/y6qZc
OYvymzKdqmM3R9KxR3jc5MZfqWPKTIEw+eDHWITu/OBr9gXMtAc3Z0F+Cj+RPMN2rXM2RF3t3gqe
sE34UcK4Y7FJelT27JKZjpF0pdlOPa+O50gypDVoM+2Jj24xgeIKlNrt0yWLMCk9Kk92Lzkd12W/
Lh8M+98FOJN3LvpVEegHq58XUCiXasXAh7Rwdf5oKqVeNKthkxOt/PuE3YqPY+8BGs/d2u29HHbJ
62TmPDDVA4i1capJltg+z0/eCWB+gw/ijtcpx4Tug/CVfTLUqhqlyJ6xJV1Xjj4WLXFXT1MuuLKc
qMMUQylrpCb9cP55MWju15h+UeVMXW1n/8S7o/pvvJ/TU/LsAC10f67CoxdPeK+wlXIXK3WTyCwh
KsnWnngtZJPQDw5h2oy0fhv5MWJuBAFuoPOISk9ZCBRMe2Ih2/vv2UlkCnZyY9VpZNM1u1/Cdm57
3QE/LzHeVe7+TOp+W/fDmGQxuPKnn4y2gs3xmcgSLmi+zSbfL5/rrBNxoeBwZ4MxMvbbMqbL6g6B
4oBZcptjE00FMkWgrabk++qO5a/k4L5aFyy+r1y/WtRzPat7JFJrrX6cAcCPrgepnl+IPu9640ps
4E9jF/lS+dyRNgBvIUYwdbso/44OwqQFf/PhEtMto4FYgXiSWoRVXAQjUuQ0TPAhIBSUdEWjqO0R
WgLCgbfHvdbgT/Qj/WItRtDrt26a7E+sVgBoxINT1zcNz4Dxvx/jtuh2dpWXEYKbrmv+u5BmcmOP
tDRKaWEPkcLr6qkuPLJ56VcBqAWyGmgoyyaurcMA44jmnjAoWjq5PgyMUeKBgHxN0s5A7AbcUTtO
mSUUdOeutfVRwd/IK6EUVJEkVB5c45uRCp6zz5a+BMMZ8pYwDIkaFEolHJ6yXKpVvI8dQrraFlp6
+XHm1oq8cQxiVrMAjUQ85NAsZmSN/MtQ7w4jzjsQAjhAHjvgr+h6YOlMj7zCKwPnfzGX9F6/DRPf
Y9OstRMHBED2XDdGaxYAvDOLWsujss+7KRGNDnsi5zXVgw7bhTv8ymZMx2r2lFL/G1KxhGQt6j0k
VVLSoabKkuuLhJ/eqmCUrY3yVR+BaQdLJdMFxDG/iCTxmYCRtMs9OqwIw57eY/5hwU6WIyEVG1Ni
fHKmgGwg3zNH1RCrqGQHVg/owt71lNF9BBlEOrlq+gGfPkNRzo3uazP35+M5m45eZlmYmu5fh5ec
Tu7JSQ3iKkRatiTP9ve58NYKSnirvcfEQvudtSI/GvDCiDHs10HZKjOfgRiSKXTvUWqOIbJT5Bfx
f5kdT60FgB+dviokUuZdybewbCIlySn8N5P/0dCbSXn/CdZHclt0Y6v6yokZh75ApKQyI3fmJ3kL
3PdyexAUOe0zZWWLS9x0pV0Zb8w6XZIwTyYc9Tqcczi6QcbbxnV37TxpdIy/TqnIlA2NmhBeDXju
K8AY3vk4h765Cbeissdm+fQuhHrN3uCYny3aHkMBt3v51BfKJWEe99rsgqLcaWHQquUF9i2ZF6Bk
ynJVxpVuTMt98qfasuauWBaBHrV/VHC8gVWO0Ih/lKbThbGIgPo3QvJ6/j6MhJQ7+BJYsrUToeO4
z82UuUyDNiYp54V+h42kTCm4hflWWooomtz56ADNFuQPJl6tPxufdHS4Tx6Syb8AcmHMorgHsLjp
J+IhW1eDDED9bYS5D7EZpMKHFHivR5WfTykW39yi2tpiUIkgdEbuzVZXvwEwB45lWOZltss/hlet
YdqVLex/Iuf4HAMSyzqL475On80Bd7PjYQjQR2t+2Y8E97P4bxU4lqO/AvwejsqchH+ctp1OJA+A
hdEi9kiMrRSpcPPN2WESPEW9dK5nRzBJ0wtIFrAAadF7jCzoqvj8PgTIDq+CvAr277nNTKfyKrC0
IK3d7a1AHbtzdmcqP8NaVSj522BvRwrPteXzfYXyjuWGHpqjWydfOZhHPLnyU19wfR/hq8vztIDr
9hEwoB+dZCwRYj8RjsRjFrHZ3GI3SR3U7eB+M9+kPP9bfITcPkS5cvnxMeywDdN88NzdeTXZwWpm
WDciC0SVvCUOV5tDy0msSGcBZ5J0UQZayr+GBPCoQWrX+sdOVMReYtUQ5Mp22tqc61yqkcLp9so9
lJ5zKwKAvAgoZqtgU70l0yBQIqZou9XbDo+1nre83GfabuaC15Jl7kGQt30Fz9nYnYNyIxtSWYgw
8IOHZfthlx0tRTv84MCmNN21uQmi5BPTYKCPqi8XBZsgFDtPnpXF+Jgo2utdOZDIfdaGMWgcFeek
glYB4mpG8Hte33xpblJzWjPLoSQiSpkB9lFmIHtoLuN9EhAjeInkXhcfch+Wb8CdjDcVjcGczLXL
hstqtHSemR5HdTajIumcl82HXLlaQUx/o3gQxDxSsyXKiRgRS58D398NrQOJuHGy71DmitenrT03
dB5a+LDCJ/82eMbtMrgVqRKheqT7JGHVGvKq8z1RiRny65yDKejnbJ89sUZo3qIwcznxPk6nZYfz
0nYXcpvSAuAMl0qd6MsXTS+cSGooeSyPyJKkScCk6xMx9ZH07Z5r42SYEc7R2sgUzeH8PywjNcL6
W+ha//9mycmjo7h6z9MMkUqrE7rZ4E/lgfpMigACbzhSkiE+irQ4om9noRyygBFiW4IAVMDcyuNV
iAe4iSFxUsryvThi7iBU3wWKrXqbzWW/YZUlESApfRLNZymKyQQLxtRnKQlC+eHPMgMP+K0h4Jbp
THrX8VjtxF/viGm3F4+XWUK+jsJytI+66R8WRkA329LL4q09OMB0qAS3eEKX4xQ/CSDXVsqiEiZV
D0mjwG5vqOMCSKCCLca4yFCmnpRpby6GntolUhkWdyqqi9H769638q1jf+1kAZcep7CGASJnDP5g
ExsdEaHueErm9xqXJwnCWIl3rjuFX2KO3t5dkxLJSHZmcX/PklwBOJqoj9vzSMh/NmJtgKNr3HM6
cjFb86KRUAkKTl03v43O8+/Epsl4j0GnDzq4OJYyRrV7HWVx2kTmCcxTryc9LgMjuZ3kiyhmVJGR
yAi/Ayd9P0BWyYQ4pvaCB7fW1Szyr08RwHDdeq9Ahb7I0r6qEuNVAkMqioBtWHXTJxOirYEHviHB
n38dF+knDHsmSZOqATSFObDa+pWDMTqGBZtIzBvs3PJX/JcmjARaVyDSpLP6W7MwVp3gAoeNbYng
udy/4ZzcuddWRNA3LiWyAOwtpOGGZ1u3E4eQJJe5aw6roBkLK8r/gzqcK1Ug9303nsAvRs1tnzjQ
uZYJfFrM8fiHNRRfrhW+tmoOHLhKfh3wYsZ6WOzQMWE4zcOhOBUWf8+qe9YUepBS87GAiCoLgu3t
PEEq20Xc/hIMpG4whxpOMTqeLG+LwRevJgCb2WQUFMkJW5SBNiM/1CCRdVcYjD0srn/uzinZinNh
gfiKnXyh+Gxe/cb7doC+IvCkIwEYCKJ6uSZG2/+OMNsuWdlkC24seEVJcdSo8t+wkMCvpLZYvDH3
mS7+Kao24RRGqWP9XAL3xZ4p+xgDdT+DPMvo9FLr6NhWPhNWs91qsM82+uijhrTcKW4ORofJQS5d
5gpuNuMT4h5gA+vLhgqLfZazY5VhbK9ry1UZgl+1M/VD3sBvyYkY07CMcpX5DAWeSQcG+kcevhrV
um7ErB6Ks6zbllPG1HgqGlian0pVlC8sRjWkw+Vj8OZLCzL5mdm7/VXNdmCpggTig44C3IWSpjM6
Cv3u9dLiZLskeILoay3VrRX9hGJsXSU0QrWoda2qzXTNJcQqcLB+mob5XEZf5kIY2PsLsrqUg3sy
Ac8vET7mfCephkXlk9F8bUOkIhcyWzumRLLTsJ0nz06Q3YQTyR33W2EPapXEqGq3Q5M2hoOUq0OC
beCWcm3ZxPTdK7u9RnOkSOmY8hN9bPLaMyE6HmLCQVBH3NG7PWtlz+zKOpj/o9AfqBaQhFgHN+XI
65jSW5qfgOZNLzn/7+DONCFnMdNI5ErtIdYV0hv3i0DEfbzNszEK/A2VepF3iimCUXC+6Z0zakeb
GiUpz9Hqy+FP78e4pJxokCJO4JscSdnR9Dydox1ylo62bJJHgVLyooUqsP60kg/RiUEdoUQ6wQ8C
6ommGA0HGuDuIAGg49iNVTctv/lwH5kz8tp+nkWcYghJAk/RUlHeQz7FRwnOdYbeb2zRf1mSAbon
UoVPi256lKC+gw26hFd8mxBUwfXNzBZ2xOq8dvawJw8jmg6w6E3v4cLx/ttyzQ83OlkxLNPpNnX3
Sl07FwjFr31qilKuIJlnoBIRkEIvWcnG45aH2XExo+VPGEMEe6r7+1HfQrxAN+U/Df2AmiHKTQxP
NloeFVsCyatCQfq0ifCyGvX9jLB6fLBxl/4oQR+B5vVxO7Z5oIl6AKyMrkNpJg5aVL8iaQxtS3PG
Qn8xx8/lKDACVcb7LlZjMk5l+5JqVuqrEI8erU1ZpcmfL5r4vGh6v0AH69RbNb3nbgjsozy5ES7/
9TVkkSAOaQYzoIInNc0s4bR+UiUtWcyFgnAhXweLVpPZRBd1xlFxVwMMtQTcG1MKHbuX62Tga6eR
aRpLDGod7Dsxgps3fpyBnQvJgdYD36bDK26fI81JPtK31c2csux6ojfBabJ8N0N7C/AKfMu2EY8G
8MzyAxSqJs0SuQ1NMnWIExR9hEdNcyDiY0SlgeoESJy10rw459K+BCjWcGb1Z7qZdcVzUYn3RC7I
3h/AU7XjHyYN+mOlA8MUnu562vldmtwzwZ+Uzt7qINkKeNQhLXJwdHNcQnbriFIBx6PMOV6G0Ilm
4ZjFioI497uhaw5gTW47hDvq3KFvIUL/kc8z9AKWVtSJPhsh6haofPrHqvYj87QEzRTfYuRgl1ig
HRLKn5tAgeViwLyP1Yfg+ZywUJu7/pKZs51JRjfHP8hGADV2K3PY02cvqCDIMZg0OLQCdswZFco+
av/kExMDIudDojY1+F7v6zZ5yZrfKTxm/mJElpGKLwVodQsdp3QSfOTUFFb/M8aomgd0bqY3R7VC
pF/A+8wG/jBgeQcvEcgH9RbKN4lBP4EeE3e48IiNlStZ9easn3zXl2n2fk8C+TttIXEHSGbio9fA
X4dtMgGE/8A5T/KYBwFi4Vf9wGhqbYnBc5UErkzSBnLigWyFjjlce+5LY/CdGa+NkxvA77tovN3O
firk3sNo6dDjszcZ7AxGMfW/KyGt6H9Zm9h/SvhfT2kXs8QGEZmwzheT5VzPm0CYtPCMeI3nj9FK
aRvhF+zLvUeUofpe7Gq0qfX0gcP23B/0WzhVgucAHA5/02aWt3gHv0iXpipb562A5kbEXTvBM5xz
lj7/KzDikTcPZN0g0x84oWlwHBfZ9woWgqBG34LivZVxWToeZ4iWzLRFvTls+T8zV2gsMhBRELOK
dVgPZUwGwmqARTtXB+ySqP0PQbm2PESQZkfR/ww5wb5SNtOaFAm1ft02AxALJ+UM/AWOT+mlrqtE
plKrK8eN4wJTe9JNKfjvQWth2/EWzPGJPYPdE7ue7ahKxLK4YLCnHioPxjrtQ4HmsK7wIU9PxsXl
9Y+qKKVe1yOwFmJBG8ELTd4WxzueMe09J126LbVngPBN1SU6l2+NGFwCBsjlK8xUfFejnGIglDQr
F6peBT71ZAsLFxcVLk4sho1Od5b6p8hR5H4EQWlHAm7iaWneGxUX0oAPqPK1t2YaYoDlF25sRHzT
C0DXbO+iKz9/hkJNtaLwy3WTCrkIQGpKAeyMFdWVWMAOUlHV9dMhNittyjFAetms0yeyiZZbpiMI
CIGkjuaPe/RNkAEd1lFPctZBBxKz+apf9fYk1u3iL8c4jMnuK8Lm6qWBxj0y1WdmcM+8lc0T0cyu
s5UlP/ZmbiWQM41goqw4Yd63WUBt++7GoOevDSpfskEPwtXx931BCI/kEEjaPsuOUjIjwBjGhlNW
VTcgTGqfc0c+YUL6Qfy+Hrnrd611B+5iJXKm3ooTQzHHs6ylXzosVYgx/Wr2SzrblqpzYU5Kgk81
FzpJrKjsAnF0xvDiu+SIVohMcGmcBtthGayDcEpcS7zHZZjVJHwN8KNIdzcCT+0A7hkiuRlwt4Xw
HeMsKVGD9lnS2ZgcbpuPML3+p9pnwwQMqQJw54ApPKck9F/3T1vQpgR3eMaOX69TO/UNEzZlKPhf
h1At5ZmCh5Ki3U5f8S9JtnZXHhTJZsXgaDnyOfLCX6unbvhvJCEcB5XVDUs5wKNDpHe1/l8Hs04B
Ws/a411mcoxvlq5WKAXtaXAFrWwAQBFIJgZGNNDJsqTpmS9qk4MuBqVmq61nVN0KOPjSE53ZrwQ6
12ohBdiNZvZxHH5hS2rasexuyrzjTed6GlcxqckUyAwv6Mv4jtlXXwkmBGWijnTcONccJ0ErbCSP
w9sEUrwzUe0q3NB9RUxCwOZGLly/FYqrEgrT1RVMsheoPkwgln3bNXBrRPVeWjkRjAspJqiM6fcZ
WhLOjFFi3aSXhwF/9kE7SXVdDFvMnFpFovab8+7UfZwVmfDVFymrHltX9XcWP30s96K/IQmSGU1S
CU1rINGDuyKTlkK4s4cZ25QwiR+FWALSJ/Ky5/hqDuNGab4vjbbdfE56IPoGqOEj7OXGdenaQv47
4ZKVgz5M3lJJ9I75W7D6femwn2HYEkzjP2K0aNlEN8xa99k3ZISTinDFnRXVcuQqdNV1KF21ZAUR
S6S2wozhKiAU1NGG94yfMefligTW8m1ahLW5YHkhVvqACToWJKkry+KdiBFPJUXZlxIrfVRGLYjQ
NEhkNNdFaP0C76TpFv0wKccaj/iDURY4uvZZGLvld/yJPB0GfU5t7mutQCla8eCBuTmnBgri4BEQ
ngqn9xn+eNSdSfqoWnoRyegsAzkAd3cAjMdtqcF46zOOUEyw8SKhnSl8PaomfZky0bH+mLG1tY1i
l9FPjn+DWhbxCottmHxyRebV/9sCCQzYyQ1pXPSuxZB7hmKRZdHb67tmstGuE76s0sXeNkoz/QFO
KQsI53uFQBvV7ZxQZwS2pa/99pdVyZhrGUEFu+07E1XCEocIBj8QwH5JUaYvGjucrIbhhD4xKjGn
urL3X1qL6oOWKk4omYAIE8y+Ax93Dg95E3x6uU8+nDmwKZgGXhTYYWEnB1gXP0ZvOwYbLfeDHASZ
Uh8nlZ6AxvFG3k7o1VDNAQKsnpcr4OpEJQ/gryr3D+3ylR8v4HgqVnEGYrmBcolaEiohbxZCC4BO
IiOQCa1iNOW/w208nIGWd/3hCTbgF5QNT0hMICdJ/KtC9y7hbeZwmPXJDMbHPeg0XFU3j27+aakj
Vc/5kRvd21PNTmOkdE22EbGEErvgwoBmGXx2rEYNOnS/hnqVmaUzul5QFhz0bPWyKxLi1k2mJZM1
HYoz2C89dULe6JtXGL8ESxEyTTBv4UW10uOGsuwnjmHRv0lr2m6FkNfPytiP+OHIzqQ0bCHqFiRk
Sve77yO72AIQ5UhLIZ1jvVLMKBIb6afT/KVRyqPvtu3/OxmaqhAdMPtNguj+XXVUkwsvc19syIv+
ey9au2JOAqQprjAuqnTQFePJ9PBX/sYZ3nTMcDB6EyLwn1Is8tQSny10NyNR/UDoiGQl9pp7kl8A
9OGU/bPLNlg5raPgejw8b9dL/MptXaKP0tKROLa+eukUp2LGXozABc8ykwugERRO1la7KTz2qUIo
MhAvEXt5oiKsGIc3grHnwvpDOf6hbSiBNI4p+cdgsyhAgYwl3kceoTnB9A4R/0AQ5oTRnVV6No/2
8JQbakg1JwL2ifxLIaRg8FCreMbaSXqYEKtjzeUg5yKULFMlWcFVcuAPp72Tiy6x0td2pBOxMEQw
amk/cbAwCx+LxRPHGir0EyFe9jdj3VqJZWjDfmWbcEYMWXpa03jE9GwkodoDIp6mTeXhBEaHFtd6
K3lcKJeCzccpxS/0u0bWmRkbEZnbPJpTruFHULfqfLQrHnyiDUBja0AO5FcYbKboMOiXPtTqek9q
T/unjf5YY+cDvAMxwz9r5cq7tB7PYr377uvcDkERQ1Tql8t8Ah4kfVt+6HznP2ltCtbtRAF6UrxF
A9C/WiPL2xoDqtFZAEBphSRc2q1sIf7SycR2MElkEL0BJwHR3yyq5mDXF5WLMGzAuoS5xx0cnnRX
KPgqSaqkZ1NiMv7Oz7NxQY3RpeTonl7tj44yJmBFBwFr9Rq8Yr0X2WsWZpV3H31IJ04ki/b7wOXl
zvRrRTien2W2An8QkmaRf5ZgxIDXcxz49BYhI+pAfjyuF3i66IJYnRFRxYuofPrOdbWDjOILeFxs
8tSAQesdjPWyXmFsm0B2jeYRCwLPFTIdT/sGhIcbDXOq9tYc5GSYGR53l6wlV/4joqGA3PU9B0lK
pByKiLO6XjnmaT48hH07GU4XYxp+sgXTeOzavwUvUHrzlVviQHQ2qEV1VRF7/YJjJ4VkviICR2lR
5kE5Et6pvPqqZX+npp6giibKk/2UG7Fk8Mhnb9efmqv7I01tprYEzqw/O63NKP8NTOsHOW7uUqmw
zjUsW+8g2iOfaz1DAymTOigy9UuU/dhrxwxK6aDMkQYrWqBZg0JlVMq58+pzCMU68jtqFmHX+eMe
RrBrRr7smKJXPTsGCKXsAVz68IQG9L/VyNKyUuRR+0rvJi/LoM+2czV49IUVWSbSSbOy9xIeG3Qs
7Zh+XX+feivk946+kmFxGVb082OMgT+fGcdbGaIyKE8OapIV4cI6STMq3YRdqs+RdY5H8m8xNB1w
mRzfB60bjGfqMYxOkNc4YcGgi6JuYkPFTi05ReAmezQ5j2yWmoINlKpKZjZfCf+LKRZaWgNZ16vn
FqKDgAL43M4CbOkGiFov1O/iwc32xnh94wO4eSQLS3iVjXCe/TLUsssqVWMCN1+4LCxRHcZK8mW9
qYPVs8RXXeP3AA+XosuHrm9vzmt5xdCsSlevYgek6VqmyMoT2Kp+8ia/wNMe72cSkm5BtARC3qo1
RcmWEy8XW17CdNcNPsEsXSc+Ups7J7+nLv2PJFjiMJ4NeRFzEO7/t5Du7eP/eEDv8Dw0q66YYkOJ
kedGkYOHSxPit+R9z/8rhMYd4/izulIBN8PzuvgwyQGVQ9V3SkHQA2nbw1Mnlqpbn6j9lPKWVR+a
zSBTDlcgsNZdH2cOCW4hyyqwijGMkCK+nEomHeSbwRqM4fLO0zK2uEpSCwXm5MXbTC6P6ZYN+uiX
MLpCuE+rDK4R1NKxwr9/Al1TWwC2vU5zYuB6WC9BXDR5UvPEDU7al6oZTuT43ne8jHuJnq61GEz1
nYN2e0jOaKhCA1jTQldLuBPY3fXtsahGf7EzGRgtdwdxm0A1FTQ8TJ+pEkCieKOXWgbryeJynpYi
MG+z/1bVbXxgc6zyHmKB5L/fWWprHOWn8zPxZ4wpDBW8WKpw3rgqTGbdBaI/hwaOK4SNm32lHtTy
cHNzDs34fzPJWVVi8uG9GU8ICfotIDnbudy+VuNy+Z6sNOUbBEuOcj494avoXgJMbxl6QLkqiXAt
t6kX4rgJdQz3syOqNtj5BqfruBmJo2Bkd7oLpLf48i3qFGWAjiIxirL+S/va/835HUj4XwjqVs4s
bhlw4iLrKpxD1+0BGx5ceK2uQDXNSyWF8cD5IEfJOAd9nJ5SZeQsguZ9BtC3rIuYJsdKY/DNukzF
r6eZCxOhCUOfD3i7+WpAnmz8Ld5gSdEtmWOUP3BFpK5rVY2cCsftj36OXQL1nsOHkgMEoEV+7XWs
CnCo7rhhlrheDmeKGIXci6vxo2iHCiJrYctQOutMDsIJWMYqFgJSGptkiGdB7xqJdCGenLkDhat/
AyYW+PTwUgg1kxSoXehpaM7ZQ8LNStKuiK+ZhkF8w/X4zxeXM+R0PpqY+kRRfNAfaypDEc4OReQM
G9Vr98hukgYVSkdCq3hfK1lsndNPs2gDUc86Jfx1d/5smuoASAjTj7fW4iwjxwGuDSzuoTC+2tU1
k+J24STqrwRRNhUzYMK8rm+r3m8lbpuy88VG4ATIW7+nICrEWeOH1G6uoTxD/mjljO/CjO1jbWr5
7gGGTkBUE+c+njsrbvmUPl/azARFP26sfoksHS3TjYV0xizhVBhy4LeUaNVhNlbyBxuwhkvu6Uzb
tEAGSdGgnib3UGQPbwbmbGPh49sOi6bDJWQ9yEiRi6Ec420hc7tIAQNGxmkNf77Ar/uB/K8045Ar
Xgfb7dYyYsRF6vyKT0meu4HnJM7T+7h37jSw/5/S/Bb7N9ipeERpsz58wQR441XX7vYkVMwGIM87
3vzv7RcD5ANQ+99B9f4jRboHVGPlES9APFEUArmojtRfDnIVBDyNC1F0nJ9JuVdUuePQ5X+l1uEj
g3FkFJ/kp/1EvY2INtY1kLdSUgzz9UA6Nc5kD68HzyQmZggx9zjEMkoKpF8TwZYM4tTI8W4SvbRY
/tqZmkCkn6XjkUl0M4sWNKcIhvnOYNTX9fMFxx7XAww0PnL2FrcvglmE26avSdPjkuEf7JaQtfid
P/YphBbmddRl7PyXAl8Xq1sCux/SSoY1rmkVIxKgIqyN1H5qikwAu7yjCib3nF5K51tigE9vahHm
Fss1wpNkREI+QUUf8OFERWKzqIrsJxeTtqch8ELSvhgKqFX6ZbQSRpux7rC86ntAqbi4ox/pI/O0
aX9dv2iEuoWABRl424WmJizxqgGMCt+rnUdXz4pNI7g6W/UAN0BpwRz+R6wvA4sszdgIHcNBBknM
euK2AzjOUp/ieHzhEfyWu/9rtsWs94S8bcvMPmE0lNykY91L0IoxvECyMmVKeJs3yNgvWUHEI4Gf
IihrGNlTlfh8oyHitmvOStSfS7CvDcOqfa/uyw+8CxvveoqTA292YgAuR+eCJaRHbsr8XifSQ8HQ
28+NNK+H8W+txmcZ7Swklis1lDY7If2hJoK+mBhMX7MZR4cAvwlJkLOLXYxAxkjTb/SBnSNBGQZf
ESIfHmIig7gJhG60zW4A268Fl757f8H5oJIyawLaNHZqS9XJEd8ggSYsZ+SZW9KS1dz+5JMVto9K
kOVeF7LiUhTzroE/zD4mkM/D//fC9a6JuaNi7Jgut1JW6hsOrTaHP5nr45XNsmU2cK5IVnIjkgRR
4SAzNM8sCK68+KWdsWsBXGeESF9MXtbnVk27rzhPqcjbTnu7EYij8gnNumgd169EzPUpkA9p6wff
mWGcewdVwNUYvdqpQ+Irmz/9qWN1Ofu9tuE++0pLRJ4j7SV602FdHq9T+M6O3ATdF4XS0xYNHvaL
mjIurgYtdPsuFokFJa4CI5E+IBr/4qlhtfwcvUmWw2YjCnaJrOH9kxWqUFVz1IN7mIwdQtalC0IB
pG3+qKCmR1MachLZYlzHladf2zeLc9XfrfCrOLvwQRDZVCobElaMfuqWvf4lVTVm7ziJ1hTsOrM2
dWrTogD/xTRvJDQY2IBC3rlQ04WmSW5j0CiPLz9UK9riyKHXJ1uMDM/m+Mb+C10jFSHxp3pkUp3F
NYxtgJzXvv4WugLpUPnQhOzi9Ohzew9B8Cu4ndyyGVNZchOKjvP0Fgm0oOkJgQ0GkGnHsw45TXbv
jQvmOWyp4cDmGdoDKaXC/YXLhP8W/pBdBK4OBB+T2cdjB7ovKUDMiMKjymK92QjtBuuqNE8+MCLH
gAzoLkyYwuGjQl4duDeWw77XhkG4X+9k+pfwgu0lwMZpl9WJ91BkittUoKgHfG+q4kyR4kGCJ8hU
XtMoNKaEVm4Gaqpp9HsCC9VqN5yidMan8mHOKmBrm8o0/uT82nJM/C4aj1uhwaOFCmKnKoe5g63e
q6JrQo3zhMw9NT9RypxDqF4fhkK+aYDDe548AT4soRc4U2IpSgBh5yK5FobmsHmST0YqYx1u3JuU
98fKMWRPyspmzlUi5P7h7tm5FNcAFUemv+MBaBIAD47fblj8RJHdtBX1nfGNJYup/XCS40u2FkYo
G4OgkoW04U39pJcau/mJ0IRq1vlspUfRkd+HgFG4NIsuBNVlWjbeF6TSaLaLT5hxs+j7+BDwLq82
wdiZ1jgAk0o3lqmGJc42KDhSh9hRrCpj+lCjqyu4vULySMorgd5YJPz/WukCce17vGHEQfcy55VE
opp2ItdUHq0gaLyXE+VhMsr8Q/VvY5USkd/vBeRJNAgzYyabrWmYgdPo+4CyW9GSo5h0jRK15Oqg
2EH6STvxJq+A+VuzDGdD/7Jc8DwkJp4cntP/KPpV/yBI7SVWc7TBmgSJYh6U2Q4IsXYq1ZlrCKN1
R92gY84nxN1DVz/UbAPC+g4H9/HggupJrAF7NEcv1Ge6fC4fraODZtP1CYNmviu1cgzCVJsBFlro
arbsqnnwNhJVflFBUysKezsAVLv01S427kyy4574iFSvDcaUkjdDoB9UWiuq6db4duyQbzaeSiwN
hsZYuk7yYWG7bLAWL3S4+Ctdi2Uz/8G4wXfDws7KNzZoh16xsmqJosVIgFaM1EeilIMB5sbpCPqG
qMt84X+S2TnkoTWdxctJKhu9AzPOvJeMgXAU2l3ZCTxgikU8ZCpYyPkyo+V3pgHAdxfJnhziO/8M
8Xeg+eMfP8CjhgAW0BfwIMY0gygGxC9XknigWgEtxb6Mmk0uHjHFJ9H0f+CHSJtTlljxDWq4RX6Y
ypSQh3fyFk0v6ZPO2kKHYnt3NhXLaWNDg+AEWNRhWnVxPcHcuOVzbL5auefO5B/JUWCFjyCKcQJH
UdNPtwY7+8L/pJUyV8mVDmo/13yEf1s5bYkXCG0DsmzUI51hurjAnpm2R1S1vbahb5LI9huUe6WA
Go6TBgUXFwUBjvnTxTZ65tUoFII6vWs/AY+uqGaxSFpGI1JSRgVqdPar3btwl4yrL6zwNDfHkzeg
Gh/YSqKCTaY/bPAjJMnGkhriGWa2Acc6xdtSb1Dr4DDUXFwRzWoItvDA/9PKQOgvZCM2YC/jaHaG
yIPTE1al+9xI/kDxxB+vy8QBWqvvESszKGfp5lt0i3EotVWa22TZgiDCFuV0ZUgBI/tX+g35jbvX
RMQwj1jiixFHfQ/33jMtENwFLnouVX3XblzL93VBRLwU/aCL0ATULSk32MPdhbl1BsqfSZL8/QNh
VeNBLKi5A/tCm6KfdDswxg8YKxLRqIsFKts6AXndIdrO/8TulTwi1i1ZRfkqEGUYooHjY+JqZJEJ
aACW/KCvQ9TsLZ0cw3aYT6mZ/1pkqmCOrssxTBgbPHBOEKrKIueeiKszpyoNeZOFwX7SoRGXOXaa
wEG3oxtc5YHScp00s5s21b1Yxw+j790/3zaeQ9fOHZ1T9xRt3eSKQdIg2aS5BJN5ZlVHSp5fMkWh
ovKznbLXsabUwuqM5TVGPDxSMVxZQfGssr7Ar5HH6VJbwEQRkXZ0aitiOtOTtlcR0dvJc9njkZ8t
dGTtK7+51R6XkH40SqX8ajgIC2PTVlzFWRuaDyyTkvd+55R2eIJJXhNLxh4xY+dVnTor7FrBMg7b
Fk66rAQkmnVXGmg1YYR0N7u4yI5HPUSPC7O+YD+3FI5yiyG1RWG07TILCaQfU81NCNFR3RaLctNP
+yTE+4N9BGx9Yo6IZjKXBgOgbOwhqkoeH4q1/4zDd8VD/TIe1RiyE/mCO/moC/gEekq8CzLIXMh3
4KtgiEgNyUIXekB5NRLPkTJKzmDE/ashaYLRqAVhVwFJ3J4+D0trRl51iZZLyA9pLuftQ3RZgTK/
6ESSFwrHax8vbU2GQ8gIczfSZnL+QwP2cNSEHdFx/3LNw6ssWP0smsDmVP51iH9wh2wLvnXm6LGW
lxR1Y/DgEj7+FNw9nYPx4q5yT2C/MCe65B9hwytqPQh1mZcqDHGxn6oM1Vh8ZsQXZFmiJLpmzvAE
1WjAGXo771J6ALZsUV6d2acz9gK+Xf00YDWh8FKDxrxUTr7T3OvBXEWCMvhzPilCciBwrd5vLA/r
wLGxdqU4Qyu6ktboJjq98a+T/DuuiKdl4phXsiSfMCy1niac83g6k+0c/LGuP18wPknNyaeAjJG7
Rpeg/NpwM00h0w/igztvymLqTx4FB9GhevUdfthcZfme/VsNx8hK9aSH1zqQvoENT3r94wdxyD4f
dz1Ae4oDNxcTFNbajPR5uouW+JOgjacyxDGdW8Pd2+37RWzT8eIVnQkVT4gltDTFegxNJpd0hMeU
Lel/23fbqI5unMlbwLz/MKYm3gGGKR0vIcl0jFg7MDhZW9Du/yAPeCdMblK7+bcYWO+W8Cqr5q5T
RmDjcBTEIvUla4CBvQewLr2jvKUtiYRJn3JD+0IneSoEPbmLfOo/9yAv/avIlH4etLT7tMHrviVd
JRVTLPSLG4Qb7nYo+51pjxILJkwORjQkinV1tIUPtapQRxgz1vkBfdp63PB10iLBhkalpTl/5vz3
u9FSYsW4uw7Le76i6+4iRk4DwlYzUBe848NPPUHJJf8qQ0vb3Kbg5NRHEUG9fNbmQMSzUHxuWX3q
yR3mtgOkadRibhs5YrlrTBjYJ2dW/3fUJ+bXDjKx6RHaOTRGnEWSgIueDfE9uc3HZRmiwUQUfxSn
BkBj8qRCeGw6tXF+vdq/DN4Zddy8wKTAwau/HTiHSlcImiBzigw9mMeoE1ryHQ2fjZIjnsR1bsNG
xCbEh3C/MtRNWfYGtpgdbjuiZ5KW3u3G6n9skQpxlGB0BCJrqiPYTtC9gl2QVER085ODTGi7gZBn
Bwy0EAXyBT0sE+qj76OueAcW8O81GeEWrRFRDMvxYUJVVM4tUftnPLC3yY0glAMmxGLKPPfmL1pz
B+/F6bRazgegfsFEL2y9v93EFu6NobwChCWQn8P7qknS1NcX+CL+JZxS+zcLeo5euc7qa0Ie4T8t
6g5JTcm0mnprblVGxk/5sqENKzd+5BwVMxJclpOTjuLLmgu/TOSe8bTv4HMl7UswL922qY6z3gDr
yTRkP9NlQbzL+QK4IdRregcVhHZPZs/R1y4gmjF7NgUz2HJ0PcjZ3vekELeKO1B1uNyUoHnqYabY
Zm6CM5DL1/k6n5IuQ4dFPaaVCDzONVk1bTNX5Ql8kqxQwQTvQ5Yk8uVfS5PHyaosV3KABQ3IDf59
QaLsqABpToH8SpSO0JkWYINfoVBXagORg09kYxVTwPbq3x4j+h+CgAANSw1mnzXm90h4/DB9A9Xj
eoY8Wnhdk/jSL+KiHPveekuG1UXXQ9bXWf0ZDcxl6jfvzdNhwgbcJvMGP/qLEGndyj2Lo4f6zPbJ
gQ/x/ryMatH+F1Ls9SDhcVEMAfueYPLuIa6/7PTokbB+kHFw4uP4N7+0Q38mCogoWpVYwSj30E4H
8u1ysE5tlFl5VLEpU/nTzWsRUx07WO205/NqjPD4QFfNrQHFb7YyK8Ru2kuHxAmJmlsJiO0qlOdn
YoQCg+t3rp7BZXaB9GkfN51AuiPNOPRKyuDbn8Pjo87yuTwqa+b378WlZ3eN2qmrMjAC+ozLm4NO
XW3Pl3rh2naFRU3RuIJxD2Pa4GERnCOeW4Bdz5GXptsVmHOBwF1GitqhBOat0yHRvVji3Huuj1F6
cvR7GzTGbJfFVs5rtu1ZGQDk2ISdCYJ5WU+79XlrHkhLx8n2c6ufIX+OXRSfdIN7mZJQZKrTmTAU
YpTgWFj1NZOkieIzJE7BndYRBtAsvJwsbGihXNnWeYt3TmvRdyTOTxtEA9sSo6+ON18CZlb6fnZB
ld3/6GUgq5avdDjSRSAw2y0IlhNgmjZ68tHLhBz6ZcgMhpoyn/gRKg2apGWoDWDcsnUNEn78c4FD
gkfkey3UhMx8EsW+aG+6nxbjsNdo2T9Mbh7K5NHq8gMxr6nj+0KBWej4z2NVvzBg0uApYAi6dMc8
mUaVV0uYrtNPIqCTx0mo8WBuMkC8VyMA6Oydah5TAiR1Svkcllvjt9o5Amp3FwrO4EQOjjC6smKN
cuS197Vwv75quWgrPJklDQ8KhXfhGDeVW9heTVAf+GuYeSlYQRJ4paa3lxgdlDVJOMu8yEu5c4YK
vrze9ZRrdMltlDuHDmZqQlFiGVTTuVyGfOMdyqFLElesfqgw72aDNMm+Syn8xeEGnX8emOE49YZJ
JBuzKLVLGSQqm7/3YqfvPgmuV4fJNR6/+DqRZ3PjqweBnbqB1kE8anhTLntAm8pdDbEf7VDCZbV9
0YQ8xqaTclXjYMpCPJ4YlcCFc5utTFVODa/f+yClpBZhQpskUe2YqjnPm7C0OeoEBMWAcPuIEzIn
vxd2TxFCinZbXuvWsc+XIjQhdIbD9YrHChvV0IjfjMhHnEHMj5BrcDe3tZkCB2HPdu5jpGG/wKSS
LMBKCEFe8BCVK7vQg2nwFbvnAgbV8nwiftJgT/Rmv9CVBONpitHRbWRLoChXYwHl/W9b//Ve4BJF
qjZfw+JNoZU7yrnDRGwRRbkh9U0FLnmNLU9POQkfOi6XrIPbGceC7XzXdzCWjVRQ+qUpbQtPZVdB
fKGSZS4iy1+H3dFuoxE344/UCqikiHCYCj5kCb7cCy8AEVp4HXAqJbOgk3TZQk8auEF6xaztQNNy
5ygGihVtPYc8kMmWH6EFM0Egoi4BBrtitWb47RoaHoHWIF6PmErSnzzE+SYqD19ymXcwfKRY+EvA
Ab5kQtpKBIldF16KPnWtbhbNhA9zF2a1BP88VeLzHkN7lE5eHNN5Zd0FzIgnu3mDR2NUkOjEp0dS
DSYgKPG5Rx9WFvMG9sBD9pA26Q3e3Ohzt4i0rWBQf43YvJ7SUF97erIvULemBZbFK38YlfeBSQS9
iRPV33Pc74ADJ/H0rw8uc8DgQlkzymjATvjiLqQjhCbE9SLuWHavyOf4DRGrFkbrRUp7wOxhrFem
/ZkOep1bdb8SpP3gWw/8BnLyUNQukzo3ICXCMpvMExodnMT79nvmER9KXpR39V3TIBBD0yvcCjDu
NjY0AlP//jb5isELBAsCzDYwZUUVeoHns6olSWvcVfuzkk7w+oBCqZc4+JqPNOEYTGFV1W4r2/9V
gF8lfqzVCjdnU0iBKEhScoNtLf8s2Rcdpxt87ISMXZUtrfl5zB2HE300xXuULlA4I1fZqX32yxHp
wUY8Qs04i5wT1bMm8qOT1+TZA/wTnmhBkuHE5sMf/hpPewvwtBU7p06XpNIbg3UCLtxYVXcclwEY
mLbYFhRWmtL9VoE+dEa94azZDxHxyuwExLkskKmaRFipV9P2l2qj9kXTP19MnnUYBVdWDpepWtrM
ElAPAqH5QOEsmXyuL6iVpQSn1ghCIhLoy3FuCowqffMYtrwgY2KCynwaqiAIrAjLqaphz6GzYGNf
3GPWGwHvuRThaY6oh1oRo6vHm7wcaf5z8XF4a2OhiNtd4FiN7Me7R3yfRf8M7EpNUoJN0TYbv1V0
kAWnfR1zSMHrSxoXAENWbhvGc1yXpchha07eXDTdvxsi1x4wqmp+0lPFbdG5dmNbiALjeU1dXjCP
DKHg8eDm/arQeioB1Hzlta4gnQxT/+tOJVUJUK7sEa8K+QpR3Dv2YBznP3DTRBLJppNrJXOD1X6M
n1Fuv2VDACM8WX5aK52AxKXS2VyNiiLJyP2GV5WcsMQ43CXXpED6GqMlveK0aWutkRiZLtADV04c
z/y8yCstvOpP7L3XTyeeb5DCmOPkV2UGRBRfUAkhsL/ahrzFrIfAZQU+u8TcduOlXSkfqXEjaUaB
mEpj24ZhK8FesfocpFxsxY4s8svtsFyq+keTIj1u5AZ3YuYBijo1AG7z5LOnnTfd3DR4STOgLhX+
BpgPR+IyspKtmi+sr48U+uTPWkomFeL6w9OJKvMF3eRa4ulBoOzFjS71ugDfhlGlBfCZcgdOSVC9
q5cV7dYwiZNHAjDoecPBMEizdabo//HJ8OzSU44//Dypx6nm5/CAgba5FFeJtllr4Gc7MrHog+lr
WeW/JCSaODdQ2Kq6L/ZtBrEssM86ulob+YIjVdNTM8UXgdH0KWXmECagRZ2NhCHBvTbCDatyrMeD
AHHGRBrk0xALkGCL5qkOsdaCTnu/N9JCLyd35ZzaBSm7Lk0YFt+10vQItal9oO+5cBwOKvPy7/Pi
MWib54KyMiHSbIHiZgDp3Qmk2/l7Mb74unHAkSC85F1e5F948sJXmPgvUz41FFxP/fdc78iYVvWA
vc+vbvWviudt4biVbsXeiNXK2uFj667wYxkxmdDYlrQYvSuNreI+kjyj56Bc/B6Asx754kBEg8Fu
nn6SN985yQMaq0891w6DNhOFd3RMuRmHzSC9j29wkUEjjne15UBlJy3BmCi3QsGJdTOAiGUns1KY
pgbrAJcHZQe719iM0PwcVI3kNJiv9CJ1X4uDcHJQ7Cv5x8pzVxh6/5KPtOdiSqF/4RFs7NJyp2mU
lDqZzh3QkVD381DSKyGgPRhxIBVAjPgGhREr77yHPy8fFc4bfcyZQo4sXYhR8zVt/NWNtspzqP3U
kUUUGfkFYOvJ7WpuV5FvcsDOJeoiZkdygSDe5pbWPOQ/IrpLt8aCEG3Kr8zeYgkVNkMlb0x161+6
EgsyMsLEXZgGo79wCF0qdHAQnlMCD3CEQa6EdbSTYIWh+f35TOZ7BxrKyoeAykE+9CjautSOimSw
pVVTq73jLjLsPDjja44Haf3f9TapHXHBcXIhSAE7LdISXR06NrzPC/gwR5kPpH6t2Eo0J31Bdzul
a55pEIDzqswW71cEP6YZLyuQVOjIjZgmdJw4HNrbvPqomMbElYHeuEdn1JJQAcxTkmd9WFGMfI2U
0fpUaVybVAbWk2QOh2EAwTTYTTp6Qi1PmPtwucnRqnH8EgkF2IxKrogKradlcKaRbP4+KZ0cs+WU
fSIIAkQZQ1na7bMgC+ACdNJ5pmxwr3uIvwDuD8sVjvTHpdYofS9B/AriqCrh3XD/+hLWHi498k28
Cd8m/15bsWgfEPeZd7dc5dv/5s8ZROj38qv7ip1PaFzUhgCSovLo0DpPe6dixBfS9HodRegWSvOD
HZJdrFXyYvvtQLqzDdylkyZHY7va0PkwW9KCGG/CX0kZv0EuPYCvd9LLJKUGWet1bvf/sB3xXlON
/5yw0c3Bpe1yNI9+aIrpo6gGBOCP43jwIjqMZyPaifvRQzJoFOVREHlXrnn+/NVZqOoiUU1+He/u
oZ7thWVX4QaGkyAadCuX9bBJvcmyvjY6Vf3b7NA4w6Nob+TJ6pwfqBF7OSXUhk7LYp6Rlkeoy7LN
BESqw7O9gTGAxKlfh2XVWFiCGhy/7lbJ1m+iwqpaU77RFAFouy6NKQVwcR0i6VCfTfhawuwxMt1N
H/L7YphsCy3EdNUmipJcWbn/iKcdRUJNO5Yhk3NP5HnAdKayorwHvVkik0oLm0IwlMDqhv3XR6gs
QpzMye+N2pQivQMN4xS/jQc1nPrXsTabUXOnkKP/hbD/uwJ75qpCF+RoP3b97J2HDntvHVY3DHM3
2kzZIDhyqlyG63Dd+yKO0WTRwJdrSWh/xGaxZ7dAKv16Ju+w0Pg1pZXf14aQ9PrxtT+700JeVImE
dqbQ8xQndGee5NLauEv2sVFAHLa31/UNE0vh8IKf3fwoe/8k7tlgWY/6wYoAYK3YgAhYCoOfbdu8
XqWMnnCsxZIc1ZXtc/cRyl513i8bl+sELz5TUYC57XXwigCvQjP3YR9aK0Y92S/BkWhijHyZ7+fn
Qjze/nKHJmdCHdDkC8hWZucrovqa+nv9+a0DWYONp35QBuO6Kiiga0ewPUXyZcyl8esSwGdlHYTd
e08mbXbYClwnpdiqxSGmZqnCQk/AbhQZgUD8X29zliO3bfburHnlKrH/4uErJroVBH5SkVioLW5b
j5GLCHKB3gvTYn6QnJ8EcquC85pygJY/yt/gK9VyHtSoWpMR8MrmB0onUxW9bbQQLYqU7GOq6QnM
jFj23TUQnbRp8CuM5hJkSGfAia1lCkW0gRKI80dgMYQer3NDp02SeEKN4v7KS1sBUhn+psH9p7Dj
Myi4DtGWnjcjDsyAfbKz/zyyTsFpeEWH5J03g7ajakNArpF02E5/e/AVMg/7nYUW0euJEHGVb5Tr
tZBhao7jnMRtJkDj2WxcqVJpcuT0WJLwBkuOTvMqbBcK3F89XNCnzgdbIRq9KgBN907+2KUKot9S
AymwCvs1I0+whxglbkVTnksJ++bmAO0pYbeQM8vagAFdFIz+RkRBRqrwK5kbYclVt922KBxuQJr3
Z8b0fK5mNXwnKM6t5xybq26e4QIAUoT4kfy2Fh8gNF01u5uBFmC65SmCXjjcTCmecO4xcPUgV1kA
5ZF5u7SMH0mvN4bIuqgnw/1UstveUm6MEnbg6K16u3zKYKu8JD7cxJdM9+vTFvZhvS1y5gN8iHu5
pHf2JI0xRBo7CL7XFqo64i+i6Cx6PfwuPf8NofV6Vu2Qf1XSxLYSiv17sn7JMNqcdBUqlY9aaMdO
OmMbnoPrXT5z6S2Fhx6AScRKbjL5CRZFuozYUUJUmscQDp3hu6hocWOfBwxp3Q/x4+E8wbNH7sVl
HCrf7DcOz/XnoHkst3TKQYXkyM12lcCsL34U41zcaAu7lFccLNuhXHLdWM0av0LhRehjPYCWpOvI
X7L7laX8rFmHRkbMOONRX8PY5nIvjOZ9X9NZfyRWy5d9opsxgW3899B5wCJi90I6vJ3gGL+M2cd+
Vrp6tsD2EQFUZkZqgWsPEp85/2KJh95PZzdlG82Hv+s3u86SbZcpLoEN4UkOJNM19Qaj4gT9Lotn
cKkhHmX3vynvn5FFXlcEI8mQNJ0HlECC/kw3HYajvWqLNSfqSZL6ShYm4Ay3AcpSNYxL0OQJ5P2C
vje1AhYn+vD6+3Lwi9MqMsMkpAayqFW1l+mMGkb9xCag8hyq77tWYjACV9hjuLzbKcF6aYMKbUj5
VjAY4yzt6eFfni0XXcq0qkct/+JdxV1vMPubL/1cu2ZoEv5R5vi5jV1RlaYX56UbYZAfBPjr4u6X
nrzTEqNY14vK1TY5b+HheTRB8ff7DmRA5Hc1hTfQwWurHAwEr9+2haAr1DzcWlQdii6gjbh6pEkH
KB2mWVkiIiZ7FZjmuOQy6YMOi4su5vniHQ8wB4Dkv4BRQpgtpQaFM98Yhl4q8kJmJ7B8FggAS9SE
PdAkshnpUJ2WaWPAjjB7yrDt0EVVJL70X2YwP9r3ZDIQjnNyYqn+FCz8khRX4z7YeOO2JjsGz8dX
PvjEoHSfwof3M2C1cItzRxJSFy6Cgs4Pg8n6GVn5aQJ8uiUJH5G3kbBNyq2HBMHx/39L6cXtoUH+
k4oK+27K9CeO/8gr3Q4n7XmvGxhqS2bAjIcdhTnGYq16IivUj5BeIyZkzBvRX4REiKROgPEjkVfb
ZYOyeZIyAoZOiUB/JDa/LjsqnQgFV/GZJgI0b6TATqiW4F2GoVZb1IUxZdF8dXf7Wtlop/sv9RJd
v9u/8q3wBrEsDTFVosemoUOj6q6GSzjsMBb0ay7/d5rh31pKaD+kiZIN0wyVMQ7PCio+d5Jj/69O
97YKovV2OY1/F0vINgxsZtdwU7+9XRBPvZyHCiJS1e1lcN+6VwEpkSG1lOP4zl2KRukxMzQHQ8/m
sCToIv/SY36L2CJ6hiGuBqQwgJqOwrGIn7PGgq0EVT/aCWQjI+D4rLxDJH5YlWE7qhy/XB/B4Rxx
P+TOwhrgQ8XCXiZBXMRe0b5nYL3X57+dIH9dKayCF8sv1MMW23ONBERW1vBSsUr5cz+SiXp5B8ev
ZTYtJj9LDfqDC9P1TE+VfmnGm9fQJ1Kera/K5WWCJ/285hr2iIHnXkb8NB04GZbr2su4xfcftIl0
iy4W6MODWDY9dkEBW1/Q2I5oR6XVTeIaUM4j3vkOzMPzGl4yy25KCXprtrd7TgJdDHfPZQZVFK3U
+T879Z8SIA04Rpu42a5bh9X2tL4Hb7UUTyTBWPr8vCVk15KuLonYHXAsgnE8tdRxdHQysDa6jG9X
2KYQCvPkQ/oNy9xnCGXzHlB0n860J447Lk9wPj8/5kT8yPT9MA+G+1tlU3FjisqEJS+mhVUY3xz7
neopdopgEfMdJVaqdsr2XwBDn2aj3C28djgXjVyL6wYINOjqRda71irVr8LqCtzzMsFuHa9hmTgN
kU8RrQ7/ZgwcYAxAvN+Jq3I8YXdoedaQ39/jgfuxk/rfQXZZGUGHlKynspLzDlSiGg+mCsHMR7Zh
AtlJgz39Ejv1bFzhlgvX3HRPWf5sCbe7RRbMS483icMXm5GqnaYYHYRFPqpUFZP7mNnUw0hgF11S
hyOoiSvn0sBYMbOu/aZWuOoQIoiVvWfTCjMUieGmOvNFWPGiUKgAJ4JBjseUSEODiTDPEk0+8/bc
U+P09FA8UoThyW0cDc6aUyTw14YTJl11gYw9gN6ZQFi3IwhqU9jCYlDieNhxlhPdYmWlZTVwEYhg
qv1yxyMZAVlwdKKUMyc0VOOdNfBy1NYC3Lsx7lBPzsKVsXbAVnsClxlMi8ZvMpJWwoHOqt1bCAGu
eM6lYOXnvIt/UL8ApSAyrQ/Iwm8Quft+W22VWaQ106ketU973IFxZQUPPTXnMJnHjM8KYuoWhmOd
xNtrndFFLFzcA/OqTWxyQV3Cm+FlHNXC3f0+Hh4WZo0Y9vd1QQWL880HJ/RPziA+iv2zW9wCAaiu
GU6wDSWpKX00b4KAwU14UsEjZXOMquIV1+vf7fC+B/HqHgR7JDQPiXo3ZMIjP/0rNyDJioEfqfrC
mmwgzm7bVYWos+xMIioPveUrsLmO4Gqev5KBr2LMEgSaniCZ/HXNW8knVxHNTRWAqAx+RbYFz07p
OgWpn6BmdpeTcfij0Y/95rLPAL++17GnlN4HHLYnDgNizEM396h4k7NzfcWNr2iDeENOudTk0KOf
/0VYq+pF2gjaqj1rHQmhiznuCgiE5VwBOVHmmuFuPzxybsN+VnC+bIfHwQH3rifUx2cvYl8UVVS9
TtginFCAaou2AbioOPDzXRzs63MULFueHodQBbr9DHIMHQe6o9GomBRiXRDF6LGd5+AZhRatWi4c
fYA4IpqW7HQq+AUSq5/WHDXF3iD88WIHNBHx3FAXNN3AE1a3QQr6zQ5ye5xV72L2EM4HM2kz5FFj
xVWd/XpjHdUMkwJOpIRvq2X9JPZNwWhjaTjIly3GnikcC826ReFeltLCLPUYKnSU2mh/RfXLqrlr
7mnOuPhU5JtbllA7H8lZPt4/mIMn/5iq3h/4MEqDj+o1Yb8sPrkh4LxYcdLPXKyNn/KuiDaaxvBR
k4YyzFdj6mZHe9MJImie2ib8gLDGQgZtyYEYYserMJs8aledjMgtJVuG8lXks9W029ouF5cpsgNz
1OTWg4wxq2KUoiT8mx/aiDazNxL/1Tm1rzUwilRkZLkdOdnotUii+Lf6IYMimBlocDk7vg7vlvm3
Q/oG5u4WGXfZmF9JNxPWZWSpTVRj7uU+2NKO+eXOrKPY+65fe9WgwJ/VXrTmVynZ7Y5R2BjQtWCb
TZEABzWkd2cl+QM6b7X4FtXB87nydOyFA7NPZb2rBswqoPaDZkJqLd13DYuhMty00wPjE4R+S9iV
4xbIeNWf3oZM+Jsgyc4+1eqp+73QFs3jfq1lolSFz3FAbxmtVePV3E0SRwVfttEUETzgBG2MYSkk
x9NzSDsaqyMG1Q+Dj0+c63f7QbUqPc+Klyw0NQihwq8123OGlXhzQsHfd+CXiaCbI/kca9J36y1i
kHZCCxkPVnt/Ze6r6dbwOUZqNSdEv992JHo9SedoqD1eN5KneleO73SXb7Lw8OD4TriFBr3YXY1n
B+JpEfv1qLS2riBXA1KdUrDhTUemiR5VqT9da5ZI2a6AfOyBPVCFBoMIQ8p45Yw8rbP+tx1amd6Y
WcLCzl85H01++ioPAfgxJpj4nwdlF0T60K2N5UvIPlJAwp8ZXUjEKRcfoxpskVnF5hjGv27ZXrzo
Zj7Y0IsKLQa09ABARFy8/2K3DfdATdlRiNBb6LpJMwuMrqDsYLhCe6GktkDKrKhhRbUgueEFy1Yh
hXyXutjV+bXpihnXaIxHk7M0tU/2h/+GqsxBGLaCJVjLRY3Ui1q+4mgyLbkeDy+uOhwUkjhFo7Xo
zmQ1f7U64UwAWErDKdz7Wuzg3iyqKXAmZW5TqFUCr7KQZGHbn8Wcnr2tGfsLsfnzSxKIezlEE/Ep
WaswLV36LNLvYe3y4Zd5R3t2xyo9lO2oVM+4K3JcO/P5vKlPduLlR0XlubPGB4FLJIxhbata4n+b
1kxliTQGjcvA6I+ytfDtD5XW5iamXKN3NkEoZcMbPwFkG0bnoj/Jsiyzf/wBIyeHKC54nfQMiFL9
cerO4Eb5awxEN9NlU5oSHQm5IXJTREZQAyKevYTw/NNKfEalorSAfVRmmmbcs96W2WyEsYm+YlWD
cYpnY4W0r93O6c4iyJp+3EI40kjx8FelvqARosgHxSwP7kYnaz4R757YKmwpQn6kRRisMFyeas1g
T37ib4uC6py/oA/4KKL/aY2RfbcEQ/RlGProbZTAB9E8S5vCy2QTyU20IqTZ7JZW9xoRhUVMeT/J
7zrhnNhc8YviXFVSf4dhz3Ur0Cj83iQgp82ASncxtn4clwLtptl/cyVrLoFyAmBdfiH+ciZ9KmfD
aZSGKaWOVJLoEXeCeC6M8dI4laWpkDBwtBe5tIL/IcuLaiNtDFtULmAjx85lzkaXOU1Mq9pYSw6u
rzUTIRBtfE0jJ96GYB4c6VGtMjlvbYmuMNrgtkAUFtcwGfQ9fgTj+V8ubdiYESwvJ2t48Mf5bW/x
AlEVoanf0qoOLEYsjPPThc4Dv/7B2nn9YHKAnNUbouba2G0WtbZCLZbDIGbCuINoXArSYbrP66Eg
vObFAvG2OmGqYkVZ/bnI85dJUXKVhTyH9YrfyiPDiVvXOqawJ1R2W7u9CCTNdQAcwPMzPT1dxzZ/
WpsVTOP9OrXsFWOyVW5GgpTBf50g7zzJzJwqsPonlal1189mN3HM2ryZrtLygbZH9ewpFEWf7xbR
0qpEGb31ZKYE1oNG/8Xxmk6GFb2O13AALjDmMMx8XtDxvXYYYwi+wltcjjwhbv2Ko5uMgSl/326K
B9m5h1fgFLfTSToGJlABjL66f8S52dyp3RaJK4X37k9K7Fbn7hM8wOr0tlPlM28VIoj44qw5bi7T
dF5V+K5EIfJIQ7jEmy63gRrMaguAkaq5BXkeUXROnbrP8+amyggUVbCHrJkE1fmA8KrRxEQuAp8M
kMN0Zu5BrAcNHtaWe18e54NOtpeKFICghgNainCMCrtFnND8OB3lz6pEB2jD1ZYpAqZQ+5+6ZAAq
ceTKcTjJkL8HjE92VYv2k9pEVYmybgXSeqwXOISv7VbZ/KAa5GcDIb/avbFPrNHnT0qY1I1kNF0m
02quS4Oh/JxhN+QjER5iFGvY3ZZq9wtdki4DoL91/qtBxhw841uCzcCYbW8TpqAeC/yWa45Bf18t
hAsdbhr20HodUYNpwKmtSbp1elP9sIa+2MIP84fUypKtU3ZMhLCGQ0XjVKckYMrUrDIfE+oB+o9D
YpGO+Y3LPKYYKe7x3DF0PkaPU8NoaMTOA0tVaLhSm4i6H1/QLN7GffdOno2D92s+SUvOIV/WaXpI
8hnn1cZWAyVPm+dw9yi/W24I+Fux2rFoixFs4RUNZnWbw+y62UbiXvA6IwJxfThfE/TIyMoZfPTI
NCmtNUNIuzrLHTt17h5FVo4Ma8hmeY0nVaCduvhCJOIwbXCEj0F2ATnKPJI1kaIwS7gOlkFylPIY
7Et8N+qq5RanMahmCtiGznWeH7T4xCvnZA/8grNfBspz5XyNVGPuMrH1EI6jdW1EDkA3eVgNtuNV
btzYWXLF7nxTKcS9SqcgfUDkUphTAjKLhdcM4HUD5zWiHGvvsKLx94qdGjmrlcZfLW1uwARGoNVT
uAVCRVr4w5baqs2fEESQ9N6M9xuI+Nli2AHaXhqltyGf2OroJnc9JaNsBZS7H2KTSSNiqnCxBgtN
kvG2LIHUpXXOA6JBge9SJNH20rMvrwdBJg9nq9NLZWdMrQcHoMAp2N4zfcvYQEuBYGvf4CdIMaBW
ecBrdXuc/sT2dZLLHlUiQvRNh9dWJWNtqur3a7m/OVynlCUg1hlVWLhAmGouz0vwPUE87d0Rtpl6
/8BQf9VBzdm51gDJ/8I3QTMo8aIjkb0XKJFLchZwtzMSsA+tE3Zi7w0H1O/agi4OkOwyo7SqnEyu
qAKcQGLK/rnvROBQ/CjBd6pCLLl+o2c7GFPecyBchqFJ8zUl4Y5RQEQ3eEndP9K7wqzzLsUuxoJ8
g6r3dvnTN91xZn2RquMVSbhwp91oxsK4Ltgcnm6e8+5JGAd0c9DshLa+b7KRSu/zJLCeXZARVtp3
70s+oxq+Tf8m3JQKmHvjoaoBjQNrFFhjjRouNNglQl8EUrecNetAQpgoE9/TEsUFbr3yxaLDEvSW
Y0XWuJQYKk1hEmka9UDv1SCVsG38kY8y8YcX5Km4IqcU18kRX/jC9hwZCoJl8m9jjoankwZMorgn
L7BohNHe1hnSjKMJXHN/8qcVFA4ERejGWFUtBGeqrdxDLZAv+c2OpsPZBFFgJmea89d22heKrlKx
/lTK7/YQgZFdRb7W1vB28S+sa0a2lHqgeGYv7iyDnjfedXCgv9iWxfBJDtyxLSEEDh8tl02bKkaJ
OCYXXswoP8pj66RLmA/1FoZIHAe5CIcpnCYUOYaoMpiswcDbiJnPOyOl7m6gcUY99UPqSGXqQ/2c
kgfgJ9YC5/LPhjQEwXkbG7fEmNpD2PIt2lVp+N8oyYWlvOlgL+46zVnExgz3En808BcM1UuRijsM
nghardW870gXsKpFzhLEAR6R3d2wH2p6HbCRyKd5FHqu4zIrn/iIQjdmTSzoM4vDFyDgaOkBdzOF
8fPMLLcGoYtvnkQgECiCiHk04YMBsuJBgvG1An81PiY055TeycXDVXxEheZaU/tFOcTmgjKntycd
IRdd3/baUtZDCQUNu46A6c6QHte9KVwYryvkxPwWsKMe7KlBEgt58No8vhSfiljT1KEmY3L1+8ek
ycCq4MosxTV3PUy8s0XgHH5eT8iXnJuWKnxxnnw1M5FusY9zjMS1uyul+M3o4XyF1Vrxqb5qcY1e
UnwtekLjHrmXxvjknMKoW3J2PuR5oRsX3YYsX+/abBQTOIA84/uReZrshdspYUEi86S4N9dcuuV3
kEaW11AIe3fsBM7LIyrQWrxX2rgnSL9Bl0kYAnxuzsfwSpe+YSCdyEpIU7LVBC/IgTGLV84sGyZI
k7gIHFhy7M1LAeT0n/sGXf8Ep4ZhTCDNABn9+8NSByvgfWlGOzI+IyLuIQORtSe3y3rs7d+IYqKG
+tcyPdzwp1eX9TQZ41TV0dysfJNNwtmcNciEUSk0ks+DnQls9Y4vZ5SYC+g0bsUODM4QUBJ7NQcm
P4zAyIDNhDlXIcDOPDtB6p2Kp0Zcs2n80vyum21iVyEIKG6VuopCdBT2+mFeGTvA3jQ5ctingie5
Rxf8Bh1RJGd71F/BtKIe8TBfjewggrVFDK13H0LiPiTQgje5WWWwMt6En6oXeM4DW3fWJG77JwJV
WKnD8Uz2yc+1/vdp+obYM/2VjCsx6zTqgNmIXp3z0CGiFwcS+sdC6F2wqFOWj4tRGlGr729gEt2H
otb61a50mMZxYe8TR9x9xae7NRHMwqHfdQO77jgrqYjdbIay5scTcJz5Z5no46O8aBGDGtOON2SC
sAEHrIdQduFoeqduo+TiGMEo54XqUknkPUyqMEmxp0GkAWIRe604iofl90s55amnWhsOK3OSNW57
RHiuOgTt22C2AXj8/KazLoEcICFYAdl2aYvcn9ZqgPJTBh4Wt8zhBUXpK61Jcn4PRk0xnK5wDdP/
4uFvF6BmYyAEbHm/xQ0gLSGAKrMPuLn1Zb1ETFFRh3PUtmHfMC+qRSKvLQ1a09UWwgsQf6a87ssY
kJr1ZaLVodoInSFKREC1UYm0owQTX0OYwlWgmNICfJU6zP9QdPph0D+U/wH+tUqEqKbZMGsXRhSr
euu2m12Y/WP1iwHymx+zx5065cIzg9Gyl9Fx/FvjHWzyTf5Due5eCE3gaSlrB/L5eW90G2g3SBqw
mmWcAiyU5Arn5e0GK7/MlpWcUrnzl35TuYjOPihPeRA4zoYHuOWBnXZmVRES/a+TGTITJpPI+pK7
CgUbYMtea3NhgJijHopVA4rD4sAPNYs8KPwgxx0LlCWZnrh+6JRz8pR02dZs/YfSxRu7o+9yKP2Z
Gf7PH/B2/UYrv4zbLEecVReNmLBpjp0Z+RIe9YRzuccqWW9gKvXcJOybbPugm82Oe0PVfABIdqoy
ho3H6C9K6nOKvzHyQEWvV/JlWu9ZSH3Xx3HIQY83OKICVyJIxMLvh3RbkuhaL6yffpEXdc+g5OO3
wQmWzl4HLSktQmJIx7cWtgfRXn8XzEX4g1GqkRyv052uG2iehooi2o4+LikvqSBa/3tOtEXnE8B9
uZ/htZ+T+On7JtQFOc+szIw5uOrSzk3JMgqhNNJJKQOQNoE8fFCIs9vGzLsl0ynNaMhuQWTVGI/6
71KYdsN0jnBEpQMudlZ5tSZxf4xn8SvAq3mo9MQxF7GsfqNgCyQYU8A2z9ZSwSsfTcB1iPJmDwQM
KO9K/ScHxm47M5BGOzg8KgJOSUG33m/OamoL6dqkHW44TaOvhZLDD3QRV7AYZQpbD6zxXQHAhcse
kyukuh0/vEm8wzrq/nlx/TDiHgoH68qRWyjC4YCKGstDi2+5wQFElfsAcZShYvpsOHQ+01P2BoMJ
6JdJO8pHW5pLq2sHhmOKuBF9+Gr/l36k0tdq5m8wtersGOVhYpz7Uk/Xve9QRumRs8z576/MklBF
HKPtu36Baso9sHd03YHI5A8To26V1WkaGU4zy0Y9OqGBefSmN93/9NglUdoh+B/AcYonDHXG0sxT
9cFAwRpLL4jmUa3brw7Bs/ZZbpb6ao7CmWyef70hRR97tfj6NcOFUl5MXVJOC23jkogWvDRi+QrN
46v+xd0ATx0YXgNM2AqlS8H/1cAePI51FMkMvog0i/ziFErhCnsiEewTTx5pWKYU6v55BAEFAxbQ
JFVXOIfLKpgw1B3obZsAYpXNrazunBtuaG1pRe2K0hg3ZWCJ7mQInfq8EpMl+AhIIAi6+YIjtdgM
F2jdjam9nezQ2L6PaGqvGqk0hFZrt2/VO56ZXh2ie3C063V5RjiGsOGOPoeJ8FJeci6xZj9FIPni
3efYgTCjkRoSLFxvY0SojwyYlg85yKrAe2X0f+GpSlT/a++yAnfhH+CjzXqDP5hDj0cOT6PTk9oW
O6m0KdLXzgbNa8+31W0rIsg8A1102o0g+t9Q6osr1XV7ahfGqKJ6n2Hb4O7dABLVclBWhPQA6yUj
hFL6yeonTG5ArKeIU4mi2woWLREChdruEjDw7slZsHar2BxYIJlvRML104h7L2o4Tq+uKTscEvn1
01tpfMYMkdLgS7R4HpwdzJTo433OyrzQM9mNv+K7M/Q2x9RBPnFoZZjvEzrxgOULWkRjzfVLrg0I
C5SmIhsGkELFy4GPAfsoOZZAjRKp4wdPMxeEhzM3RAeyef+UXjxyrgw34bGVVXDLA300wk4Cm9+V
99ffS4h0CHBMd826DcRRVWWrnaGwHEgAQx6SbUh4KolmrprIMdg0C1cT4khUz9fUTZUlkV/9nFgf
+4votP6GDg1Oc3kZ4FYB9MAIlN8qds+U2Z5fsrNatRerp9AseRFtq+PyZWPhu0a5pHhAoIZKswD0
flWraETQj6HwxORdwn9pq19mAduHbu8tafzW+0P6O6UevboJbLrYdC3VljwxHI54+xb0dAOokjRD
V30Ek6faKBnXlxxrr5bTER3LEr9KD4/4i+XgpGg+1jiRX2UAYqt7M5+ARDsrvYWEKpgU9uaxCcD9
FymwCyFiAMoUdtMdbxn47T27CFImNQ6Ix1bzK+WEvS2nL0pTqGspK8IDL3fLDUd9C39hBFDAisw9
WhmgXYbsHWE68ozVOeO9kMuNXclDqWTNy/hjlsp3yvktdc4/Tca1PBUue+x8Dl0lyzBoibxCwkZm
Pqrm/xk+jtjoGzHjE1/JOrRTqlx2e0sKGfqiv0PKLXM+dPARij5vbUsnMU02iK23YOfJj55HT43U
lvpouCF89PTLoI+wU2KXiBPp/70oXJFMBCDCtx8Tzg8uFkX3z5UqmMaZx8aTQ/ldQYt8XJD4nvI7
Fk4b1xlSADKCxLi4waRbXaK2dDe4bNzOYoRHS2ht0a8xOot0TMm4bKuc03wCB+FJGKAxwRg7OVFb
56dTfDHcLRZ1pBBCnwCxNw390zSXxjTurABqPvxwgo9ymr1oDEXIezOjxJQDe3YPQxr2wwBZhsjY
jHYDZ14fG7qHuXRzt0rKdRpRyC8XHOs+VqXwf2EZX7cy+R7XA0V536/f5bzaqjyhB570iOGN11OL
P+l5BMPwrH+M3+nzNP+v8LM6Y5EawlQtFma2SUMUxXU1O6wERqNjHvUoYP+aYbKIiuk1TH94Ngc4
WO9nftYAnGbG4SbrnCmZlO5hiS2D0lqbTxlqfpjr/qKe5nCMe6W7etL16gBANOSdlCLUPgiPkTgz
u3HLAyr0Q74Pg43NmsoMl0XsciZ+42aKSIETochUZIcehDCrGbZ2pr8aESX/6eoQXXiKSNS6PbLX
lq2cS5k4vcc36swxSMz9QfcUkCzDdPFzgOcM2uEN9VfX5HyZ6soIGEIpv+I6hX2WFqvZPTxx3nGQ
9Nd7ZRqLidW49OYprO0/2t2ivezwT+Cq0TneYuH3e+u6yiQCrxBHdfa5T2DfaeUDCTXGCD3ZNRc0
8aG4pvERm4zLT8cENKCoPwv+MLkDJmkH4wK2P4mxcbVkR2vu2raP0TSS4CRKWwaUcq8tivsnsN6b
7xrmj24uziQCiHbM8d9OZOj7yZ+aY8bfq+K4Vz5q2go3x5b6vgLIpBMuEbrjGpN8gMXjw9rxZkyI
dN4SIPKMzdy38OeZHJOEAcu6FTq91MeUiOzOrfdlXcXC9hp3C9j6EAWs+8/YwFFZc7mN8j/Xeni/
y4F39qjh85JzgO/PD7JnMzCPYp2JydDjI8M0/0espbcAv45dkGZIc4y/NXWp7NgWIvHSSXG4ds+O
NS1gU0keObN0W0tnF5jXxADA8SlSfyq8aCwQRrij+kJgCeQEJZDnCKMDi7E0BrfvG8ZUgcvuETUI
fmKLRh24gweMo5AfjGh31eZidRKN6reHhPxJf8NzA7JKYUjdGTdJv+tNBb1sYiCB+EJK8HkWuN+Z
7APxC0f1QCgE9SquF3Mb1hmsnXLRKO0oNKTYUHkey3omRKQBPmfFJ0tEuyWZNWdfx2L0AHJJrE4k
gziGarmHbVynU87rqQVEIUBZymHAioIPLbKydQnC4v7VJzsuSUat0CqTiXm3bC65kW52NWlHRhL4
MopxnHrAQNYvY23ttkvWAyUwsijETqL7rr69kfjOUypOInoBQTWkc4nqRAKei2hneEfTrGAntspA
O5Wt3RIulHemFXSvjKCxhpsH6bnBpr6jLkCr5wnEIVCbA4sToLRpvduoz8Tfrg/NiIGQTe89vpmv
XTTvODaEZAuef3osYOGJzgTyZ7SA6xC1g1Kb2SQu5KFpFltHsSw/fsA8miX8PVyqBGb79oknAmX9
x0RzA/kZ2EhK/YcfqmRf5FVzKq6JMuR2Wr1wsAA32xQNy6PSnh11f8tuH7DrSfpR5JMS5Ax70nMZ
E5LXBEkQAfcBIayKvGLhD3oN1sP68kos8v+8SRebrXfri1n6TPHKp/CZ+cio+HgoXdugVjO695BE
gVDOv5/awb5i8HbJ0rphRLLXyM+C0416rrbWSw/7gVM8R6a8sZsE7EWgP8sr/n5Ek1gttJmzzI9w
XqVShUs1b/9B1mhdXe0weL4o4skPTfdpLEoMZSfApLhpG4OQS9+XZwEyVdeh96BW+bZwQZtpLIfm
fs2qrlCBFjuReeVSbwYMiNuy2+i4bVOzjikmVE+PTYoL8V8dCdA6mVz3T8dYVepiioQuZxEse43d
sTr6KvmGtm8ScVRyVj8R9EO8UsvabWTCBPul82Xeo10kQbFFOGe8lKfNHl2DBE8x1C6fh1+f9mbY
yz60x921pQAYnvrc2FCzGUWi+xxVydcnpu/RXmIlm+GqWMluX5eiZEGC2k58/iDIvcszztIHMGLR
kgSpJP4RoAKcK4dgw3aMA/yonyPp2WyOzDM61+sFV/GTqzL7WWEKJbZqyNKeDvP5z5fS0qxO86KC
ciyIaFVhVfDIPbpE6Ve+BrPDbwWkHx4/2pckmaoAMwQaSdS8a1rpkyx1Pc1zc/aQZmyBVe5yoHiw
JS2HqZpTW8lKYdyheY8wstLkZDw2pImtWCFnYLTPD4YeJYfJXpgr5cc89ShIINLDPLwmZUQ4Hw72
yqW4rEt5zsstnMDGCCxDii1gSlqNU3I4O0VtbVGgGlhRJryWwMmDFWmrKBXLA77uMuPcG52ZHM6s
FF5kitrtSnAPpVRNBemElU5A0SLEcUysM/ojojOzU7PbFz70o+uI00CFUKsNzkY0ZsGiYfDhHenN
VuRznl2AmLXPqQXjMk11vI5XffoawxjVfCVzfW8DyslgyvZ9MxeHjd4buSAaY+DpXR0HlsVgf0N8
aq8VALUL9JGyCGWh8o1OaS1Mb8gSOZbeVbgDoAFscJJpxt6QIDlmjx9uJnY7L5EvVfvgtmp4aasZ
Ddv854vyAHnfFH/YuGBt+2vCl6kreGvgdiMakwzZvpNKvRQ9KS/gP2dYHzZJIjcsVg842+0t6rJo
J8+bVMtCAhfDwieV96WTZC9dm5DP5+jAFREnr+ERj9CXXM7W6iQNo3NOFEonAMyoQ89tUYQRfA6q
VV5EQ9CbphWrDLzGO21yGU0bcfzqVKde89QZjS4VCF/Rob+hWD/GgPZ5rKtG9qKlzdGf/pN4/QjH
5xgnYYJaaQc9gLb85pa1I+azPKKgTDiEf3xjhj2o8ir6zhKMQBA7HIRUgheJJyR9C9uragoAu+hz
dnMYYszFTF2Qv37jHkVr0IE0D7Dd5ZuRwD/dhCWSB2GWRByhJrEyZMzN44AAD6B0sbsZ5xNw+r3c
qERYEiqVMG4X/zRNcPzKCtNePKZ0QtjCkQ7F96hoBZNxwenIxJo5YBdgNsT9VbPSR27V+sNyV+7v
l3N2XRmejsnRvCAX0HpuTdjeiUqOGihNUiN2NYiUMIam2PIIhOkwTcPxQiJaKHE72F2JhiQW3z3g
15oMkF4K6u8xpDSjcL5JG5r3FLHiuMqBIdrY76VhZLh4IXQA5U/RZd0I9cM8cmK39n25lJb4l0Ls
p3LcNMzOgN7X6H2SL7G0A9dwSuB9sjtbabatlQMHLnxu+qN6rqrXCdogXR0cglS3SciECt2p8Ano
u4EtDeZBm4v975z1Z05x6FXvg4ChlfJzQr0apj7ndW7LRWN+elUNAH8nBDLYL53P+fovpdCCrnu4
Z1Dk1qkZ6gpECXbcUPRJZ+FP1r1C4rkbglcuE2WX4uWLw4jpZ2IRGP3U30mJEj4OV57RPUPyEk8n
hJQBj36lZLLf8LHf888gWMSdpI7T8mG6zYqu3BHqvjluyVXFwYb5JV2JeFnlWERAzpl2RnmKG6eU
cI1BWRzw8hMOgw6gW9SEmnEy9YK7iugpxqQ227NH9ojmBePTdUeKu9Z1EOsPjDGJVUolHFW+Ll0x
t0aEaFZJ4fdq0dsN8c1RHN53USJEqTnB15dwFinzdSktjoDq9oeFX3JmysR8VHJ1+dgnoq53ArA4
7l+6MrNLl+DwLLfdTSQHoJ1ijuEBK+w2AGN1QU3mJMURgnjId8b5kNmQX/VnO4CeUe8di/56qEs2
mFD+DlGiOI3E3ZsGy07iDICFjF61o5gx4qU7UvsI/9yckLrnoBUJ9O6+PHZmzGRVmcm0KTUofB4F
72t9P538zFS1NwbAVDDNXXCsi84pzgPBzjAMAKqcL+5hTFhrNokin+hS7m79JjAeiSlYyVjLxe3i
Bg6VCZfA1NkQgy5XePQxeDHH619cHJck58Y9uDxNgXTb8O090tY+rgXNktXHHffL0V9fiijmSxxM
+lSHrCGO6dofsXs+t2jmOpAes8rwJYM+NCdHLAyGxNQojtmFbRQhljiIpPdy7cpXclccc4Iq4O31
muJdYUpl+Zp089vRMIU5EnepvpdHdZ8UlBaJ4It1eC54G3GY1NfZKkgRAUGOBjF3o3bqw7WYEmb3
SQBi9GDE1sph+kZPRIhR60PC9NP3Lv273Q5D+MyHpE8UAuokdmDMJqjV1UVWQWmTm1JEN8gDyqAS
sMnCg4PhzMOYEhhs7eKoi8feVwEM3nto2KaePB5T7nGpZZk6RDKIZZYTptWtqMZN0rwdhunU/pYi
lMvaOlKOiT0EhktBHnCCYD29ocWh4VWJFgF9G5P+dBKFtaZN8BDBDXazoerA9K5nFuJSaQz66TBP
6mxLlmAx/07X8YUl6xPJDuWv7POmcbMC+BlWpcxdIoWSaJ1+uIMpNyewRBoHIJEQF8hcEDsIUGLX
jrPpuqwwJgQxIeRJ/zoNY8lZ0clwyrku31FiPfvdJQ+g9ktL3U98K1+Ddxm26tSi5KkbEVl0uBiO
yv11RLop54Vo1JBN4Arvx0MuxNYVBRqVTjIj16CZHA8dyib3AkGyo6Z7NIjZimHRnO/AA3vK7U6c
ieJpUcHa6hUqrpBNpY9h13Tq7+9RIhejlVLvAYHTiEyPlqJTDu3MGNUqhEj6kq0LZ7LpXHvUcmcK
yFCVeu67t+bgW1GYNhEhzeHnERnpgWTVPjVRQ7dYyKIgg48RtUO8FaWTHATxztQ9msieG0pNVGnW
0XWIlfu5wvwaAa00IzypMiviSbVk8aDaPmtZZmE/GcW4Y5yOnluoq0rz1LDH+sHuR+1fz8T54XD5
Y3U0/rf1MzvdxAuHCMqeMNmOj50QEwCo62h548k9AQA7KT5e5dE6ED4tkisJDAsrcc/aj9X6p2U/
mk4L127BpZXecvDAmvJbp/gT9ryNO5iJyKPBf+OhwF+CkAVvviYAe2IQC4iZT9dK3nLPYBe0c9V9
mILROpnSav594W1g6pywL0EFR1hZbKciLOfVoDYnxJGmiShewT/GbDTrkE/UoAePlDs44wEJ46Hm
C64AryzZpNhh7RaADLTSbly1bvXCDUJSeOI0/RpFu2uxVz7tdeqquBIWnBXMc38HWPaWm9hMKSUW
IpSNGluq1HET5PxEf4gmutlp+3WL4zhbDrqXdzylTZWc1pJ3tnfyfwSkyhS0ASF6NYSfP9OLCcLk
m+5Jit10aF0h9/ccu3VtDyd1+ii0jibzUJUmAoZO9Zqk3MpptzqWc8F8XzkktG7xWXTvSlBI4JQc
3n61ocUd91GnUh4svAUCpxgt32TG4mOcRBF8CdO8mRhmNY1VrdqT1Tla2igpD5JPFiX3tOqlLXW+
gNiCV3vlm7pQIrFpey+bW1wUhkicqjjgI4xL01M1/vdcjL8vzXfyro7kx2Zvc5PP03whS0lYaEQE
YW7BVibhx0xle7pxsq9BJaWFIP8WqCPQYVgfzAy9KOmfnu9bR9X9hp22XPBC6ks181CnfQSb8tRm
939JLLB47Q5l0IZWKuCtIUog2lUiWHKpWvMmjaaLM/vDkjj5hhImQjr8jCsltjoz0NfZbu2mrn3E
Jpd9p6yQR74KSSeD0N9cbQIbw7qk/OXO7TFzCr0zrwbJWmzFivpvbpVV/T9qmRa0JJ23KiD3kcjr
vPFq716Sfwm+lEw2yyhNEdHC/DBIX95Hbxij4hBcvBBhz08Rz77MbJBwvcSRFSIFoHmvEO64IttZ
m/34mnLDqLUyXNa2BKw8pIPJM2vucbOBueSfti+NfCzezclgRKt/9QhgYy4WeSBJdh3Gl0q3xH2X
IukDuY9PZzuhkdsq/jS05uMMTTNm7OvzT6HfZiMm1E3N3n7TbXZ35ZIRIxTVw72zBnpPoHou8DK6
AUOxkYP6uMrVCBnGTPHSdbTPm5lgiWpyCEEXPioNeV6Gd8hFbLJFcSmxZ2PsdwQTYB6kOsfTMjS3
JI0K801ziOMSou1QWIDucSuyvYgfW4bhm+H01padFw+WpN+sfZhXddOG7veQ/omL9++5LitsTvEm
uss9GXzbIDrKWRDx+whJh+/JU1HuJa2Kp8aGAVfsFZpG/Ev5zgvNtbst30ergZfrYPBu1xH4h7GF
tC1fty05UQSiHwihH4CgvWvVH5NsawZ5c5Q8iQoOyQalU+3TkY+c1fSQUqSeJIHpuOAAx5mo/EJO
msIjXtR4RHpH6rEhvtCmCxt2MfehT7m3smq1b4HhjwnsODef2YLk0ai0bLQIaUwDBlWOaTZ9pJYC
bh7Q3rPFrmGvXOlqW9MULOeVOycKaW4Z/o8AX1ko6oxTguwsqJDhZfvO6gcw0/rTDZPZrdQnmzNk
RHTihjxGSaNwxtGkVwHhrcSt1DqYx4OIVasN3iFYRsB1Jeci8f8313DFDnAXbsX7BcazSBfXP/tJ
IarSUqXxkQR0JAEBf4xqgX2fzuPtTb7mBkyRTZBCnUTHOonuro+vm0eTqs05s7IJHMgGVyShPhUu
cVXzjQwfFL/ABDY8Thd8Iw4OWa2fmYijQVQ3Afq2nYmymudMykis0MwgVjd0dNJ+O0jTRcRESKo0
DGyoe7GTkgHJ/mCb8YuKfZ7Mdr73JU5ThyVE27P0pXv4mi+hx4lr6q0I2LkOq65YJD5Hr3E4Ai0l
leQgMcsSo0FLJg71uu4KsogNhsIitXrBARJ++kcZS/3Xtk5LzYEH6mY6oxdPNZelQiFZeU/hAx35
INLnLsjP+Tn0cYJgQFQuiOt6VcwVgG82ZwVbtpsD2kNzVcvRSWM5CYMVZ8JvdzAtrqZhTHGS5Pz6
tQbIqw7kVWwuCqS86C58OztgJQ9+9EdSSMdycEYevjGdHjwE+904yXZ1Pv/JY1QRfBjpFAB0NMux
TvOW4QWjNVP6iX7gDV0t676rVJ/CTz+olt/zI9gYdVZW6mfst309NphQFzNBI6CI3saeIBhG8qCM
9+I4/LS/IYJjgbbh2liDfcNcPHEWY2YGWon+z3lLWSeN/tMECLRWB+znqBAquQqWXL+TKNNQvNJ5
vyGmsDbK2quyNBkxWx5OWZFId7j6oav56oDiqIMN0MBc0VQWXs+XhB9rpT5Ffd7zUqbukchZ/N4C
lFFQ1b1BWhlVJil/Ch3MY0DqvTziadEBHFp7egooifzZ2XctwstxmDcZr6Yix5djpvwYyqGg9BEd
WtZ1BdVi0Ob5udZn3acmgc39f86AktMrTRMDN2cFvVhFO+avs2MG4bN+bR2i8MIUSsXaoKCSAiKJ
UyDAwgshVCocKgf/JQ/zUASs5v0oYGOyrbUb0ddB5p8Wo61Cz8xEBHnGsBhXlfF6kHq/8JFOf3U9
6+Z80FdrrAFvaOM3YDC9he6toKOnxroTsgT5EiNV7mXhDDTBpk+slbyWCKnwhCDKKQq9P9yYGARC
MwVvWcc8N5MyXUSCxypwjPfVNO4VCSCz+IvFlBU1uHXzeMcvaq/p/HxwGkCK0Nco2i2qKwHwUYD5
qe2G+/RHR8pvDo85UA1GtaiyaXBgU26V4fHTu/8gF6rg6g8wBGom6OCzfyAOjGsWaHBCy/j3VqNU
IyLQwJ4Efn2zeYVh9uSvBxvUyV99RM+fl6p07inbj+kKcAnAAtlAfxbT9OHNWsZN5f9hEBtxAGR2
BHvb7TOpdQ82LNmRdhWVmn11KZDEsoMosLVcbgR1WLVsZixCLyQKfsnktifprA+lokpYUh/ab3P8
wc3KlkqG2Mx7UnmHJ+KIxKrNQQXp2GzYzJSargkmrEtGmvnhEgRhsThoOwHtt+w1OhCnxjJ+xfD9
Ui8mS+j1sOrCmCATQ2B7HrbQLcH+2hu06zHRbWXEz0wQdhekAnq2rMSo2v9QJaJHoAAT6zHZ6auh
iDBSp3AXWXSE0tfqOJuEhFIkPqRdyMuVrrvfELvKLLL8/cvpSiKnyefcxiZP3l0cGzxVlf45axzs
Aneov0ZJ24izvRSoDmDgFT36Wb8AKR8QGYHWgXCs/WPuTVvc83I/PHPuO+YoE2N797C/VnKfWRss
qMfdhxVkGctm4un/VhLvW0UoP3mts3iQYdbl98WA5SR8a34qVPal5JRS1AEDN1dOiBhcp+D5wjfP
lamG9LPHAuw1urQyf8Anp4pYi/7Iyz6kJWmrUFvE421urrGmjcsi+JeMvKELXnciE8ww88Qsp6O3
wv0oQT1v7n5DedXSOMIrqvbvsOkgFzKkZ8UjvPB+84wP9ZLQSZTf2qWs2wXoZyLb32YHdmh7rbUF
Mjjt+aeZhv8dWviFumgyorcM427zx25epUXm281aHb7whT0As//KY2ZH1Mz7+Yf8D/j/lWGAs2mN
7siq8SDB0t8h+gTJJZKTIzy0L3vBql0pX3DbLjvwXQgWsMGs1qy3x4HTsPxBf02rmO7yBe9DYGDF
dg5hjqKjEzrZFRqa9Q8Gi08F1DiQVBypptQP4nWjWJEBPFjb/K4xe6f17k81ut7C/HNqznOkIq7J
nJXUnKr2DyCbgKq2TZ8LCzM376sVZWuQ7A5uxJUsZQRyyCZmOTnVcH3RS9XHAIr6WxIpcRyS8fjw
PBvoZHmNAy1D79SQHLYFsZaB0PTHII22dxAvNChhe4zxGO7TWBBLltAAQzs3GTThHvOJA+XavA2H
b9nNIBiA1isrliBVd+KtZDB8dQsCwlwlufZZQ40rtuTOvgs6Z4WXbJtb58D65fQ1/NE5h3XEFD5z
+gwRxeIfiYRJNP94M+17U/imtpurMRbp4jE5Aq/hqBYLh77aFiWw+UyE6othVGvHtzdByFYjdjIY
pVi32eaI3gSxaSBg5VZFS3dIvh1souYQB5QzDIA7zSKS9uqsQG8LXDy6n7+bZe+jLsAmyEGssZST
gmLjNzSYgA8OG/V85106rEGQrviFrL5Kjqi9QM+ywLu0v+S06MaRpn5iTS6Iz1Z6aiw9O/OwUKcu
9FJbXq3q/DOUSu1dmt6Ik/fSrdxpPPw2KTYMfaLIUIUHRvu0Ifm53QmItlq4gTUp6LMVMFWxyMZq
+lhfEduTApktMu4JTXHJPfCviq3OrWADy3/XtdEonsScdfVCFUrASpu1dgBXXM9BZrmQFJ9sdL06
kx3Q0hy41m8MTAhGJVXdJL6RhUkcBJPYd1jnTJeSDFf5Sa1a0c+FARFfB6AMhYkZrV5kUvZ5hr1s
/KCkx6lWNWBwJgjpzrsD+7agSJXpzYUDvRWnoigMQdP/rk7RiyoiB8StmNxFl3zsVBxFI/id+yQj
BkcDqfo/blenqMdyqB14z5NH2AAY1yPOsNcasYm+IORlhJcya7DCD+v2Yvd8SKfNDa4eLiqtOjeq
Kpot8lCzd5iV4wegDxNx2EFisF9wG1a6G8Ovc80VnGB0QSd4oL3Aui/ipTZNw0dtrLXVHo4RUO5P
lXKrIRVCBuglA8wpCKfStkp3hGlQ28jTqC8869tntbJmClB80muzgXEBa4KGsgCEu/UkH2cHBgjN
zCiop4AaRa6FewUT2PrtE//7w4yb5zDBCQatPuHPkjC3cYjNcJ2vTioFxx/tovYfY9QNeMUpfhTh
baMzXUc3iDnnsapP6ol2Mntzlo6y2UaHyjUwLwmn29JbS4dVuy7IznH9PxW/UrDb2m7+Cc/Q0Jip
HFOgO4IvFsHleTP6wwCIOFezpCDu+O6BHKkUpwBYiusqSL6nMMmDJhDwDNM52Cng6YZqSF4H55I9
6saAvl4/2kr/Cz8YlwEYmhk2docu+hkP+AEbfqXxkuHUKtsKxEPAcnRR0878WsZq7TpEI0Lq8g1Q
Rb5XvwQd4+Xwc/09GL8srdXVg7tcLyHUJUFjsD+MQda+RMtaERHgzNrqfHggfxfShl0pMg9BxYD3
BE1CPm0gwtRoro2PZvHFE43aFAyGPLE5elvTpItHdwKxhy+DWd7U5V9EsA+auJbTwccBglFbpC+g
VW+BnHVAN9z/vEup7ac5TmX3cUvPhHBm7A5Otax14KrTemZqPLOroBES8kwFaCv6dyCKFBGPtwpO
QvhOQOqHndCQkf97c28MCP2ELHIPK5r8setqf0nBu9lX1gAhFf5FdV7qwSOdkUhGu0nnMsNBzDlY
kTEYyjLMHcHIeqrqzLKCwCrZBRFwmfxUgyXArCq72wnZJ6lSXQ8OGjgjckI/3wPl81F+fB3Hv3hi
u+awk3EsUu401UL6+rNG/HrJe51imMOfxRPNGqmECtnqbZDABgqFpre6SVE9QTO+/yufRDwTqyZv
06S8L7tCu/UOiaW7kA7HrA89LB+PGWdcw872mr5oK/rPqwC0NF8V0ICJReNGIiYT5XGNK7yV+5HJ
V/eJm06k7zKZxnv38PIwe0/33wd8XM8TKnspxK/TiGsmKPcsKodnleWIKfIYFRUOa+DfXxLGOwka
I91ahhlynp7Y7zaKYw1KbPT34pWAA1NKbsK7tkwq0JGST67GPHssLrjphVPPZRjfj/fXcih6wnyd
RIKddrrxW8TrlI/L/33RkzdeGQBMiOgy1aLyb2+1XHo68mD46JAPxYBApq22chBHScA7E0IQE7Co
57QMgDUsVC7qEb0WYWZwVwlUY5u/v66tlESFGPZuLHlfVgrW332z/ZDOQNBfmTDm4fHcb4B/3iVt
0pL0nF9wO2WsmLC3bOKUuRPZ1cfkskLEer5XJEDrWtzznSEIH+1qCYoAtU16ZaeDAlO3XfLCuahM
Gvofs/I5nMuL4LXc40bMQcwi2m+17YLfF23VkN7pP7Gq4RWQMHM0iQL7SOJ0hRYH/OgtPBIao1an
8Wa85xtW4xvMaZGp6d5i+13fO33hQ9TYW+sSyEO8tO9a3YeVfSCO/zxZNPq3p5Hg3IQmfiAmGacH
yuEEZ9QQEYd5RYn7SQKFoSxKbdVEPnYZB/6QpR/lkFSin4IVD7j4/DkdRVojB1mMyffmZMP0Mdxi
Sx3kfUeTGvVdmNMX+r7oD3c6prAJhoGjz1VkrJniLnrzGaaDJ6/kkXvhalmL5EF3f6X0P7Gqn920
dVdh6tnIqyZwHQTViadxcrQmAGp1y2rnELZwes5Srodv7ZD7hRaBjwbKPjixed94054XxpUYCiuR
71WM8G82eHcLjm44bDlLFvWhpId4kD0GPOlR5c4H50liPRNR3DPohsQWbzcCHQJygqrvSwKSB6zA
xMrEAi5dfmJTNIHsyPAs1bvcmbc8q5E3fsAKcaRViiD7uIaQ/mfIce0px8OdJ6gG9aWYpXptlNRr
MylEFqDhsd37nWxqfGJWiErijVvOYxJQ7EYm6SHiVfEv3F5p2A9G9f0/wR1kymoS9kWZ6zZWeySI
bwryo6Uvm6JiIdhFL/KEfXQLtk3oLli4dvN5uVekofkZbtP9k+cTt18VnXpv/Yb9Wm3vh+m04nmZ
n9p1sXIxkuMtsumvzJqqtf0HNvSB2YARkTZZgXYfa2UXt3TjTCkTrFbHa/nM3KrxPPN3owez8U6r
AMrGNun9cXiLwrzS3OLihnZj+bfedg1QipHrXniyonz/muNMsAAbJA3kK0iyIu/wr5NN1h9WoCcP
mSCUR80p+LuCRRip/5jFuGM5WtVxO+3dL5rJnHwS2Mhd30EzO2NblJ3/J+qwFMMz6ELmqt9NUItf
IpOv6T9CnMLWd81Lx4FiR0wjMEBCr9y/jPpsved849OCP8P3V3uTV/C0rCvl9evt1+vWqhe6kwO+
+VS6LEJ7KE3LYbQ2zwSy4jlVISLakGIBoFDHaBJYQRV3VOObWCCfO7Pa4Ee+/1p2yRpeWs2hnXe3
wdeS7iXY5GRlxoPZNfqlkGql/5KFoJTtk8PcILRYvEPA/WoeqDKIE551g4o39KUO/TFEukU3D571
yV1+R/iB7ltOh3GCtn0T3UhZct9S+9JVNB5akS+6lOs08lhelr1PQ3dTm56/Dq854KrRDCRWNIBZ
fAaRiZkjjxMARDLVfApQXmtQCzJrdVNgwPlFEGk11HrL2T+uv34Tf/u2nvEKwOwxMlTmWSz/awwM
6c+MzfaYAwSEwM25qi5UqR2lO8LRUCTP370rfZdu3Fjq/OHzw3ANjOEFIrcbpng9h5Qz2CbIlZ1c
a6zENYSE/diaX9W7jUSyx392q+mrqG7euGBoJzniY0iWnYhxzDnSeaRecNhWGUguRTOn6wEJ+Bnq
NBLjEfZ7DzQg+RviCQw4NKz1O2SXTCe6pAm/72bZYzuGAnqg8TbWvfabWkHN4yq7YQ/BL56Hzmys
VyG5OaeUXsF1JvIEg14/Az8LD1kbwTyJha59mgLLwynK/EdWhcOyiEFOesy/dS8ImMJG7hCU3WhQ
l/7aONpAepNMYtTnB/510W4jvIUMTKsuE6xYUM1qfgCKm2OsCTGlYQMJ4Sc/XJbBkUrbCKHNLOG2
35ilEEkwBME0xeYupNspc9BmmJmaE+VIQUHSF7s/bU6HHW/TPAenI3WxLfxd+yxefmTRtxVob5is
oZTABa7KlVhOFsETF4ktc0uYc6a8EmphmNJ+tEoD0zuywUmv4RcAV4YAm4rPnUU5xTUutkMNku3B
QW4hUSmRreOYltu6vHFYXzhTHvZD0711jSWA+Or07TRuA7EGiKHmsdhFioLQs4RmHCsBSrcgYUWS
thYc1+RmuMNHx2JofFG7m8qGKxLpIrrbzYrBp0K/h/GVavD7DiZWqLmA87VF3e6vfPpOhlqBeHdq
OiXEVVmyPKNY0KpsEcKa95gWZ5XVDY+Ahi1h3vWaWluZFmXJryNIi9fZvUmdslPH+6srPHfB3ttH
7RdRChDk3zfpclLczLnsPnhzQKNJdBgw0CRXYMCnpA8OcvDPtdliLBcCOUNozMs8h1yss2O4vOkN
6fbwYHkfIBUPog7b59hp/HBC1j+9CEGbc6VUrkLKlmAk9AqtiBs1Lpn0wIfLqxbqf5Cqiws2Wtll
pV574gEo6aJbAa70dLKDkj6yk1z2XeFa37QGSK8dQo8vxWVGaFBbL7tHH1uC2td+qgGUfVarXcdm
Ys0O1jDU38Hq7ETd8ikhj9bh97VmOT1dWEGIQt8UejcNT4Egh4Tk8Mfuqx5fLkySQWeE7dNcer3/
zh4DsAYzLiQeN9nBeV4gYRvW+VtOMBpLOJbZB81IWWDC3ZIkSCuBk/abv0XjeD9xUDo2oAQSiDpa
Unah6N58vtB98/7YTTZlWJmk4UdYZxvKu4La3t2S46N/brW4Hc7ic4RjlyuSozI6gZxfW6sDxyTA
/WaDTbKjQOrEvjMGm0JCivn++YrRfu6WIu68JKipD+a9pjfavOUmcELGDAw+F6iV1EjNRzs62T8f
M9RchdYgT+RR+EqvI/87C8kw9vZ1Os8gk+wxyZsZ6wq16g8adbFqNB/X23rP9Yx5djiQm6noT5JP
HJP9kF4JUPGqk+ASCt/s8OTBAJWyOu4EGj713rEiv299COkifzxt+PuJvBaYQNGqZwUZrzeQnqof
aJc0IVam7iIEH7hf9oKMf9zKRzqVh+6pMDngTLGveJaS9Hx1/5HeRPBfSufG1m79m6FxStoaQWLX
JZ633aTgVPCFzEcrmmxHz03wvcIj2F87DTIO45wQ1dip5haRETVMhhMzDeNZALS57wLlkQMhtEgP
eeGiFE4dBzHTGKgNIe71SH+EWDp8i3afcGnt4DyWfyLG9PEQjQabZmphlfqW1Yr0zFnbH35yUcAe
pwO2OY2GDpSO9rKum69W6a4WKrt5A04lCoh42TwIMTNoIra3BYVfCw2elFV/tj7GaGqYLUK0z9cB
s/9Mi4STjz0vOX/5D3qnSbofFXTyHiyUdZAKE72olX9fx1LhN8L8MA9YuMOgtJDWJn4zkeid4I8U
hSW/Zo6fuz04BmWmi5JS2ESJgpvAjQulGPpSz9V/y/xOojfWZwhXdtPMbEgTSa7O6ZihtMfoa1R/
yTrjSRnXzz8Ca1FxolmcVPc0N1wIQXeaqwg/EGkaEvB5U3gmHG73cNJmn77vU6rk2qO1ro8WSt+7
C67CforXh1qFcgg0zK7NzMQzUXhG2XSoFuviopsKcUzA015dvvEGwYFJOZf5R9HGFbvwSQB9HwKt
F23r/XbE3e8ZQeXaMPFUyrXDz+kDR4FAaKjk9jagsM5MtLikAHXNTLZwdPMSui5EYfwvr7Kd7D+e
OBG0yaU1QHrTKV7loq8fBUXj04efilZ3YmM8RU3jxXu3oVKmFUwR4FHyBxChSZVnjwTEw24d7GBe
1OJ8mioD66oBQgHSX2OOWfzhEopBUIAylb0hGpbOlh6tAeXvwTMDPrBgbRnzXLKsVhsPnT4wi96M
92HoaFGh+yvE2TxgPB2PtCpUuQb7UEvkRTRwWl+HhrmszNW0QYXMT+IvgXpidKKgVUQvXsy7P7XN
nhv5IMY3wq/O4BbNpBh+C4fZkY0OggGXaeQlY0Fnh4+NnPOc3yunF8UTaqFbY1NEIGqvoALW+8fr
TAsqWv48ODhMSkdaVLnZx8ajcu4l0XIXRcNZKEzZ81bSSkWj9BNXoFtsqFrqZCxYKS07P76wIvAF
34oDcWKZfe/veaAnl78au+EFBJTdQD8rn3fCFI2UjovUfPrZXSzRzL1B5fEGM+SCq0aPzrq4SmQz
zRCPM0oLDHOEgkzZ5GbBwIi4Xr+8IcrthLpup7Ga/RSjFb+74JZbhmi8sl9Wk4OMGQ92y4h4Keh8
hACKfPRMYZw9GIu9EGw7E/gfnbJEQvXrYnK0T6m/ubk+JFMr9B7eY/fQRnRkenB72x0Po+zUXbh2
BOS30caqr0Ka3OTwq8YR2Nog+rYFd+Tbygm6rVH6k4A+I8UuTsSDlJkE/E3hSO10XFR2O8CU2oeX
7BUGRkCfveKkcUuGp+AB3x4CgCI8gFjcKcB7x0i3VbO8dOppsnyRJJdLgBrPq6mighj8Rzx6x538
y9o2X58TF72BVibmS1KZHHBa5nQUlhfX6o83GIOU6tB7IChHODkw8WvrLfGL2Xeydp0VbjIWUWSj
oAX9QnzxRw/8u4RsZMVhHOAi/veuqR9PkIFiqXDQfJA0g3UL7v+jBuUptmlYCbKgeR2ZSyGuBNTc
2a+bbaeFtocqH+jyzompYY9jbcRTCm+pT/OQvU0h84eBuAJcy2CqfMQ2QFdNQR2BaU60aEHoyJoC
IHLjk2dTwBNOW+LHKoI7VwWfbMcvp3muFGJ6L7j8c7YIG1hCBQy2e8QKkm2+HEw9sN8hKpeOl2mb
t6nxWgE1ch+M/vBUxY0J56/Nu3tHCXCBoAt7a444O7pQ2Z8cXEYt+wNPVXE5OdEqYG50hC8XrUXR
tsIqbHDnIYwn2Fb2uJRD4wrqxceaVqmDqJVFYkOo8vAOmN1r4qf4p4TRohzWLz5OhZo+/DNhKcuw
M/f8raYF9AllzIOab+mBgHW41r2rujILw70gAvmvD+LbWHpQiKhAjjDPlnKPUj3fd2JXgi7N8euv
T3l7Zlh0wmOYjCks96PiM0TnYceiORygGQ0x6JUzBPG4BeHhys/mqeNyOc+QLsW3MwxsHFvXnJxX
vCd4+k5C7LKnWpeVHaLq8U0IbhiJ3tLuWxlTkPZ0AkVysg+a4i6ePB50i3DdiGj5igMwli0fVpi/
8sBzMPgFGiz/Lnk3zwN257pl5CNqcE9qGnd7b3QDM0v3S9Uya+u0FcykfCDqSNtKldSEnY+z8FPq
N7Vx6HNshQU/Cho7v6Qh9jZww+SmVaEP6+4CEypvF1KL4vBNbOeRJMsYSy2nYd+b9Da5hKDwOWOb
zVYzjvx9YZHw6vBhq6Zpnuneg/9KQinowM39Rj2CXMbsysgvPW84sv38L0Wfbj2s7zOzOwlv/SWk
j4klo4IwQrwccrpb2oq/4Tm7Z/t4N4kFSCmrWfA/h2R26+atXA7wvIUr3kaETdIV6wlsCE0Vih7e
8yJzFUjdkClLLPPl7H2dYvfS27XfObIK5F9/dTEhWBea0J1pLpCf0f01KFWx03LPdlLD5tN5sQHA
+wut1fGboLjwBhtlAJ4cpc+gBWw3Yw+9BbZ3GIBK6VnRcD3a3s9h6MD4lZX+udPghwhH6lGgPjfC
itUINCVjck9C7Ad4g0TC9pqaiGaaNYDdCiky2o0J6zCbcFtY2c6bvgWeaC48oGraMpayAOe3Na/d
8P4to7U0THOlMJ+163XSJqri3f+4/Lm72gxDrETAt3/ttGW0xeSLbD3rw13nIcV8l8Z1HLrHFhun
GYv2G5lk/As1lBXsKDemHzVjhPK3jzCJHRK6UtMuYMnfds6ANBldPw4RmRfuDH9kLd0xBOqErvrM
PTxowBgOp4IvrM8cNO31hyixmxTTWZm++DKNQ8TJEB+08EpXVcxN6WBsIZ+MPxmngYf37OfSs4TB
f9CCb78UEoviza8fwBrx65hlsWatv7QBOY5UAesxgHIQdwrxocecnzDt3z0RyxbH82LZAH9SDgxB
O2+wzU0+I8fWC3C5EuZXWCBvpbTq/KzLMa4ZNfVyvs6qtkUbKNnRzyZYHfQurlHfyXNZnAarffqi
P7ajAMFraxR73wi603e1BLWLfCH+NazeAu0dq7Sly6cZ8xOChT7ZPRJ3wp6UpMdW/a9K+Xks3fGm
hhyFwDG9jmWxyDC02j2GeAycCNyZyaIoQBbPkcNDEIsCZGh0ktPTkUBPuqA9skdfKH0k8flaSOE/
LFANrjfrJZEdL8OKc06YWE5qcU9zBsHUQ3lZcm5oDHgPnbcNxo3L3bs5pcb0c3yvYTAp7HhY0WQt
TMMj+TWPO/S9KZ65aDfaDLZx1pMCOnkuZBdP1UQjBsaP9ttr56tSrY7RGAVFaXo/aXsijdMKpKod
9w3PojasUV1/Wjc1o2/S372h9Q5KYpCZEEXmgBqxc0W8HmNAX3LHZlAU/ftUJigasHKtX/stGA+t
SWbu7R/rCnE7/7Bd5mvHt72HjazJXAmGzvedtMMQs23D/Vyo9vELYKiAiDfL0UNxupx+Pn6cvnf+
2W0BtymjFz0p81IBE8aEH6AJF0Sx2F2trZCvds8GI6rSmB/tJxrW7sigxo++upETN9JTlPCtugTt
b/xSEdrRPl6HNC7GMoNdbTrYDQp+xzIfuPxWEH9RIQUoHsa0wAGCkuCN87L9uwqNLEvdw6wuvtt5
v7GeUe8ivOdoCn3ShtYfmkbl+sVrmvCKvnjHnzrSFYP5zpNe4pz6mV0v9f7ClXCAqQHIQqCZRS5Z
XULDgZ7GzSZM90JhuFI0W6RL0iIAI5QHn2sE422VSu1f0OJ5kGaVhk9+6DzY5nCtspC6L8jhbEB5
eg0S7NBoVCjDmgmJsZBzx4G44CRCz5R7VNQzl+M+lXi+vZtrTlI/FQtzy1nlQPiwbcGmiuAAx7eY
2MDegEmGtTjsK7E+RWDhCTFgZTKj6WOk0x2VTwBSkRrtwEVkLxbExFKLLYZ/ky75tmHAZP+LOrNm
tRP0ZF5lcPl0S43oadnnvhYJRj5ft/PqRJwHW9gS3TIbWKDQsM278tjtXHU5Q8DQ0XFXD2ulbR7P
SGuvqdpmLDB6pE7vTAhcZT1s40pqJdqqv0lzQE5iwJg5HT2WhCR6D+DBZDNfqDg+T4BEkPyu/FK+
uS26Xysht6lBYs3mFVpWxY4HqFl+cT/ebCapT7ocOyddbjxYebTGf8Uv1MYVuRuXGx6XqenYCAAS
ashVU0u4ARkksluT9zbcgDsnjOoLpxIJF0Oltb9Rf+ISUw2yQtcBQBNtbQW/+HCGvkrEaJZQoGPz
1OCZizcR8DLlOpUx0JzciSV5VIlEPdwYiFfJNJ4aGZp6ej50czRUmAkOw8wNCLoyujrXwXXHLENZ
iRpBvcKM5H74DQNtXABsI50f4ZbI6pVJt46FjkCAT9MDFexDqcV0NRq4xKgUE/6jOoXqQMHjLQLN
3uFlZFHDwwWF+l2upDwdxfoY/1LxGTpvYEbemL1utbn4ffyDSlWctuIL64H0QUhW3cQeX+akVRW6
u1HACM9+Kq5W+UqJA+zUAyB6DzlvebHpkxYX9hbbYb8DjAOLZgz3ArgdgIRDxkNM4pO+7/4ZvJdN
WUfNG8LjM1SSpctiA/8QxIjgx9oyzTK/AllR35xxcfkt/QrdljTOviga/FFv4s/ROywlvu5W9h/G
fwMwyn8PpMolSlIv245Bd0VyYCld3uS4rW3lSkVu+/k1Jzf10b/FGlZivb/2N8ijf9lf+iws4jw8
HVRyGIs+bT8dhkStE0AdyZZ/6hIi0+7SAR9y6U1WfId68UByw1MOEnuzqME5A0/OC2kiTvgnMj2f
xEMC5NeTqMPHx8CjjU6RaijShjgMddDNWctuVZqgy3du7za2kVDUL631lmdV0uNiLS/yWkkeB750
GW8kZthFPoMIW21VByUHWjozFu4q65JzJn0fySQKeAL0BBhd8HEgD75HzXjc/k2HQCs0R2zTdOXf
b0c6rI1yYdC0yljZ+lS0SSmsB+M/nqYjSwfGaollhzcTUxkys6eaILVr/tr/WWXlpegcxRnK+vgf
pI5JVjhs5MxOJ8ttgmksKNaxjB3TamMdz5a55kJalP1mM3TbuBPm3JWyS6oRLP6ScTMLtJ/vtCyD
SYaGim/TjKOYAcrK7ImtZeEFaE/sApQnoEXI6YJeMv7rTDO9ToBfO/7GAbYPP995Gcb4kjo8O42z
rau50th2N17qAGL2ncmxx9sA7cE123iTsnA+E9uM2K635ezaZeyqD99KxQfn+Qli/l3q8Lmppfyz
jpp60bLIdaQThN+482aMUXhLFGMCA4qHVNTM2u1NDQMSQUxL5vsicCJ9r881kIJU/af3p6/AcUAC
i4j91Syw++zH8jY/zFUdfPAhG0U2jF/BvwmS9vnWT5Laq6+xT3iBTmZlm49zTdXilZmHpPHe1mlx
HJotAYrsfj+X8VTtJ0tSXvFy1fWe2R23uJcRbKBklniCmrXw84VjHxTdSSBFi8ff/Xb1ZapsE9E9
/dpGTgJdNm3dJUJm18Oj4l64wiATyKKQwZ815l3gKKDlM3kI7tPKvTXG+EQQIcVI5ZkiEH5pFfUG
u5jHX86XTY46SMs2hDZ2ae1I6lUfa5J/h65u625y/MaxDcMXm3aeVXYr7HAwHZhFAaPjlIcbYF+n
/dCtIL3A463Ar06cYix31t1zcHHa0izAg7AGY/Z36XBS25eTuXWsgIBv6eiVsIAaFZ4bAL5RRVZs
zJQ47cMQmhABd7f/IgVYebZ5vcsiPu1KvbOE0MxfzJFTJkU69eOx9hB0DUY6VfA1kUGEy08cSZ+L
aBI4G9k14ctdGSCpjBSkWP9S7WBe8H91bg8wXdAn73EvJlNyMR2/4T4jrcPVdvAXmyYTI2v8hWs+
psF4iVZfEmSEXmG0hT8DsFYeF7QnRKHCoQpxViZGRL28Q2JeGkUwX/WSWrY8JV6Ekgu4cG1H4RlJ
BkRQjNW4bLcPT1nsicS3x+i+YjdJZR+mUzfeGri2wAewosWq6N6I2/3/zaY7JR/yLaf9ln3AC21x
90sS/B/C6e9EeV4t+hB/8bwc9fCv2bCJ1U9Bxg+T71KqiYvHo1KUbxXyDsXgw7XV6BhyOCoG8eJz
S7uHIG2EQqv6jn+i8l3vAOqS/y4gacggWHV1agcgit/ur4nTqz51OAr0OecnF7yL8DuZlCjCXYT/
m+DYURgPjaJeZcdnoyCMAy/IsxnJxLSPh78GrYX181opglyJwSlRlPBCP1+RJ+Y/o8svXHeWbefL
O+2+DElQzvXYzwYRY69r2FNPE5j6KpoWqvtzxU09Qyf5bkuJa5PSwFhahAfrhe9cG41AV48hi/0W
KaViGTxG1pbb2fi8G6+3yrsbnvlC6vTkGfpK5pBBBRTF0HWRPogd5fuYFoWRrfAudrAbg3j1K+lq
z1zNtkhGw2WRGbyHse0uxUNvqapvAnWSbx6MORuV1X3Z//HPQkUDapikMVNHBXin6u/A6yAtXSlI
8al9lOwe1Sc7YhQL3NVpq43mM42n+tCSG09lN2Fob5nAKn0TEpdYieidj2JCw9CosrlxnVDG+GCT
yp5mHEMgdMc84ovNQWvKG/QiDLspsYlpZBXNXjgTOSJ2VL+W/ERXujjWtejf6EYWDZhw1MEcDvsg
IJlbeYmjWtlOXR6JZkU0OVukBAKDx0sT8yRGVHqtOrozA2SRr/5wa739ls0fUEOkdoeufNJbNxVD
bl+njupgIajXuGVhpW6QsfyDjT0zT/U6oKTiLxrWp/oeV6BewYhBrryIjvxvrTkC/waSoBXc4vmm
reT6gZuTwQlLQxiLBHSOBJX17VkM4EYU6NGU8UyTdkvcv2fueefxXd5uKZT5G0Ak9VrfTwzG6k7L
kHmFGn4KFjGER0MQVNdfm60sqX40usbQ8touN/GwpKhBQuLtsyIj3sAP+vhUQXwyJ2nMJ3HMIVkZ
oEcz/MtNttPpuyh6Q4Cvav6BCqa0d2zgoUxMxJ3nya+/6x9daTsx3CI2mgVZrFjmNOOBKzdeoJJL
HGoU5Oiyl5wOyZk2JtEnXG0VifbW7N6HVtlEckBUPa5ie6R15Ni2tqcgmlaWbf3aXyl8aJmh4rLG
2Y7rfI4IQwT0tyWduzU98B+2enuV67Cj6Ae1ieBg4YXDv+7ZFNsKePe0Z3Chc+gNgqcZq5PJhiOB
CKqHRkVP+PO6t5Vbi2ZW1GzDyfDn9VpFDA8tza+AOPgKQ1uDMxAvDsXSBVJBF+LHr7sqU6WGDpXp
R+h55R79B0Pza0MWK1BWL5/rjpWeOMkLenUJKlKSVZEZaKNrDOYaRLHtadyJeph3MFcjstgC2prm
pR1CbApRjXp+w9Fx+/jGJhFGlRFhTcltJp899Q0hhxB2t6BczH+HBpS3jgwXckNo1Y6VTQaf5R/+
MOwIsd3CTJsgrszW71lNiuilpl5OORnuL0dnEar0o3+RDd8zAkTwkyqq3RlMIeVuLNUX6mbNKOiP
xNLPlgnNGLhsuKj+nomLkIzZi6nvBvnszuItyF9HXfhGxitmzErfm7Rg5e6dj7lqrkjWgKAiOv43
s5sh+OVQE14D2/txzVmpJSYoNWMn50tX1IF+Ywt5GYSN+VP3kCA+LcqBtBOkd39vgA3VfSVg7cHN
DCse85QSD500YaCJoD9auPsO4uulXi8lmiGuEYGc2dS246YDmeOc/Rwo+2/aEb1m7mN2ZQ6aFlVJ
DcDlbJbUtVcNMWIcd0jiYeM4b0mOPeTR4b+sU2HACnuBItKsMnk4mTq90wdCps9i21J6yilTmt14
jO8NO0q97eVWV30rfXkqAUkeAnckDFCPE92AWAmKahV3OgVFq1MXvaBLbMKMU7h8YjNqsxG0dR4C
ef28uxSY+WOu16DeeKCRaKjPNIWRQ3tWTDEluPuZL3rk2nUL4y4wWJRIm3lC4kRJkdbbZNRk03Xs
k2nmo9sBMT8LAZ3g/d0hDow7uSZdDJXtwcxo5+JMkC0Vkp9GKS86IOYIjS1yva0oE2lG80wAoTw3
QPlH0tO4cS1c/qu5qkoXlrHD9fH7KqTEHcgxgS4kG5s6GOSkUuHJTkkvRBae6p69rO4QjBvcRF6R
tu9N4TdACLPujisVc2Ez4L1oHQVjBv0JOAGpE1PlAr7H6dDwSURJrP8qHv1ym3yWp7mtzbUus57b
AXa4vzq9bHBxjI1WJwfVtGTNfRKy2P/5XWxL14goDAtzXG5EYWKNrdOOLC7U4lx2uAMbdZ/PE00k
jRaj84NNPUuz7OrDxQC6j/78j8XuxQLs9HgcOqb/khn7a7X9XYlxAtpfX2XIdlQt1le6XCw6k9LL
iPe8FkiuI5l04rhbtAYPe34Ddxfvg4pU/wyyxr8Amgvrbtqan4of+klfdczaUVvFozSxHxP8wlb5
mH6D3kYR8nWZYH6H8Luw00vgekYMF5rAh4B9PCreSlVK8kfHI9BZhWV3i+2aMPypppFGahkY79L4
u3zvCz1poG7cNZoq41YMVRCqEAAK7ji+62cChLiNVNIWya3Pq7Pqdgd/a2j44lv8DJ2gblPNT7VU
GcowJl4ivEpcJPhpawyQp59FL/eVIG87+R9wDRA/jNjOrgl0MPoc5YRF3vOobfjgan+evekRUIR6
IVZ8JtUocScNix16d+LhUEfsUl+nZSbIHI4XIMDQ6Pp5pXa5F7UDFYt7Pw1FTzk3LKCaf06pBodZ
N4tCyPlIxi9I9+2KfFOrLIVYEQExuOjjENTggaS9NycARIyrJVmXQ1ZVuuViHm5V2cLwJQ6r4kOh
9727aK3fWShHUc3E7TwY2Hx1UHR5AEZ9OMlzSPgVhvhGoRG9AFXHe55fqvzq/ZvDlH1KITJk7axg
h77NUe+jTYOOk9cKafuZuosVmLAwoOzyt5XT5gyuVwCcRYsrbXOOqzajHGG7Vjcxxs0veI+fqniI
l+/icK+Vax/xmNJX3e4AywGtL5Dh82sXN3Jb6WQnK61WqT3mT+UGin11bTHS2LTd/hWxpRXbQrMi
xCWeBIJPkCSEbQ8RqV74OumDRjAse/lRisyrtc/tM67/xd4AAdMWbp3+XmlXWB83d0ZdV3yPRhhO
Jsu7nEFrtJdoeyqWqvrfjMXkjuKkFkwAr1PyeOBziuz0BZLeaBSCAOD0urdNQ+HL1xmMHYikAj1z
mSjumoJ7BU9EU0E65ADMndjBniZSD8bGUUYRw0aeiHTtAqk2OD8g92NbsoRqIrV1s282kWzJmBPi
v0cvFxyDyYGT7mSg2j0HYdx6cF8RirjLTVxOPSZmlC8dAzX4lkD0EO129p3mR0pT0PmtdvGgiZMP
VElXcGNXPTsjR6OTImVZt4C5MUOHnZV475VtWC5+hGZKWqMu8VBZZvwcxZSJ2eICfkj9/+uOXC45
drdh/4XjkAuIdygYjPwZGsn1v1BnVVyy0JNx7PkA/G1wdnRcrxn/f6k0xbLD90LgIUjK46i1p2xv
T4l50wneLZkt0IE/qZs7GAYX1d0FPhu/xg9mElMwNGIZwzxQVMwFoUQuubAQzC47P66a5Tzkl6iQ
P9F+0LydKwmjG0X9SgDUgl36pcBZtcF5EtqCm4uba1hm6EKJqe/NOJgLgT720RxnrqXWZGFPaGeG
PMPeMDTWaO/eDxVGZ119Ic3B5IP52eghPC5eMAi/ieEjbP6uy4vv3KiTx5u5Sd7c0KZoGm9NJKlh
6kWHmtOvtBuJF3OlqeFEx75SZ2VkBc8FMQlmvQkaKBPJ6IvXWeXV1ZgoIpVcAVeKO+AQbFk7taAI
HZLIzKD1Mqp1ntgUP/lsj6c73pCiGwfIZ6Qua9EXf7G4wNm8YKsQ4M8rGYEyuvxh36fezdA2UCfi
C6WCRITdcnCH5x+dUplEQFdVIUK5El8JgCCcJ8jPydyAjWJ/SmSJaYdpkJeAd9sH6M7qGwA5o3+3
2Rh5twTTS+EhqzL3xpANe33QXFaeboV07LgWo3wHjJ123hBYVDCBoEBIFovftsxQ2Id9k3o/OLDP
LBr399ZnUTCqRyV+rdBowEtc9aEfWEYAgx+KWLSkbpJGa/kpq+fo67N70ICE7R1jxC2rT01o9UiV
q+i9CpjTqPHPwgnI42nPYVG8BiQ0UlEbjJMf+wLDgj6FfFbmFIK/bgfPP1aFrLtbL81HZ6OrlLri
OkVVcpaZmF7q3c3Q4zfkBVZpmucC+TR1R0+Lgx7HqhWPqmqKfHGDvN6IXvn5ZnSIdDbU0v3uqVQR
NWL2qxCvbgdKvfvFc2Ol5oDhmnoGkq22shiyJsRZZIpMxtBg/y6OQQF+pptzohn+40mES7uiqb2l
oQeMB7s0+quT6xmL64OVxpzfs2UcYLBR/YEj2Tbe82rel9B6zc0ABZB31efLOZ3CIudlrfJ1iDj0
+8Ra43wzlDByhRyl8lCzo4FdjWYQBfo9hljtLcCVnCaOtnVRwLNjvQ5Uw2RDYWdHxdnowxb4+sPa
pW6N85cR8jN4wLIlSkM4nkgxnNzdYUYl/mvLoTWzwpCUfyE9Koc8x4puaq+WS/lyPUnf0NeIlPBg
PBHYosbakS7+SBSkz0fJUnmhDnihfgLSQbC6fpj8FYmvUqRai9hRFXSfN72WkccMiHsIxWgloclO
cIQZRbskP+Lqi6HRezWau8ZapzUJNpxD3H7ASBBx6kG3byf7BoQWKWQJ4rgnJ6CqB3bU5GAFRHsc
EKupzaLxN8Mq8hciIcnDp/u09bBeSlHNRyzjf18HGsTrGKDeaexWyyxWoSq65A3wm7l/kkIj1nfF
ZBOOKTMpgR2BeLKXMA+OfZYkZijBTJXkHnPjMpMCZskF9zJ82V6WyST8+6GwHSii1EicnXEaR9Bq
3OpFHxY4kqLN+RNchg3TaEwSu/6aMHfHLPvY1zQdEhVsC2xtx1pDERSLKLgtCfc+jvFNNwjt0fkB
k5v83xM8l2UqTjD5ikTyz+iD9yRAVuaM7o2l9AhNdLA/c02DEE7JixqawHsO2+ifEnJx2/4+P07C
krH5DUz8515BwAxZJfKMbHUXlcgwHr6QdFM3IfzXy83c/F3Uw3tadJ2Xf6VP2n7/ee8Mzd3yqL5G
4SQXVIRAFyfzadeAy3l74t/tSFlYgNY2gemBgld9SIlEG9vREH0E8BoVT51mfpgNN2vlVHICK9af
iK2hbFnOfDTF/xzAS/GPmj41aA6bfdWOeFRDjrr/GuReBpkSlZW9GSzIAu4nf4TNCu45nzT1RAng
S+fwDv5QHu8N7P5JEcKQNZzKgKxYi68wiENtP+pO25EJ1PgBg2Qga6PGXV6upRUKW15gbDOjAw2i
cYMu+Snqa0zhS0ZaCkcoXKjQg/tUOPlWmtIOBsitIzqlf75VByia5ls6DC/nUeCdtBymuGSN0SIh
6yXbk+uw0plLCfmlp6oyZyB1iWBrmogq/D8cloIIFj3Ftpq0AY3c/rqdQqhY2PB/zCQGAFludOPR
x5BHSq1uHWWfhvjHDCwEh40Z5yKXnWG582VoSjYUPAd15oQP0xRl73JXG6JZfSnneBwt51ilqQc6
cetZpczxuj0oBjlRVX+h6vg/T0Tg/W1OWH2u4nB3IlvJgS2/bb+I4Ub6TA8oZQQfXeKKf/l83SBj
ppOgLpKkU+3J4OjAsh7GtXzwQa6G4Lv1Q+CKcIomb2EiTVjYVdZ/PNNEI/IxSqWqW/ajC7dNEEi9
z7pXhZAABCqZBi3UQdrd4wL0hIfD9fDoHt9go6mVVgiT9+0dJV2o2HAdG/HRJ4alp6VrKpxNKb8N
yamlS1XsoGBobBlzDSU3bTOmCliC1dSzJwOQuFJ2lP5nsdgpPlQrvVGjzOLyI6ToQ5OHKp7d6GuU
kFEPsJXYYHkt+fUvPNc1BDWupERQW9UqIuwmXCxlgb6p5Rn3VfqVs2XvRNoCwiVKKCDekfgwRd5I
+XCAUWPoCfxC5EHZ56DcyZEJvFAllFa4rmTRwq3SgS9vz+K1AS4RE4RoAF7J5bNgy50LnbaV8VaE
6IhTieth4FmfXEeJ8nhdg+xU6DIHYcfNUGmy3dihYbS49HNOE9i4qurdScysLWzwudWtxHtars8W
UCuf3TqHs93XHurz9Sl2K4xsRuSzZOcCZm0g0kLdcXncdzmB5Cb3TYr3AkhAG0mhPaeCZfO2PFwl
uALyz7iY018htMF8zWiz6NewGd24jknAWFvOnQUBN6X3GXSpsb5sLRS5gMa2rhSquXev4G9n0HG5
7f3vT3qBw/A+1XvH45Fz8bCiyC19XkY/08NM7u8g2iOzrWBVyFmc5b90bGYg9KexbSMhDzW+GWov
3XlQS+nr1N1skTMbdYriaVC3z7+LNdj3DcDRh3nlPzzj4xR1NiwRt5qc65RjRbRHREuIWXUgJ05C
/no3BKNcL0P8fqdz9G7famq5fgfkqMj8Ae93wmTdiL8BbRbPjyPRJjwIcY3qDm3XaAApvKdDc94U
zdjp9w1ivwajCaQ4NaUxYMjANw0pGQERiIIQqbmAkNuA5qoDV4/QBanjZv4OaL9siPgh43v5omGc
zGEmAYbyq7ZspDsEoKCVrZTV3ji0EXQptFzj7hXLVXljXehWx46E2DxbLHV79T+9uew2LF08lBXM
HhKP8OxJsm1eSlJPVGCpdJqop0vaxyUUprKmqe6XtSCf3c8pz2CALbLAqsHtd0uDpEhzWpnm014C
uvW+yHxlnUgkbLr3TOeI56QDgHWCdU/w/pAjgVFpdElajfJ26LvH97khStIDR3yQgrohA3FU2Owh
+/E7RFpMvOx9I94TYhZZTL7DOrFq3dV69iLjw2xSuLZ0Mps3hzgyvzgaRRes4Q5jD6fLEt1BBTLP
CR7CFFF0EGq8LrQkpmzdZUcRvUpq28IK+RXmhs4fFGhhdhoQ9QQswre/wn6Wle3fhAuKR+RgC5cw
ZdeIy1itSzYYl/5bc4X2s6fcZ4AeJhCLKRB8aOZpXJN8eKECQ+cXpsXQ3fRt3XdaHbHXogkvjlZn
AGBxVRH0uFMk3WK7pSkg8gr3IiPCSEuwJ8ulUVs8v04T4Nxa2G9fULP0JwW0L1AQcQ+uPCPsptL7
cqujBK2MCbOyFI+OwBw97neeCj+J518tmhWgea6WhF1lBGFPHmIqZ6tL4XYQSwqYg0AcX7/rKhWy
e8Jz2PKSuqAAFl+vatx/OR8NH4FEAKbWsFMll+KNW1uEyl/sAMsxWOWTLKBs2Ap/4ibhQ5ml+i8V
xVmPMaO/yAvm7CVf+HmAqx3Uc/FoGvY+Ih2YVgCcCMGhFo0BN1o3Ss6mxy/7ZLYsnkaQgZkPKOqM
ypOAbuW7cuzDkfOCHo0lQv/Z67VtYT+KDX9b0aL4BM158z9kArlBZr/iKn3gi9aK8qqIqRoXlI50
9E6Sg+lkOXC8x2GN3hhlxf+jxjUHto1TObBG/kA9mDPfnyBkUrgyKUrnnYsYDgRFLwjo6w3Wcvb5
y7QGszuEdXktSqBqLmgYY/H20OvYC885MWDvnFokXYc7FKlmdXAWh8J5rCAGGBe6mDqrZaTZThdC
R2LBAJzquMG5D3eXhMPjXC0ICAPbEAPkxhFcgwB+epG97SVXs1WnnSjLz8eDRUuFuyfjufN7do2p
gDm0F2qY60YS+J1V8QnYmr9SOPIkvwJ2++GtLdaQwLGUmCcOO/0g1CX20+Eujt+kV/suzW4ck7bo
OqnTHTd3AZg2kjhFfEF5ZKE87KDj+QKSiMzgwOBvcqacDpEzS3bzxGoRoVYlvq0m0iHGB/PWAYD8
xlWeVHY3rQ8XAkwDO+OGdmsofsXS/2QVIQDHIorI6GkuuJ8uEDr4nQrAr6+GFI5KL8IONO0XRyur
j7AYIbelERbdNMoWPsLh9fdiyEUR3lmG8zcl9xa/8C32zCV+rlyrAHNTXAHtSZ+fU+n2DM++xrYZ
X4je9XY9rqb1/W7ZBtCTsO78L6TPElTEs6Y9IFb+Z6AzPuquXlqWxMLvKrsb7NG8zjLZdr+9Ypd1
VZdrl1ww51ZVb2ik4wpZGFWssPHImFrA2TbkUR5k5UrfefyzeB/n24ILgzT9IrjnEZryMrRYMEM2
8tGG0YByBTgfFW1tNi6hKbXGrIe5GcHQFRhmN4gfYZiouUV7MeV7KSRXZliGkxqt7ggf0tYW493C
qgvGwZDNDNFVbXUuMaAduINltrzZ1XFEzdGxExvJ3m5afs+nXXxqMurYcs0HiNDPTkHBFWllsdrP
d9PsFQ5LtMTxVoc/Elc/TrOUcf0wHJ03U4qrH1m63QmIMX/CLBm6myIayJDY1OHFjMkw09DLArT2
00CToi87aGRVr7qpu3UHnr/5VKHMKDD1lQLwU3fsLyeIR5MlZC+KRMGWIFYcavko4U5YdgW+qWuV
dm6+tO9vnH9qyWrnHSM+mu6G0yohuyo6Xwn+1+/FDtmC/prqe8ManYbQ+qnwLFXp996/EAEk46Od
DNW4jIDkv8Jhmpmzsy5hlBi15ly+Yn25uRu7stKi/aO9MF9bFJBeAjQBiiWDUq4pYnbPzqky3SuO
cKmv1xwXJSFRaEh2fIKhtn0piDgq/SHUrwOTrNrM3LHTUnj/9bx3lu681PjoiFHTZ32tJBJNCYz2
qfD6Ila4V++th2SBZj1LN3E62F/enabsQsep+s2kTk/0yDznG7VQIrA8m5d2IK7vIk+/ldyj2IXR
8dgQKXMMrI7R162RFe4K7Sue9Bb1tn4CGeEHV50nEST0rYllT07zHY5truRtWrL7zAQchgHklIab
p8EKbA9ls+4zMD5086MvrU3pM/mtcLAUgYo2zrhzY4RHvHLPPsb6l+bvcZhz1fOcoad/Nr4jIt9E
WEnqjr0ujY+qKi6cGKIOz1I2l7Rx/RrKIvJ0YbCR8gWSxa6GVaGs39ctleUh5f1ZEMlC/hWl7yfi
il1RAwCulgcOokyTOA2GQL0nKwvkByLrnzICkzkhPeIqWpddyFyvV7ETJT2B54TZuFLIz/5713cH
rypY68qvbsq80iYLy4iz+SMfa1D1qyEo+ODpz8EyeAAHVHhBElH9J4NE+j74mBHX0IpE92f6V/BQ
gqWb/pA0V5tzVwF2bMPONgqMl5oi2bVXPvYn9guxgxcm8FiX2J73SXR3PJ24JNkozvXrL8RpUD/p
vf/mD8Uu6mBgZ8sH8yaOLTqRZlYIC/FeDUMO3Kf3WJa2xalQdQKenVquW3wVyWFxk6qDAMt+mRLu
x3HtEjy3jusc4bBxrVgRdT3NIw3HYDOuTNwi0IWxpSSkNdSMr3cmdt+D06lb986xriTQvGATXVwV
e+VwfCSTW+MUN135uj9F78vR/rPo1siBXHAn5LMeCZT28Wg8S1Tzf6sVgThQ6tbFrsCsFynaggy0
ePMG4ipZ9R4POuBBW1eOdOcO/wuwKPkouVh5JNcNPoIK0ZgvGtClC1NvJncdG9PC8CYaw4rGeeWi
MLfNnCacH7D8iOqbFbyB8ZTlP6N/0A43lDTGE+OUL1vPIngDmVFDWLe414fg6u57OElF2+0s42Vk
tTAbm27PMLap/cB8pIh35sqUySGy66mM7QCz+qVauItO43H6sGijHV068ZgqOwwqEreQUEtWPjBQ
qfQj+8Ldw0nemd5U4UXiK/H7THI/VVdGXVnO6PGDqtJsUOfGWvRv+Ni+nWpzK/zcP0FEhDnWJrMC
LqnzlILE95hK27+Hh+UGe0RhBM8ce0BjZkYRSxMQgN4F0xj7aMLjB/27KTLUcdJZslF2JUFUgwMU
sKpY2V4x6KsBVU4eSrzDteefChR32s1bb1Ggi0IWA78orgXk4wNhq7MOzYOzYv+V8BL1/EZ4c6zM
FFImrf7Fvgq2SIZo76kUPQjaOqWqydkAGuZ0ec/Rsdukpwd7vvs5fmvz9KncyHWcRhR52vvlPekq
ytjK0JP8d2VjojOVtHLr1/sHaou8lPUiyZdf4N31+To1QlbbF2OXAgGd0l6UCFgbaCJaW+6FqZmO
H/8QW5yEKL1oXSksnQQm27wztdL7vw1apOPBh//x98RsbhGp4rzdWn068hsyxoezppDyHgHq0lHL
tYUeh3b05avN3wnO3OW5XDTgR9D4Ob25D1+QTiIO+UZYE54SCeOEVwPFooR/258eqMcDHUE03N2B
sshpL6jEN+jpclnpAwEUa9jGoaYR2zBa5TWr4kpuxGq87wLCqEHIs4nhtatjRzWBhjDUCUcelSC/
nHuYCZgivkNUbqxQzuu5MeKhkr7zaYu1Ri2+O9PWsAC8ZWMT3H1J64j9r+PLQ0jZLS/v6j4mkRip
LDdSEUxOrHVG8kkCik2Np4fZKMebtvWkUlRIpHDm6gb/LH2PIcu1x3nB3RVKk8EZAth7Br53c/JS
BLeTtHtqvk5ilUJRT4e6J+LJPPUIhBwYFGBf9nfhtXWSD1942RIKIuNxE0SbdLQBPdkuz6ClPPi8
uzovc88KHMgHxZrVSv2BKzzxPNwKQA3tJVBGVFHr4LPYIBL//YmZ7h4F2vrU/t83BHDRDkmDjb8P
LCkd5VLC/uTKVuXlgbCMM4jChtjarnOC2tgOGVKl70H+q+sjBO8kcheICwFr3MwyEUeHSVmAyag4
4jaOOTSsoglIZGvEgMy9jJYSkzg916w0tsg6MRXILFhJbQpRfh0ROlXol4AGl6oLNPyce6ZNJuLh
g4bs5LhLt16w3JVCCA5b0cL4UZIYtxJWb6PyuYi/21bTBSKtOPFKq1I/vClXQy98Y039NZms/w/x
IueeJ+ZvbzQubILcEcADx4M04bwtOS+LDEyWslhxEdYnx1J2KkZYvDzMn2YucMQcSlafyYzdrQkN
P4kMZrlUiW87TzCK9or55N8Yd+BHmKxnOxVHrtf0FM6B4LrlkL0uF+trdW+6+LXWbJrLXJc4wAXg
TJ04WUb1EP0ImmbTmdW75H0JyW9FqkKDzedqZVZVngHjt5alCNpeqJXXPxA81ihHr743sEtjedj9
Vie8nRkzXXlyBCekhKMi+urk9VHv7QlbW5Ib1UIgFlT8Jb7hCpzFVe3FrPBaJZL02x1SbGknUmSA
Z/EK63ah2r4RmjPCQeNRoosIgRs/Pq8+iP8STYIfCDAz89CB4cX4UpQGwAGs22J2ATip+m5IZO3G
EtaQfexlk9g+7FuiCq/mZVjUhyis0clCfb8xEUJJp1Q9n3p+JpXdYvh3QO+lVZ/ruERKbBrH6Rbg
OixwmOExQy/LeOFSF5Bc5TSyZbN6GZ/GJ/bGSUjg0+ufCjP74GPrZsaR8TuyHlwh0/akroTaky+w
Z55nH+w8ogOvC8/XA6+9seQMtdfqHsNnDwYYikDSSegxcNNzX4yR0M3dKz7mYSU6nY0cL6rnJuTf
7rK2nnV/hxQnMLZJh0ljw0QjyI/wJhcPYoc/BCPpSTKo4jdTbpD5v7CYFNUvCcSwLqMAttRPz+1Q
5FDCtmSxg5g5BfOHu/W44YEXsaF7vVMhdCTrZWxydLdazHVHNIDr+SZ9SJBKhaMLt5ZlqaYXwwGJ
TVN9B+XA2h4SRjDXizyxLM5Uqkl/63bIULumLLpci4d/4PMhtJUlXWudSGE0EgTJrDrIeTbPrmOt
wAiHxrlMU/ZKY3zhLenQ/GkJElMVFzUE4IZ3Qh7uLii4dmssfeu1vLrx42fV+rzcdNDRmWxiiY8V
kAmBB/Md2ie1ptNJttmUWPTJHwZaBcFWxz3675+d6KtSaxDSlFl8E5f2qQ0006+0TYB9apFeXgZI
CFDpC8Ml13dyiSBFPkFbNDCDRQ4zlF//MIYsAEeW67KRXqlIPL7+3JdhkPGIss0wG/M5Hf6xs7Xg
tWEod/fkjAb+ZohYvB4eeJMOZFodAz9dORk8QM6qFOHQNl6lAibR4dE6pFyAcbadas7awa7SQYEj
HYKs5eyEpT2mn6r+ORt3wRrErZY2kwSnHnl2AK0K6Le3H122HyFqhHOJGdlq0Mf5crPLSF0CBahT
zeIIV4c0R+KVz52bb/EZMPbcPqUBKyg/mK4gKBsZFbCPnfpX7pphtCAeL9tTHljNPxJwf0fmXj0E
jX/VIvP1ZYpbzi3v0+aRTNm/2aohpcYATIAWbtyqK6aBJCX7jwzBrCuoenBz0eVJdzDPfdx3HvkN
T7d8LmVduC+3pY/tiFWJ+4PAc3nCmWTrmNCFDR62T4xzKHsvEQpsCmgAN1n6aFfamvU7H2k4GJ6o
LyeW7HFy5w084Q/oFtEzK7UVe+FRp2lzP60awTpT9hlOd6j11zwN7eH+yXt8rUGYTfDSZODSOA1D
LIy4+0wxee3arob/chGzR4e+zPJ8Hh1tfai78c7rb8TfysMtzJgnM80uSWwcBANy7ADYWKEcH/va
lkItmyBbiMaHYFQ0/9CWgKAtsAxp9QP+qWAoYTOQ3EASVCRCo2HDPRRPztjtdfGPH20uPRD+QVLC
lHoI4IP1fNY3DPeI4Gdfi3wBXDfPGDoO34zHVK1XVpj35yI0gAhXx++zK0TGdxn77CyhntlWdXB7
IP3e10VGBjd3sYg3aohI41+aWfD1/4Ue2DauQS09gcI+VSFJIPxR5Ch1IDpYYkOAolm41tZP2Mh7
V5GhS9PVDG0I/SEZjWSHt/6Fr3Og+ne70HVxcNWBSLrQiwx30Db/o6xEEYIhYA0DFcCX9CJ7m4mV
IjeSEZFKWjPPPcH44oohCuMKhToOlwbl5RcjLHHTNWlf5SJRrizx/qAP+MijF+CYV4+/Pb323PE9
XC9XXJJVguEXmsDulT3Cl9HJOPBrO9a3gJcyEn0mEeQof+oa+MkJxu7DPzgGbz1gNDFWPEe48avI
kUQO2Yqe9F/G1PVQBdoINr5U2rn5Mz6kcRsYa9oXRCB6o/iGkJ4tGB/2kED4la0HB1YCOT9ROe39
c9joWp9UCMWh3bpoBOdbi8c//SI0kEmYnpWR5jWTW2+HS8EAbHnnv+SMh642Av/lt/gTatKblYhz
O1en+iMCUNIfKQwxi/xYR3O62523dLhR3l1WyD0YtOlgxZo4vHxWZmST0jeIHzljObOPjyQMmX9b
liPVGHvGuIA4oo3X/mVqna9x8z1GAi6/kIG+DgBegMWzozqVsTcNuxJb0As07ek18oTlrgq1OmDu
j5w0FKVIcyzuNfpc0e89Z/TNqWdBw/uHfl2RqKqnPNOCHPAdMK/6yfPdKbwTRKxocMTohZCP9vqb
/f0wWkeEMUrtKoIB4R9hr8lqriLVV7C7XqEBamzeDhVAjKXqonwvBKZW8AaEu25Rj94vB00q3Gw1
VQOcCXNLtKAPo72EsQFkjJJJVcBuS9+2Opq8iVPRMnFe/YY725wsn6VD+qgPFyO281G7Sly6kKbs
vKU75+nd6fitHX9eSv+u/HiOSv8qz2odgYiagYfQwCYUpkWutGwDEoz/+VFn8DOScxF7vwyR0nqP
xzv+pK5L6UQSCfycpEpUAcLRJjc9Lv/jRNUqJhi+RZ3MyXjBvM9GRvA0Qxqwy9jXFOAaslniEkmO
7nETe72+Tct93L0ZNdncq7trqZCmwZWbPLwg7KU81WutzhyS+bZ5DA4IF4HshbH5+JJydtWvqWGj
9qF+b/bWohv6FTgW2JpQYPl/S1FlCPiNCczrbeUDuocCnzX1slLtXYITnMXvVY6zp33pphDMCuTj
4eyKC51v2INof1WYIH9eBuMFfd1QKwMmrImc3ykVxhLVbrG9j8EbUOtUO5SLzh3jq7hmm0oEtnIL
H1saY6UGDaeMYP70mroUbxNNje74sHiqmTqfYoCZhExmu14XULZrqijhve2t7rqCefKXIByazjfZ
uzfuBNEZ3IzanS9+m2MCHy8jZNUlsDru/KLNz/243T8rdSEz+mkQidv4zGTSKN9DySwLHAncfWsd
xZpTo4wop+VVNq8PzUrrvTGOQ+pYpojLTQV1zuvh1J1p8l2BC0HfdvNnCDpfB69K6Dl/K26xrFQE
JQO+IKBD0J68hTJdYBS9tPIOgc7bKrRI4KZdMVAfkNG3zlCmASBTAxqrYG3miKlSD70CV+nXbwLc
V6DjuttnVEgYmCTwcQH5fj/O14rfqinYZntahM2merbaadaUfuSvZcm8pnn7nVuTQskv/Ao9YCTs
n0NnvSXEYXrMS+4tl6KTaLi69sk2vhCfSm13CGcboTZZWoWRXQItA04+mcag9bp5ATJdKo2bRF4Q
Ly097bDjZGZ6OhqTB7sjOLaeeoB+c6rajAYYw47RSjEZDzehNiqs3zrDqM9gepK8diwzHYUNw4Uz
TNWfATCATXxJkwwcTWsBJPGz3LvJ0Pfe/sjJ31lZI6aBR9eEK8++gmGqkW2jwujLRctJhLOt4pjZ
pQNcFBJSHaBFtWioO1HvHEy4ck5ZPBOyphadnfcTHHYdYqhg1Wb+yEOu0QLoxzLsH3tJj3YnI1eK
D9I/TXZWq8RFeBH7Wc8MYoj27PtZiEzcuGm63bzQ2JlUrFyfcz1sk/5aNShIHeGVit1SM7WXgpf+
0U4oZxwtvZ4XioZ5CI3JC6fp82bvslTMOS8uIANAwHNsHqahRwdPUfy0q5cn0QHSRzsJ4hZadf9m
XM1EAxFN6PGflg8d6Vew1y9pmcaQ3qAFs2J4T9g4cbBfdUeDIjcEwNH5MvyFcNYGACNvktixmybq
oZUYauu2uiu4DZ9Btp0bXWTUnb1twIBa7cqdZS47UV+u9KH1ODSR4wUnCW8us6YYpj/KsVTMCw83
o3PvLv5Lws76z2FOH9SAjsFzJn97/I+3kPUrXKkRtUI0d9CfnQ6MnFLZFqtWeKZ0Gab2ezwXhOM/
Qhj7OFz6ulHOp333NKve189KSCGR9i5bIlVYgswmcalOD1BtvCkg7BOra53DC0h8f3oT09yWv5R4
56UPwqG+UquND9swpUIkpj7voSkGMyz5R8nAjGQ5vYAYoNithYe5LxNXpmXddMuMPEFUCoeaQz3N
1oZTSGrWtydVG0IvlHWPUTlS9w3jwwmwNjqfumzdUObukvFCkGZ/qXXL/Gp/dIfHNaWtoWTqNW1v
nyCVpSsCC3BxlrQFwMG0KWoPLcNdec2GJnib9i79wM+d2iaAKvMZ5JHltf8qUJFuaMa4WDF1AbaG
0YkG7To96GnjdO+E/pWwRwlEXQ9e1oinFt1zKLJh3C78CMwlF6utS5dzWDGpJqGP1cfGNno/+yPq
nuMNdno6I+nrR7nCWcBxHa+mZ9kahqueXIhLdtsp1WPuwQq8e7j+7NLjfYkVOrGxgKzTHuNxtBRq
EkJMfO3IPuNZ4KCTTDyfqZMHrphjNW7aVE6mEUbb31hL+S9y0bMtaq/W3QfqSiBfU5nrtWrMAvkL
NA5sQA6jt7jw5rHkmJ8wTPEDaVfukpSUHjHwhd1X43Wtm7WnaSCrlEFuKgZFxlydjKnVsKqR2WOK
tUpaqPYprTVwiUnNhdKuU503tD2+VvlspSpCFO9U8ROQyHROxMyp0HLt2IHpNcRwx0oTMR8aySbm
/xhb2V91GZaxG5cwh2MAOmFnWLztnUrOQMo0mwypz0Vg4b/D2Ar/A6ZV2Te1xrYd8/YDG8Tsg2d9
HSywRE6M32gQDiRcHem0Rsvoa2PO7Ed1fLa0MuwL3Je1LckqkEQdWsC7nTQWkx7uBdfdWL8MFH8p
1zXh2qzidSTQY8ytJSUPg9POH0KeJZqDwJKGfQqFocTj9GgPwXERWIuv9Pnznh6fhyid1MmFw+Pp
EniseS8fs+ugO4T46UvevKI/nPcEU/3+vBVPGXWqbA60YNCVFDXqx48CBpOUFC7veAj0v0tBvror
nxGrgVSImxW9XHFJlKfxD/vmqWEANSF11+mJVQI4IhY0SgpzQZrrmIjU3qUE8bnCVLI5LnS8QzHG
9ciNmZ95y+3aCICE+FDY6V954LoCXUXq0jeZr9nvMpVl7Rmwh4kbjU7BAM1WvjS34gWlIiTyjyCz
V1L3pjq6h9N//1wve29XCl/SO9OmNqEcBE3fGgYutU9EsZWjnyvmkwtQHHFGs8FsgkH6cLMm15rY
3K18sxabBWPoGB9VPN6SDJqzBkGQ9UUwcDmSKoD6biSI3wetZ+bsbywH/Ke6lw49QO0ZI1muH6yd
xCb/MKJPvN64XB3Q7oeKzaWUX3Gte7HIOFjfT3mfWB08ectiGIbmZPArPAmQ4YsQPqM4NXOHQA9T
O4+H4lPgkfGaIg9C51mhu/CH27Wiidh+4iWbL/pAM15+EZRgKFH4Yc17PLp/tnBLU0yL+03Obl21
chJidKwFY1tdqZT/t97bs8hbcDtIOtO1XnyIvXa9ph8RaaLjU7T3//xh5nR2irfjsrrrF6Imy6OU
hju6I2mkdt5vySPV2GO2t1UCGA83Fu6ilZkUz/nY0jtqP05cptanzqXE/LxzU2m5xr0Ck5agiDEI
RsqmMeIayH+DikrYvHc7yCTaL3FuK1Vbb8nGF9Y2FOFbSOkFcAnQDoGJ1k/FdooWgc4eeEuh/Yj9
TKZ5wgAbrzFIQsCOOuutJKoxUE0OxaV5WXNFEgH/oiDN+xwUCQnsQoltzfczf78Hzd7MV97TDr05
zuvxlgxX6J8XIq7OjaSnbnnr8rXEQrGP9iA7W/C6R9J9L6B604HHG3mvCddOfnCGJbrVjq2BmGf5
4kpSAO6+ONF++RQf07GBD/Sf6Xu+2XGinzXwmTRUFh5zBfDDAxaPbHm0eI0hjrouGpQtuJlFqygX
1GzEm3HXrhnG7CDkBbsGAQNLnMEEfL1fiuc20pnCsxg7WKRVygsmk/ni96hatlN829AxrhYvcZCq
1M3rKBejlvKwdqrhDVWMok1GP1G0ou+0tKoABnLJAtwfbIaQW3k8itKTUsHoP+FKazGeFqZRybUB
yqRIJBBrS6DqThSfPkZEV62RWkTO50J5MXjOkalt4u16Hg0+Hm2UcBRMXV9f2Zq/MKx95XdDFvFw
070lz2vzWpBUh3rbXrmafafA3TppK0Vz8QCt5XDjrFHfIs6or9YzZqKyZ++9MB80xmK6WR/l51Z7
/8AZ4sbhv1qE8bXNheZA4TYQwyI4WrAAkGlFgPNRiVOy9NDOuUpoKggpEt2/SxDw3cyo3spObYU8
ERcuSoGAZsB7ghiL0LPI2vJygCnas+BGZNkr0mWlfUKcUjGWHROVt4fwsRKduhMmyLHYMmerjMEu
n7o6XSk0K4yYosqOwfHcrS0+gmyzZ03Vo/UWuV18QCXHbQpFqMS521yNx3RDRD00W/GjD+77khjb
pCU1d8ghcFy813v5QRS0Rbg5W657lRyWvrxyjQetYBsEyaHUbtC0mQS+wNPKg8weTueZOUgfsebF
Zp3vlt/2SrxObLFPVjZk1w+AyLVXdHrBm3DZ3DNhnIULpCnl5/PXDYsT3bUl36xIxyCFPLQnrzD1
bBN8Xl3XkdHtDAEI3Vwp2u8TTTIhBvc5YqFSsSRsuLj00+FA6juxC0mlBQEOIeF5SuB8e1vVfDim
m9Vl9mManZAR6THeFpa1wy8VxHRqTpUsNj4NwpQAgrG3yrwfX7fxFhrrE17LCcn8iSaRFi+PkkoK
EkbdRfmDvuv7FTw1bbAr1cEXRpDkkakSgHuTFklt5cIbjqa4Snf6tGvDEH2stmDb2PLuJfEz1xaE
+EMINAQAKxT38js78alzxTSK66yWspt92U74HqOISElVSsXtOcmHRK2ZMoUIsk+8fVS/Csd4rQck
JNyG9C++/NeomPhcIasYdfi2UkYLewVYinq7BEIBHVBMwS6jj/al8HxnKy9ss0jaWb39xVC9mjil
PFrwIAo1Sw0VZum+jcufR23MPqkHg5SZkNY5obrJYVim/LN2lS6JcuEEYyjdjAuoacp9kqg+5TW+
+pdAs/QnJrnxRiazs6Az4Ke7hDr/tPKFKo9UTmUiPpo23CiKGB47UDmCKs1/Tjc3DItVhg7RdLCb
mk0geJj1WwDjM7WXMYOk0W+buqm50agYW3A8+jVjAAvc30iesno4ibU31wnkpye2mMxD66w6x9MP
+ZPwXE57EcPENc3LINFiv/cuMVd2fW6y+9KlNbcDzgAkBSAMsGJUHFR/QvYx5Y/askpEJcmuJb29
TrJNf6JHUlkcQGTX60sCLnb67jUIfWO/ii/duNvxS9GWpOqWBZZmiDIaxy3jybRMuVq14g/yhqlR
sjCj4fkkkCHJC4XkDZ9CowInB7rH2elq3nvFDz9cTcq2TqpEve8OMKhaWL8y2JHTgNhmmL2m9y37
peiVrNk2qZwxpwPLaC2bB97mbZ1O3sspGDFJZDj9ALJb8EdsSVdATmuZjDMCd2b53RQheHKAr4AD
0c/A8Vh4fZqCZB/5RxuByKDlLANut8XzZchyTYlEhWHZla3kf9lExDo8OnEytYOZZSvaQpZPKY3C
l5EnJnhps+nbJ0WbO1nXaCQmIL9v/teGEvJp+Metxv6Q+SD5ogp0HSGnJ8pmY8vEC4P0UQMOYeQr
ty6zUZsMKf+WB+0yehv6S1ayxOMc8ErTHh0ae7M5b0j6Eq7sNl26ptKCZ2ZDPIStFerq/Ff6i1s6
IMNVZx/SU3XoJTC41pqwn76X7Xzn8JO/CckftX/glzYcNquAKHUif8gKRGedQVlZMERnXTyN3Mt9
epoy2Au1yk6z64B3/8RV+DluNE0gZjnssiqp60rnevp9b98U/heSJWcupWOCez69daDSM2m5tnCr
8pSBRJXiiWn/mKAIJy669scnABiL3mDIPgcsiSKXMKRTlUn3st+iQnWhYAKeQ5khFLVVpALom2gh
aWLsosCgI02AaQrYR3smHpZ9tG2mikORuznoYU12feSx5Eajiih8hwBgMMuZgSfNYUPRCP+ALm9W
bIkreZaTaLYoOMKYQARM+yZgJFjIpRSBTig+2VFqYaPNcy7jbypvig2wC2E8mGxVPV6Xk+Gi5Ku1
q/1vEuYbg9XZzZKeDc9PGcasHGBtrAw2M4uG6PnKfQA13+ItU5bSR4o0UIfsyMGXcT+C/wKCTkSg
HpWtzZk7grLcpV+GHJAVaDmUTi0AFGzMufiSFjVaQBkMYXIfaD53DZKAIZBWVi7ciU0T0PouyuWF
EVu9+VnB8YyO1zhtXvWemxGPBhq0pDnarAmPXKCbRZ5gttwifbMfFuJKbaR8sf4TXPpE/g/F+DaO
0FeQuH/jIJECGzlsq9WOmVPglaTJmvlaNfdfUJCgFHsRKVo2cVGcFpvSKnNC6PrDYXgUTIS/xXQ2
90uLD5wAV2hhqP3rbid5ZD4jHqlswbD1LVlswG93xy+zCZ2nmAF0hMqrI4g2Q4QSPSPIA7BvpOS5
D46dAxedw0GiPm9OsF2Mx+grHUq78s5NnFARsqmPxID/TzSnXjQFniC9GXdfPS68T5gUQwnCaKSX
KPHd6RvFsS/cFTpK0RY2uAIa+GWTyH7fHLTa7tAbKQlA1IGd4M6uswmqihp0grVz5PwedqhBo3yE
RT7B8yW36rihy3YigIevrrFYQn9QLPa+blasm6R4uAwvueUPP4K6uz1ibp51bkcaALYFuvWLodnz
SrSWNYcYI0VZChDULGMqs4SCzqenEnTjbdFK9i4vkkZ9gk6QGwHaTofNPbQ696vx/RYEWwgWFie9
z3+VJ/sIAXfsKIHgdsBBwPbJpEkwpBzifTEg4IbeStjMQvPFLOXkAegE3i3qivQ2+m8Tv6cbmZnh
P2juHbwwEddqVWmgz27KRcnbnQZ/JUcv377zHw9j3CMg/wZhHD7Enx49qS4KYrrgVrx8tv1ss/Km
qjzU/Zi/GJkHvyh0HQide22VTj0Mqs5NPSTs0MyV4M37XDYtWSIzyk3/4fIttevEtUkHxYAFio/p
sYoGL/OZb0//HHFYKrhAeHWDC1TNKEr42HTxrgrJMwyXiuDLeshL9fY7qH4qv0AiKmFXOA5IyR28
P8ajn2jlz7wVfXMuteayA6giNE081rE+MnS8DgHiQUJ/0o8odKv87DhjHNVf9/Yt9DSq8n/Vhl9E
43/1of/qWjx5mEKOUwLVSVz+XcKayWi++a4RzBCBCp6h45w9ZSTwcG9FHLbwEvBmFtYqP7hns54c
JbeBSGQQSiBOMl3rY6IVWKeoSy/QLYAR4oTzvX2DDpRnLwR+Pl/3OGfp3+n7lT5uQNtxYdPmCDOs
rq2A96PQdBScC98/NjCqzOC1O4crVyX7mHGoMGi2thoByBihZ3z8PsBHxNact0M1JOCq4/ej0iR5
UMIVeqHCwpNGt85qWYJfsiWAIZCveOS3/QQFQG8AuSGPD6DO6YQTIFlwNKSEd9COobeDFYQFc2St
tMgRCbpxsnpiQUs8ZuMILZv3K2/rrVULGgXy3UP8aH+tehSLf9fPLl/jGVNbmmxYzq7FSW60yBLn
gGYvOLpXBaScxNCoQBmXVwVXJIZZc/AfVE2r+UPoyfa2DHuzYd83WKS3CkNtVr9fCCd6a10K11MF
ul1A8+O/VX7JRfkxIF6I3NXKsMZ1w6BSCk63lvyiSfLgxz8ITWgMdhyLqvlHXezzsWvPLKMG27D4
2NA4NDhQPo+p43Abn7Xd+Yp7J/yrDxiN4BWEzVF46hGKH+0uznxlc1xObylAsmT9Ey8SKwtmGc9/
f7oTUObPQCKoKIRNj9VxKK3U96K3CPGmzF3oMbUndctiF1Lw1FZQKoVbXBGqR5IwWZXe2Lkd50aL
NQp3Y7U5DDl+4ycMt9n8yEsZOGOH3Ty0cJXjDC2FzCLcQxAnovfFcwW635KFz1Sooxj1NWBsav4O
1DKbMfSjQ/6Sk7/Xii2DzyQTVuJ7mhlL4AApaRvhO8rooBPmHM6y6/IUDjMXS6ckosnbCeAdAaXz
PAURp/Zp3jzhJ42OR0+nZs91+9/oKB1wpmK5TWsVitUKROQ4RLuxxHLJU8hH5eZokdK+fRIVFVZH
YtS/jTyn0D7zHU4lyjwihGLhkm5VZ2zu5+MzWcSwrs709UobJBAKZDWWdedC9sjV+Dbr/ndwdPmf
fOZQXQwWxvZYCvldK4GVDFF4CqLlIaA09U5KgSM86+7/sc90p7qtbT6ZpdudqXsD3Vj+0lpKOSk5
fZjJLEjESXYwKo6c6BH3pecAGM4bCAwziFWWVOQUQDeHNL69mSEgnwkBTOggLxi2MNL/Noh22f0L
rGNv6R1yqhfVRKOGN2Tlid6CEZPr5Rwv8+vtqqhpD/A/vQIyG7Ls/+rwX5/0zTiOY5CLBAZa16RA
8ilohKwi4PisBjvWLj/IE/EmNUcrdvGm64MQLOfWasdMiPSFOCe2Q06jK5iTJWr43uYpjwORkoae
i3zqiJTsqsFMdERAYATcZ7G/5CPOmsYGMAQL/xLOdUPjb1dAaRBVc1jj7lJF5D5WBuaJGz93rZH2
7PXq9XVQApLcVoaO/6P6q+CxvbcrSoqSISE/xUtrG1rrY/apHGBpg2GnHRjowxT45vm38AbROmJ3
dVHNgBuCFLRxay71Gb99vVfo0xp/bIGBXJhYbVQ5l36e1q538j3Tw9OHfy1n5M0pFGzmPVPhUlMI
hGKfxwROMg8YFjzqDShlII8fxooA2idxeqSOXHVzj2D2T7xE7MvJawxN8VURtW65IIU7WtGSF8v2
2ocqO68snSztBi/Z0DPgN0IpO6fb7RDrTzlqWrqBEye3AurTljkoW2X1UVMNUAgyoe5zrJe3E3V5
8i9cdad7KTh61QlCpXMeQptiZsllB9pzjtA0O2CT8/qpPurg1u//51sTTyH/OL9b3JdGVNig8jNq
BWDzvaFJqVxziRccNffZcUREQmULZILNrVYmgZrp8WvBz3cljrMrXAqL0UrHkiRWRcEzhH5dCjor
lzVToCn5npnPvjOT2+B6Am/5G7fqbh6To8zP8vXHtxqvcy1OmrD9qU+1MV0VXKgDXmTwgVU5Y81W
o4/qVXxCoDYa6fOso0BcJ+LzVUuYIZk7rM5hb6Yzt15i0MW9HvY+GZdMZbMxGTUL/9fzMs871+Gj
hhZCI86kCqv9FZGU0nBLxWwiI4qZqFGcHsfZnD+IHLhBTGiY7FHshHvd7uKW/uy6Z4HenQR9o8+g
bEmY2eG/8TUVS6j/gr3Onh9uxp96wrdOuxd3aE4f5Teq0M2gcZCvX/3XpCqQjVmQJO6IrvVTSBJp
11ptbNYfo5WqCAGl2utRvZRhap9Nkh5SLeVCvU8N5E2xmxA6+tGFm+9d4BnXrI4kgxImkJwolSOk
/DSk305mzNQJZGZyO5aBHsr5/J7RoloEtVrN0c5FQyCxJgKhMfLdeSITAXi2wAx5ZnPEHoNbeg+E
noidUOxtR8dNyS7tnSyXf/jcCgv6yl5VjIj6VLTXhIby1h/wQCZsXZ9O+KvwNrIta4TqgkL2cfgp
4elBNtm5RYGrukSNrsDsg3361YVXeeUrDvbYLva35QHwXdbSmYPjr2W98AqOVpgEDPjve+LGBYP5
HQu8GsbRnsSAC+Anqw7DSmX+rRpqlq08BnJBGVnMm3WvfXNhFEuHWsfoxSYTGqR8c3a3fnCYASQI
4LygeCAnD/yCOehLEtL733BgfTTbZ205jkrgw5gKV2BaDveY/qmtZ4WcuEN39W5ABQs59l1XEeui
NaFSgn16C/j9lBdK3+QQWhas5QNewnunIySnIps8fvhA3smViuuBZ1y9t5/PhuHLf/+CfSPoZHkT
IuvoV7ioSQWOXVRlqjDXfSlg4K7/0GR+PeCQfbol49du2oRuMdQqFQWAm7LX/d287VziIucAviJQ
lsinFlc1X30WPVwcnA3989Ll2G9oI3yDHO9z58NPaWshmfBbohfUUT15VfC8N9188EJ1kY1t1rvE
9oa4ay+98vi7h2oxaecZseHJwROyC1Woe0x4f+lTV86E1E2uRSh0YYq1/1wg6Au9/WKQLsFdT6Eg
1gxwHUWroQUWEL2QvEigbmZsRgWkP3QpXwxfXTkj6PLvJNRBrWFddW9Xzl+6NQu/VoSy/gTgNhv/
7atKcrADboi7e8W2e04JOovnfhgjWsZJNLByRskuD6QtGyeN5/Klwe8XG4pgnmlSR+EdivQUUBSK
ZztKU/634Y1JgGKeqYZDZVklXXQRdeGFJ8ajxa08j16CtVKfYOzfnwSHyrLQrRBiLl5pD/nrzMam
QHTLR+PIr0L5GrHltr2sqFrDEfjN9o7+WHNUa/wCxAk9V7AUcvFZYU4YaH1SpzsvBhpv73o7vwfW
+zfzshIE1hCnk+xwr1Oa32K0+5GLGfr0j6A5wiJpc6/sZ5mgF9leWsUVGgpJJ1kpRWK3NoUAJ6bH
lxDQrRpJm38nl9WPFOZqB7Bls8zh1SLHao91UjT8+BEWoa9MvokJfCyLmAclVo5rK9nfR14XaLgG
yF5SSEZOA1LiZYJG/iGELKRwhdmOE2zrzfM3lJe5mPXD5qhVGtWBYPm5mBtKc1lKeGeO2PjQ+wWj
UnvxVavQFgWHPOLze6B7zF2HAS6Y+FhaLDyEepzt2naV9b56mLpXm6CE4/OjLxGzWyBPGEft/vX0
bmr+XNkpTxQPt+wSBYU5AvQ0wgi6x7kuTF9p+H3Pe+pqLD6A7C25gtNxjrKRQLHebSa2LxD3/6av
vcqznASF/5z/tfNfZMg3Z4+FPkCc1K2KPaHIUakvLflsSefHd7/DKXfjBR5oPSjtzPj2AdKhpUtU
UrA6QY5wBVCT8Fy8zbElibyt00a04EwYB2PIt1sMbGwACyJ+OGr14kH8BsesIQIkdOGISEP0TDG7
sDTOWfBj7LwqsZEfAtB6evbu9DKbrKBa7eNRsdTxP58e2qt7TCVgn4AIWX8mNYOb/+OqGhTO7mPY
ltYMxMTOxHlsDNnHhsRVh+r6PlT5sxoJP9ikKZuNltylrNoj2TEPCDv8LRXSwqU9SXg4xid8vZmM
m3hWyde2Edor1wY8TNL+jFjezFyHnA/ejB2HOSRJtL/vxLJYPBR8+Mp9SobDlvP5ZrepIBaIW+0C
43sUztViIAZP+U05ejUOJjVSevIWJtGMJyZnSnUGP4yYj5l4FxG1/l1HXXTJGxk9xTPj2uO5fCii
vQ14ne3X9tbf3VRHy6ix+C6K9+GBwUajSXOXWOHI87A625VvRqBdavLM3hAmy+Er5Ny0WPeuuihQ
AIPugz0NUXcJdZS3S976TLR0YdnLTchPNO2Q4CJJacLRLCzEWVsdR+C7ID2i9RYUiiBHB+9FBXGS
LNHHDkESGr2sfPsl8a9j03d5b4E/rkzjy6hJhLgHKrHFP+aiEM/tpM9w2tABrCzwL8HMCGd1zNxz
em1YBTbyhDmHYRWnO/ZFlhsl9M6gYy2mwfwvWI7dw0E1BNFUYeaZsJLEV9KjF14eU98IseCQlT2Q
Onvy4QUR4H1AgeTCqtYkzCLeJYQbagIPFaUrSfMxuEGOtn8Gm6nHac2yaYhm2Rd9qV7xPp7tPNqX
Osm6Js3K8y1e5CroDqV/jd+gxAD2DJT51+aFwt7t13pyP3FO5ejO1p/NPBSJVs77j8nWAkmA+eAH
O/LJ+Hq7OieedcYYWa9xhoRhNeirHzyER7vglcyUumIm/kZGb/NKw/spDN0JWCh5NC7mGKDaNxi3
1mCUkqw4GEuyDgL3vUkYvrdl/DAQIYWiBA+NZ/dHBoHIEE/sFRLC1kCyjDcGqzdmk6IOccON0NSW
tUO6rdTaiKOOULPQ6DcNYiNfz4m2apROv/w47PVmuYAva1CQF+ySaSxsKTUOTiMlCD1fb4gZCR14
5OiPPjIe2wq5Yl1INvePXmPrBx5LJ40LWO74l8/5g38O+w6dq32hwN3sIGNodj+SAsCYL1heyson
T4kodC0/wnxWIqRSdJJSbenqlAR7ZzPyHAeyMX20Mwd0ZnNyf3Uh11wo5gUDHMm8aRDicOLIwprd
J0BVrDbQiX6i/HhpFbPtgsQm8zpwsm5PXQXIitRFJN1pk6AXxck1EAZUVtDnu2pp1Ot4pi0zzfw+
R4Sd0SXe6uV11bn8Fb5+3yfX22dtmj24dw4YZmOAov2yBsir+RhnVL4ch2f+7/n1d1r/bP84MNMa
J8WKPgaOxxNIkXyJiydGqffh1Amtza78U5EFhRknyclNpu6ZGGCdLXICA364Xd5RC8d49H9Ai4CL
eZgSMog0nDc53IWmN8ewu+uLFmV0rM0IDKwHDvVuHRq39Thao25M39YYS9FW6GkJiVcOvKhodPSw
UyiSNyPsVfs1AWLQ+IwT1s774o0TdtkgywRifQsOxqfQPolfqn5UXq9gzEg+Ayns9Ks+8UGyfPbc
RQjcMOy6g1YewIJGhqEzk3uuQpvGcHUrQ1G4ZQDaTUnHRRpKJ+8aZdChy+eV5EdC1Cbg2V62b+ls
SvnMdVZ2/NU+dr6mzYavILl/1nufWGhrSLSt7vLz3ZXuD7FoRUstZWmtS6dqXoeKrAHqRBfdkRpC
/hG5URGqkXVPk+LKMt4TNJEJcWe1DfY7BZb5VvOY8diCI1viLYLvBlTYrsiksW+WPTFl4oKx3kVt
nIgjhAv/mMcDyVO8NtCMpOrB+6XpBPV2vwyRD8aWXykxAghgTwAWmXU14IDif/ORRXiEpKGnZUT8
N4miGeD7Fw1WEn+A+whoNd+OY1owV/sDsWo1hgWpgA4yQ3H8uZlh6DdKx1oNPDMwRAY4RWAshlO6
2cr0WPEE3XuCkuMYIzCLX5FBU2V4eHmTKw8l9pnXPUGAhNgdZu1gUlKxUsrxXYqXucoUyNiccbiw
9lWG/2cQnN+VI52DcoRrq2YxB6NPGyQelkd2n+KAESTm8ZhISBORdsi/WaQjIg0nZl6BxVzBgA/J
s/EjfsnRKjKhLWmqdrdJhuzKMhilod/1S58XyTnuAnu3RS2vphQU8cc6goOtUVGrz4WZfhXP3zBb
R8nJxMyi6lreYUgqyWhQgrWM0a7OOCuGw+bJJRh97gFKLS52m419d7hkyohWsxstYpKjRPCZtNRd
6H+KgCY4kvptljd/dBmkXVwR0ATXsz+qMwKRbm8amgM+ycbqwXz46YIEEI4wXEaxRFs7mNgwCRNn
7HDDzy/Y2A3eOM4rFrvISz8BFjl/5wTXKPhIyMH1x/CyGfUZ7FrJ1FmawvjC4rKx+Y14GAIeho9S
XR809CducnYA0ME6WsLb8IfFkaD9LevH98SsO90PudDPr683apVSNgjuuXtThas1PqYrtwSSOcAu
D+y1fpWH5I58AQpUEMzdN+r5wj5QkHSD1tgYulGvqh/Ks8/nAqHie1+fT7b5w2q/0GDsdtFrQv5w
rpgPOodFrEyyAUDhav7g3OKUxWgZAhKZyYKBJbDDqfWs2QEQkpLsrTRMSt4NMyiyxMTuXIfDqRTL
HXC7mjKsNdIbXEkOjCz18juxTD0d6NJSAH5VKkwHiDgC+etykpbWIFH74que+CwcEIFMtvDr77nj
oTvIgPwIVq+1OTkQEQppUlimEJ8gVdjsvlrvxSRD9VzetQVKaGKlSTYrOIj80XQePbdZ9kJLW11c
i57HPXH/C4Lc4jc1SYnZoYn4YZQlt0qcA1RfeDViFx+fW2nEr2lEwX7EzBg9HpPFbNegl2OYUTdh
gCB7/qskPm+u+YucnX+GY6qeEbwhbaZkCfhL0DTp+FBb9FvIssPy5eWo+S0ykcl6ziRL0vgB0kt/
0HCbZytnBmnBCkvPGDMad9C7FjGxz7buMzxsPKaV5lSKwra+Ggg5k6QwxP/9L9cfN93OGFatiQD/
7VQR5kZJnc5qUqZtxHR82lwV+yKk84M6vnNIDa27eSTLwZr22iaIveXA/Rp0UXVy0hLYdH2feeqz
cInROAqSIbDngHNjdBirHSw4IBeszdXIV8sjd3pONNsj87TcxODS1SjevCNuSohglLGFy9JeQ46W
2ANEuFz63TmgJz/ZL4q9j6+bL59eig6rHdq1DxMuvJrrGjVCt8RTcLh58lxARoca3XqH1veWQr3p
+ckX/3aTYcN7EtwFeKm5DN3lIcef6Go9oFrb6TjM+gNy2wgIoJNhshbClT3r6GkLBUfPzEEapNc/
qd489mQkCRJReIfK2tlq+ZKH3C3eDHFAdNt5rNQ3R+j9S4s1AUVqwd28TVgcr7c38dybqO0905R/
abrrugwVOuRk5K9DQg2YFaSGw23L/gxyP+dlpXu2pJs/68ddiru5cxTWIS0/cFHrDofHif+wwC32
xF5LmqlAEdttxHe4Cz0AlwLSgtMiqUS1dUOdRmHwRIoce2205C9Pouy5dbWHirvNUG6yjdz31iWV
Fal1TBaVJukxeYbHGZhMp9hTz+4CUjOhryI5O8Crm4j5frPw5Nwe5E4moDv+hznVH71k4OvfOOxk
4AfYKaKkB79+DMDEw5SrGT/1/xoPW5hPVLz2Myj/RAAT5SupAEiGCkpGwOCFhD0ONec9by6IVMrF
HRViPy7HD2No6i66DHXbypAKm0dSaCUDXMbMRReJ5mTZSOzTgoVT0VjUDBEiA5o/NngkXgaQYvtC
/Yn7G974kDO5rvWJJz2Y84n1Dc5ArFgD0LDUOm5dZqMOURGN/hHHLXTU8dOMDJnzIK6wjb8BSwmW
8u7ZqnDsDBPRj9wiezOn7xHBfkQQUVdZ/hnKCrfkyVoQqOYWeR5o3DJ//RvzuCjI33bnlFTaNajF
XHds0u+r7o2lAWrZeKzlxKjpYeCtsGzn1/VVFRysHR8vswwGQ6pDxIZjcy6Y7W9suNF4hGaVSXCL
Cx8dIv/KhCGhOLROZSTWb0E3e4VHPp2aL7kTBczPd2aojlCHniVo9MYLO8E3R4MH1lONknfJRov5
yUJEgca8iMOTeg6A8ilRtzu1Ax7qobSKPzDLpGtKX9MsxOfKyiqJh5PHOV1gqVV9upKjLRkXDzqi
9FAxayigdZkQbQ8AV9jPYTQxPlnl4S0nk8hcKOFFRlTLiAzem53jDwlsZUhAknctueUDAMKv6UIo
QO/452wQSmIQEKheIEiOTBO7nu0VFCDiVf2P3Tbp83vXrlMTcpG2Y9HHouFfYrAT2H1YAeGBGVzM
U9C+T8GJrHnk1LqEtmLnwhybPPpKGFUYkKBxSPp3qzI0RJGAUAMGonMyLABxccAuCB8mHxREAZPc
tf/A52BmljOZruFNNjaevU0j8MF38LNkHR2F/YVbTtJqmq1qAGu63SIUMpxIyxoOlkgClBYQP1jV
DIC6wV1or/vt2smh+rp9BZxRRHCg9tzOHMGbF/zuEg0G3959zSc84jw8pqkw5qfoe2Jsb+jf7r0N
j1d72e6L2AuVzUWK6JAccK7wNztFTjbQ4E4BCHftXZl4TJDCy2eQxUOhlb0y9HjveOHFaEXN/F1A
Gp/F0OFVpEy7FX1BYtZA8JRIoJMeStm7tCHRERPSk0CmxiUR276JbuhXqGqfV33eUnJo0QTLABkL
4QTT86uqlEzxjgbdukT+uWf6bpIwBMuj4DwjV/HeN6rmCXdWtPjUdZ1KPHQk6PuLJrBoIzOxEDEo
V/uomCjA4fHYZ4k3W72eOw8sNxP5CojfryidbL4TrruUiMmFV+bZIQoH0sw/zCwWEFaN+NG37x5M
3MelpF8lhKY5eSfAagb5orBD4oVazeAjXEy1ggJ9YOwGmRYtxctkwlLYhUpg8PP3mwFjMPmu+rtg
DX5ZM+XOhoBc1xK0TJX+iLFeAx1G0IurjP8Tovlww/kU4PIVIS16VySdw/DMkvK8dRMfn7xUD17g
PJx53uR4VByhOwCWE10WyTWNkdyKMHGcLAY5ElVheQdHmOyMCT0AEwERSJ0jhyWeOkJ48URvKfKQ
qqERGzG+rRDRD2IC0pFEeDoit7eY9tA/Ktyz+2wyHpA8EaoeFwCO/kqaP5PlvrWzxh9hk49Jzfax
eZ7jqNgmVfqeNrX9+BVLsIUzYj85NEnvVp6IwJTkR04Rb70my/TbpHimyxVpZqXAfPSPzd2cZEQK
o4obO6cCvOEGgKk3fV31AGNgz6Zs7NPewLMe4NqP6doa7LKM+/ktmjp0oyTID0V5C3ONVgt0tYOJ
u99faH9uy3ullaHILlVQGHHRTxgQ8sydw7fDJLD1uLwzXhdHFKd/gCCXjrAxQ1iLOeQz02dS059z
VPiAYbNuyD50Sbf/qEPuY7502CNme3r9OYedAzWmEUKcIU92bg5R7Qtc3/w9JFDPQC0BpE2WEzWx
xxQB2jFSL5Jw2Rt5B4VjxVc2HBiaqj18tphjlOfmxWrySAJ0MNmG5gsJWJzOQ0zQJbyH8VGA6ECc
fccDEKiJN8vlUhy+wcvHNGv5wwlepH5cYtKO5PHOL+zp1NnREPbpX99NY+J+KMh9u4ql0OXRukAP
dGFjOw29q+tpyRpsSFTpoKg+cv5eGX+7+qN0BilxSj6y6u3LA8X+gy5b5lQ0wiE3DKlmoYNRd2/L
B3Hu1T1/8Ef9jCNMqp/1o75lDV0mEuaN+pFItGfrrHVkDF5/Fy/Qtbro6/VSy2qyXFuEmy8OpwWo
UNp9reNl9S3IN5KiEFc6cf/KxNN9WKzcwCTb9J2OpyxnlbqDpO1jJ0uxf1ZVaQlIXlkkm2B8jC7v
X44xZwLR18APcgy9n/yKjL9zJ05amQN47OmM4q0TvcDP6+Sje2A8+/fA2XtdxTYiYscTvlbF2tJU
lZyyql2CazkHl8IDfWP6hZP2LDyYw/ZlPwKrhvhUi1hUglwr9gspqRWn6Lyr6qLv7VZUjtumEKx+
CDSfMm/D1Yj9e0wx23C/ydsEyruH7klhCWyyrKkw/AuKuImm/+Uht8lA9XTNmqQlwTISip2BWtBF
NgYakbijf3yBd5Z+fG91YPbSLj+3GU/tSG8ojNzByBykkwcxmwuUDhpWFrn3lCoC+OKJDPAXldS/
sZ4SJkrh7NWNGpxpFH1b6BoKLti3KMw8xJYvEgVl2SLNReNj2PBFMbEQGhHBXc2J8U0XR83VVadR
vRWP4pRgbI1W6v9vcNnlM1LBmrF4V0BMOG/qZhJK8Veh+ku24MUkBL7h3/x1tTW0a2fFTwGeGjps
Tj+kHR6VGiUPuDhi342vZXUNEU7ubk4GcoWzCiyCr5ll4M8fwEZyWNd1hPGP7loepuLx9UhlF5wb
VIh7nh/efPBC0rbhUOBOybN+bSxNbjS7LSoXcdWYC6KlnKc65IX/8WUfM2ZxYoBIerr1KlCp5cAE
YMAf5hg+fh0UVk8BywtHXV2yCJhfxf1S/cgrRsoEyn+1eHo0a2Rj4KNhh61Y2NBI+7dQf2Fw0uv1
pRSSyMaoarSRz064t+3KsMdfjMRZO2vc/VEwiEAEj0Oi+tFPvGiqLbSSGMqmircn4XlSzMzGDSA0
YIs+BIkA3pbrqVhOfIYj1yPirEqlK5CvqdM+0cQIQQzSpeE57hRFdNMF1jsyQWS0xNb6LrSZbDy7
eXKV0LNERFI1JQauA9u+SFaVJqSFvJsPlV5IGuewKPm8oCyK7vnGFaTgW+XJte0cPEFRQvSsvloM
7xazcJhtbmeFsNlqi4TSmz+DEkA5mIbO5WWGy/QNxaUgvIsAdn6zCwApeM8nounNno5/3tBlAEU/
pD9AYaELVQ3TV0vDtC9TW2DCYfF8hkGzbAyQDeo1M0k6cpSo8Us0mEGf/kLIDAQyk27fPyaGRdLb
4f5rkk71pc2Ty80VAKAZ2Q6wJLUNZV3UT4d/JRKBkXyjG56VeaWBaD/wJTrozQ3JGPNuj6Nde5rI
SRfPurE9dwaahSYadzTtPC2EXpfJkMRp8u6XZDDkoY82EJf81ivsuTWnKS9BXVHpkEtSpEh6w4Op
tW4MQZwqFApJn4jKMDHon76L4Dt+HhJvECRNY0WytAPv/p2nBV4LMrbp9Q8WwZ4lALhpHa08G/ZD
MmL9qtsEGOoFRDTPN+fS0Xrfyg1wk/nGIxLcE01+EZYiAfY9AEfRr9a6dntwmuDD/6eg8BqbNtYL
nyvmgJH+1LxdS//L4NVbIdkXI3u0V9jJ8o5jw0lLH2Ny/2hZ43no4cFSo2f66+pvhJy7k5Fyk0Fl
eEAL6P7lzssi0COYSF/Yl4axlEZkNVxR5ePJUAB7cNhOEzdKcipzJLAI6YEoh6IbQ1FEByMOLoaI
HB1NiQW+kLK1fg+2GxkPpOA/MwN4ax60cy7E0BzvX6B/sQ+RmJvSKWUh0JroipSTd1yeL9q1lWtR
ukZ37t3vnukY5FOzK4K7t2PkFKfqWgfQeSunIvAWuZL02Rd4qrhEODi1BvstmD0KVLKqy4iub2mj
8IjLKwS0OnLIv7UsVgGLTU78LGIdMiPqndFVDOBq2vBM5a8U6J3bAnc7bTtQygu3HYCNPEq192RK
uxUrmSxrfwa2sSiaGmwnO/hr7+0WRnhcGL+8wgmQxb64A+C6uzQy9fyC3/QnTmT2WbU0aqkaBWXa
ARWTJO+e1pHe6EYb/x3TXbQoJz5t+ovJfTxkr9ndS7dE9E/Jg+nvyE2ZipUjbDkAOCY+OgdX2rs0
0+VuuHiKy2+AwEeivjIiaD+I2+4u6zVPelzLgqh+iUKy+LixAWk1p4XW3I4YvEQu5czEZ86TImLy
bNn8aspXq9D54r0e+8P171B3qgR5QdE8Ckzt2cE8Uq0EnpQlEW0y159Xzz0cwNtvb33dzFg1n3Nx
bbGGVa8M5ZNp+65rX/Av/M2IMZ4E7k2JVCNEsWMsI20ON3gkifetPn5CzsvL/UH52o3y49w+l5ZY
43oTa/wILsPdCQN9uZM75OXXshgRAdkVniL9rkA/racD1CkEinzxtDdAD+76XnQsITnXqT1NIpEL
XSebR43DZ1omzE40hhRwBcg690j49kcX2IPBtVjp7/MxOS4c9roVr2e/BlzSmtho/EHoqitldgOD
QxbNfpOnyYCXDo8uZoklIIYcWfP8QAlaSkQSUuyBXN7WwVypOgn/MAmxSSnQ2LfyP26MOxcMv7hT
cjAnoiZpEGBgmWAdAuYXtQ7r7uNRI6wZzH4mBL2IEScpVQEbcDj9chcztb3xVj4XgeeXFgcW0QSo
Xt91mz9co6+SttGJnCuO31q5um5sujkHZn+zkfBDcPOw1EqqEEdUzsZ+IWZXseWS/d5mVWNSvuTP
NI+y3pXI4gJylPLPwjWTAeCZpDh6yTdGiVTyg5xEx08QSPOT0gPeBgHJrFZf7wqcdKjerdhgKhCq
t1G+nYUcItfQMUy7hR2LY7Poh8O68rmTRrdbl2wb3GdvcgOcN/eM2OGltxROsnTZ73caoa11F2Pn
kRCa8jr2nne4ICNgZep1iji0uYUOgFGcZW/FeO9/imipd00m3zb6jA6a1hW4avCx7LpA/+NSZmRg
idgKfTvXZbwcppGzRBVoSEbuNKLB5y9s0p6PdD9NG9PuUMnvxLPy74ATmKbO158063iyRkBckyAw
p5DFBd0Tp2r04aJRnBJ/PTw5/a5p1kq6NXILbQw/cfyn08qY2vITMvDdK0V3nCW+wc6Qse+pywLe
56IXrgP8SQAd8/sw6AqpXevyZKRVTIiizAjupkS2yhgwZyq/jn2eUOhzJfsJBiMDK+5v+UGQMRRx
48idt8rF54fyErEmH7PNXMKcZhwbrs2wOpLzRHu/b3+rExhUpq4GJr9pwaBucqpd7kx2r0U9p2KW
drCx67IL644P4PsaYfDrL49pX8xV7iKP4Tgt50tj5BVqDJ5e7dINEjhrNQ5/zHErdVDWXZtmf7Im
96egvSvjkuacTROavVIB2X+c0z2VdjQ8JdHkTaj1OWil9S6yZWPMPAwOtxeUlHv6IXcM6JRgOjRR
NVG4M+Fhz+3RC8IUSL3quiz8JJ/9JT4H3uE8TPvC0oWeu9ztD26mjSviSox+/gSd3VvKNZPfD4Jx
/Gksa155H1TGCgYZgK5OHcDvB+N3yNHyiN3H5rIKhn8wp/q/5X1QI2aLXWIfVN2HZfUhoi2WEeYW
MGSR1pEvaRaA5HYpGEbcHpt9hTznu+GUB2/FhWddeUQGDlfnt7GtIDCCDbtNo1H3/zLdetwW4Moe
P67r7KOQ/lA7mSlZox+WrS3l2cNJvSjCltd3jdSo9Pko0h+bLgH3zKhHuEKVDj95pJGQb5jrrz4k
inIpa8unEVyG1LKa34kbb2rCP/ClMKLdvp+fZsM5uQydVn1CJcCW6DYJjZ61t4JfvVzOUt/tamMS
nZ792HtqJF7JQdoESJyCPq2hwxZjQVND63UPOjBJUMOYRbQ0ByOUAhkE5H5F0lHt7OSnMzvoDINE
fM8eyHkfyntRe0c3vEL9BK71X4zFJK7DN37uVMoGqM3hXkALL938ThoR0yTqAi6KUqv8mgijqJNc
e6yQFwqlgpUG3Csm446qPdCsvGJixv76AhVu12ENK+EaP8TeT4bVt28VDQtKIBb0Xu9+vLXnFntl
FDMsCJsn/Xks4hh0JKYF2a6e23OHU5+jg4kHDNAwebVFlHyZlxCREeZAxSvumtzTj24gEmoQQs02
aUJYkhtu69CmvNuxSRZRcaxc7RvS4G81PntxmIbWRz5aNV0YpjeGYc3B8PayAfPq9ggKJQjRejaA
ynZuwaMgGkOaMdMNqSepowohfzDS67Mn1xqaW2EvIvdk/lcitKHeeutp2qTTfaSoX/sOiWPsIGrU
OHUiuqH+uvBWQs1sC2+jrVDV+rIsfW4WleiSvaYpOA0uSUni5+g/Qxr0c9Gmx+35dq5fFPCzuJ+v
SaIuW+zN/mvEfDvhpJMzvShN48OHe1ZIwqCzfHeWdflPuxAUrDroCHXBrTQ7vvM4GzRr4R05Hl0e
mYJnAFKzLNsXTyz6obJpKBlsddTifEXR33EX+g2N8g+qjvJuSOl5yme23rY0THEjB6YNEO84kRMu
z4zAsJgwNP/ZXJMxmYNVXt1PRD89uOyT1EeTjD8ugzTeX6wi2VIxhJXiEkzuJV0ecGyr+MiQAikY
62Pr1w8qMeBUwAywqJPv7YMz53O3LKWo/yZGYcjQjMplmXUbCiOEsC0k9GIRq3GyNXAolYw6fTD5
7Nud5nt20uYpvpF0aH/8tsXjxBHniOBn8iREmVUpcHmdWFSj2LgeNeuPT2oBT0zDEDYx4AIHRG1k
GQhhh7Fh3zaIbyMBTxr6u7zcLYUedVX5pLN71ZDpFa6Z3jAonh/yLgYVhdfzu51VFu/LUpPgeQkb
UtwL+KGwr1vL/EFYtAatINFyFiiALCC2WgpMuSpCO8kmI4I/zA1bHiK/uFOwIyOlXFWE0ZypQCsc
FgtRjSOlSJXi/G73PdAsuO6RfveaxQm6/gXWtDrMxiEuCHFW8UQJS8xwkE3Fhzq/abP8v1NdLT+5
qD6XFhHG/M+ujCN9eOzGLvaAAxRFd+0dVWPFYLrBj4Gt0kPk2RkV7/jh894gsazrcxezxKg6FNwr
ySZjNStN4vzusXcXTDYH50EVe7uNRAMAJtHdMwmTgjsnCF50MTb4kiC5YwvU+xBdRVqB/QowuRJY
aahOGhuwBZDr8xAY7tytumj19RLo6NT13YlPa7VVsfGyG5nBmMBU2R0lj1DBW9J80IWQa5fvqdmU
NcGQZZb3CPBu5uFfqa5UeTkA+5IJanEgIyPt0m9fPhxw7H5CL/lCL6xIa9+tBUAyOg/7MxQQidwr
kkGno78rk2ZLKV+HqTm0T8zfVaiP9hKlBuXz20orptBdpwPNCQjoICwYx65Wy2rNTXRYO68gWLqt
AAjjGkjnrQUDIoLM37A9gyB2WjMKD10YWNaPled9xJxmEiJ5Pd/pDJGH3iJTbMuOyCLpCADTUAa5
3Oc2ozBcClzEIi0UdVe2iQ18zauAifiaoN4uGCoDrXbZsJZ3ZikP8iLd8xTJ/W2fl7NGzsSpE+mw
Vrh5cioelk9XXN01OtKO4AU/O4dvUC7VOCcsYEtNY9m20pvfH2tNCbvSRMJDr8PcGcIyJJVYDbyK
qh20TPO/S3GFNWf+YnR3HY6fgXm8lFkIoiDLPXcZISEDXy9W/RxTBRH/RXAmTaPFxpej6C6JtorR
A8IZJcFpxribCFGQEH4LV2meENyrEPhBobRTRKT7lOm8FyteSf4gIGj2kt+O9b66IfT/JGghh4Cq
LoE3KAuZDOXZQwoL0j7Hpkz6qmDH9WVzrBGHr24GJFm6Vo0xTZZJpYtNvwG5SD8gY5Ir0UJJhn+r
VQ8wxK+K1+LYXJzqc9ssCTk+FeDUltT+zhHnl42uF51c8Cn2hnCW7dlQISl2+vgXfhq3soL1bt5I
7IRTo0HORq/X4UjKxAmFk+JVVyDZdW/0kRbpG761mhP1RWVCbpdc1s8SgxI/PWrgdnpWOtenfWUh
AbQSEWUIPuK/D6/Axpg5O+dKCAEqFQPzt30hiJ0QYqLMbxFsCBOpywGo7rbSdVPd+CtLTL5GwTR+
bAi0T8Vq6UlX+hWb528q4X59oOWU35OTicjt5My9Uy0c2EIiYBsScRicUJNOEPZT3uWZwjoF1Eyf
ifrh8X36sJe1Iu05WHuBMjDg4oFz2DnauBE7Q9Pu/zjP98L/si/ia9AFXE6lK5A5PxvxL0NlfbuX
wbbO3pyGJQVHBcC152NfwI19p5X/xVZNwizsksICmlM3Ya56d14e2+ITfY7GJdoIELq4pvJqvzLI
z+b4AqnFHvx0BQIEWLMjOFXSQ5jmj4Y6eygkKXsmE1Cp5gOmnLwOdE2Q08FsT6FQBLi9FuMxHKfN
Pc/z09ZCm4MshPSA03bONY22fzjW6ok2KMJZeNPvuVQziAuRnN9gjoe10lyI/s5BzCwqF0mmit2y
KjVSJZlrJZwUIxQ0qbFI9tR8y6LPdgDhP+BdvE4GV9aetuF8ZOe+Rsh2oL+kdqlyqLQtiug/SS4l
SLekoDoz7h/dB59l55qErCdKa8Mkq8kfcIwi2V6VE42jlOi2A55Az4Y5W1QDxHQblVO/DXPNi0AI
1XavG1Z2sqRjWbDS3uDjxTnqonV3GITX4X/IECFhetooC9i4GPZAWJ0xsjx/sqtQDYkIEx+6eVaE
ayX/WGz62dxbkhyQmvYrI1jueGDQAW13TlyJG91H2JWV5gcSzLK+lGTCvd+UC0GSZM677lLRTh5n
GioDvFS2JPlF1pllHRFGVTNvAcHiYNmo63TMO9clytj1RfxwYWYouraLsfHwJ5CRoEHyOTLoUT9/
zAEhJU3PMPPr42SHXz6F0j65+MpjbHS366YTpKIGv1xm4bLex6mgrJdK7h186HA359WRCQhfaPZR
OYltwo9/i2xkaZ4wQu4pHr4wveyzfwZw4KMxlVj0RiXvZfEguh1Y36ovrvh+RbopL0PzE424ERzY
5QDPrchKh3D7HbuDgu57oaCTpZWiQLYAFZ0v1cZ/emMrOW7wMMYNR5EOkJrTcJ8IPJrgBsxQrywd
f3oIHqfLicKb8kwG7I10w6CtE8Dkfi2DzkA6eDwiX9wH8hSHdIah93Z5w8Ftzy2gz3zQhJdaYOmr
Yus+RJJwbNUY/uxLGeJTclJc/cIToa6FkAnhXhH9uD0p3Z900pOwhWnNnvDIvLQXriBiljo9ofhh
oxsDOVKbH7ViBFamx7lR96938l0a8N9i8qhiqJwjvfF2A62AO/S1UKLp9mvu2/BFWnzWzP2S07kW
IJ6qQE38vp9u7DrHzgFah1LZla+GKySRL/36eTF2TCqQKl6YUxZAWJhuGf7DeWnxlXyHmo8T50Fw
sFkyLeWWX5f1p6944eDHE916jVXf2C2jZ9W25JSPN9BwYwDYn5Zp+3IRxkm/4ZDU7himYHMl16n+
5YQNrt/LyM0VwutMXcaNanWzfvEpZj6HtYzx2CRDwuAFqaxQYGPjYVNwYp857KUsfEZU/dbIZ8we
xlPLsPORE7Vbxkp/SLQjqrRDIGK8/sz3tRD5nHOEPkNuCKRJ+M/4mnf30uxM3vehvfELzHgEnqJu
CQBUgDZu3B0miz+oQs7rnQTnROftCKntnO+H/cS2EjMS7Me0iw1YykeEKroH2X0zBLj0zQOMRsMv
P3vFXth0bXG5G8+qpCJDxKZPMb7uV0qOiC2Tf/2f2Zs/PthD+LRexIEGTBWavH8YvB1AZHD3vn63
ohfqw8SEYq3XuzpDia/ihwpl0dYF3xIMh+pwBtlOe0juxgZ95qwPCuuAhnykkYi+Y5HkiCaSu84j
Ori7Q1gjDmEoR8xpYxb3IDH8nHoDY4rTDZ8t9ontqsM7EdSvC6O1xux6DvffmMlsV7Bqrstlcovk
eDHOalHjZ6Ufr5gdL/EcumZLQSwHvwFZmZlEhJED5koHmvwbYn/PS06O5f1e+duhs3IG6LLtc0ts
Aj7DEaJ/UVzs1kATmQvDJdJxT1Vn+NY/aJZ5gcSCEWSMHW36JRWlXK60Rv/Ouzy0SZc56Ag49F3H
PS3W1rx+HFMSxewef51cP6FAJ02Gt9zwdhci+6ziP4UL7z1DhBuQoIi4KfPUWoRmmbXNaTimhLbt
YFa+40DWDTtTr78ZB7F3D00y3lb5WuO/4+S8F6Ol4yUTpVHSt4khJHMytpRFYc9XfzqUsqzGThOC
eX5WICMpLnqN63Sghh/SOuiov16OUfYBJ7RgQBdyo30YyLt8z38lQIhqGGe1jHtND1ILhFlZYDwZ
0+xnxRkVF/5ItLY/PfnS4quN5kI2X9IhnJfQBGe680JI/ehdBwgcmIrgWBdiae2vy1pA2ssoi67J
FbaMLnS5Td911gFqJN1eR7QjOykIr7TyNNI5CI5njbvaKDMfNFqhk7P9L7Y5sshoYb6gvsUqvn0a
x/6nHUXP/c0z0eF/N5kA2xQ5V2ad9uiBDoDVQoz3iukv7MtkCWxoTagsx7Q4jly6FI0bhs3xmm53
zLnrbXiYFWnYegFVKmvGRx2gY78YSSCzwJsWjru0ycpc1ZwvvgCj9lltNj2OzZ0nsJVthEmnn1wM
753evdk4k+KViUCsh1Bm/FfSszAW4GkIKDYCZacW+utOda8qxKdy2e5gFBCXuC98epwTCP1HGq7V
Ip+mHXZrC4HmstxGQjBV/cNlDrwz/tAhl/nm4AzN73c8aZe7d4Sor1/Xbv5LM1d7YeCWVQkQD3Py
yzX95CvM5txmL3r+mFt14EIDlQBxUYFFE4+el/ZBprH2qWjyWuKexjbjJ69Teg8bn4tVgn2/6lcY
gcKSAnwEoRFWcN1Ndx703e/1DYdJCGPSLBaXQY8lAcM99VKfIWmfZfNrSavUoqhhE48h74TdjK5p
EGXrD009/x3C4s2lLA3wZym+GdFxums/7l269BZZ7ZJPqt8bxPKyBW/tUN3LFCAlqLXTrT5cd4Cm
FbLEL4F4RvaiSfpUlYjh/dMMHUqnrNmmV7xeGfB7yKxeaB3MuxC/kChj1TZfkws39AgLMdViKUwe
3xIbulolnwhZ5y3uwz5gY1Yo6txpDGMVHN8+4ITk9s37o/xmLJ7DbalbDotWS9E6gxKSAVRxK3jy
O/2cSYBoeLi01OYjoCstBEJDBTlbFsWkME6HKbQZJVflwRQFf0vKAKtZxDJy+wldGED9op04YdC+
CuALedAXYF6/zG+BVSRe4sRfI09v68M2swUNIXWwGi82dia3fSuLKyxx+nPR5h44w9g7ZOhIhKwo
0npd60+6s9qiOzZAasBBdemIxniWVQu3pDTDjtO1X2Ut/GUi4Xz09OTJbAlwm6MXsdtlJj7xQRU2
MPc5uEhJdUmir3GYyvKkEz1u41jIp+fFhhuTgvzJ0aq96tMjCAOJXqXag7HxrFFzjVPUHQrAcgeA
xXIcB8Yf4TFCcSCjYRtia5Hjng0g48PbwcQPeO/dgCsRl9lb95H/ntdFpfDCAyBvuwhCdy3EVXea
TO3G8bz5hs4wOPCh7s/kQaONGwilomj1QucbesJJl7kINWTa2lGPvUAiRlMfBGmUPM9MSVrNQE+s
gWgWW3fjzdo3SWJF2ST47CmZcrnn111+sVjqbylastH4dPXT6o23a9XZBp0PnLjt3qVi/icdoHSp
yZhMmsdrKVtPNTF/yr9yMGAhbDKVcW10rTWAhNohQ98F/yK3CaeqZn5j77JaGBFu1bNLr2M3mn96
bnXrkQ6U/x3s7IjhOtkeV6cVNNEe6VMMFjnpqwz1TWddwK1nbpLtfZIarGgy49k+SKqgxuc6EpXe
GPYuXh28bKnURBhw/PL0poY0CTdsAN+Uh6/fcEP+WYgkMVno4A8CpWx+yXwa55S39isWAxcwUWnc
LCAlA+Gj9HIZOjbXH/+A1rd4WBU0BhyaWu83ry0Z0bIkxfI3WryxHmh1vCAc+hThhaiLCphemklt
pD3k+hK4ajFxVIj5gO5YjYKAh2gcNgcZb6k05YH3H7vByzWT1BSZvnk+eYyXNsfsXDAbgdmeOPaI
/lMoNziZO3VFfxgGJwI5s3XuwCbywkXuyS0wgc37EXLQm/3D5nGeiAc/ci8nmaBESqwIS6+yuw2B
welb+d3NXAJLglnYj6J1JzSiy8bm6iLQucrWtW+cIMYLovGKmTzPvilE9G6RoUi0NjU6BumOf3FX
/rVwdLWuGbkHH5i2/Nv8slSgOdsFbJKQLaEaJdQBVZitpHBPz59+zZ9wmWFM2BvKglPwOuCQB7TH
3TBe1O8pi6LYwdULV9/hal6hTQvkMOhHmj8bayQgRJmoNhCNzMx67qE8DoLBlLgeRMIHAGnizv6S
HyQmhzySue8TKvF9V9wzcFqKN7VkZT88Fn/9gVvFpab+29qMJgHl8Z3wpNSY06z+bqr1g+e9zTiu
fXrUsQGmqC9QgI0ppIujZldoNx95LFkHxDE8Jn/JVLUijzR7y15Am95icf/+QfyKZ7khilt6n+GC
Nr1gg2DDTC7qHWi7m3kG4VyHzDXK4vZTXaQojh/Uz6jCCIasCpgMl0nwo/fLDT396p/NQYcuvJwN
LJYrkyOnn/tiwUpAQHKrSIuSlSEALf1ZOethtoQ4DK34MVeUiqNNYR5tnJBuyGjO1QtS7tTIRaea
A9ylPjKMXmWzQ4aqZg0YBVfLrnqGVL8QqUIxQQNb8ygeWIpOuq6WTwCtTwPOHUd6OHnVyaBB+hpR
80zP8z9k2WVcBKHBZ1bymsnv423TKA5TOdVTkT0Vq/sEk4LxlgH/mm0ZehKU7GnSPXkeoV//DlOn
faI6fAyHnOm+hsltDiKcAmZaprLueuZ3Z8EBxlBIIWQLhXMe2wUmS4pJBFKMnJDwmnNzTJlVfnhS
PentCfgzGqGD2jeJN+ttdAKcPrljgmYSBsVocfvn3hFT0e89yPWnwPmG6w1F5yiYyfXoKr7yAt8n
O63d0YIJVz7GO4AG0Yql6qT+OhuD+zW2Je3nhw4mpdoy/+2EvXQ01sSywMcyPbUb2mMCh5TlKCWd
AkLrSNLPbnI51D/uGt1hJOfy67YxngdORHgpoQu7dKiVgFdOuLDFjSu+UIN+Mw+qxAEwJCZmRSIQ
R2IC7KnRiEpvCPy7Fxk0qVtw+2kP/NDzPus3UxaDnv5xQfCUo3sAbIU/Na1j+bRGb0OPNx8nC7+U
cuqW3FZZ4ytTt6a2sGlxHG8gBTdqfAjjwc4W/4w3+63TIH6lu5pgyE9SqUuvG1SBDcrD6opuGX3l
wBUVJ0ed7Uoob9dvGPqKQ7Y46JB+Qv1r+90rqmmHb4IiJa8oXdBvCftEcgLlYDeOW4asrv5JUJpL
IPxf0dBgBTFU876R5lL3E85skXbRjfyFx2IiXR7AGSluWT5WXLs8hvMm0Ii8C4NxM1zFQmt43wU3
ZS2r8KjFpPMq6LOF+SjVV0GY+HWznx0zf9yQXbHEuX8q2UUi72z4IOcOXE9R5AVDJkX0idKb+1/e
EVCDFA1qbRQjHwqxT69XF/5NFugtVXxMkevoU7cTLH3ZfvBZg+LaMGA9CQkdBo7UhXI9kHaktLLM
tCFLPdFLxhbLUZoLWP6s6Z0nD9dL2rSwEOO8MnY8ltq0LdFxQj8vAofAaPpVeaCvRLaejMfHVz4n
f+PSAF2ia+6gDfk+br7PTfsXVmr9RoPOogTQwXa1fsu374wUtgFewIaY7WXpZ7E8VTbjiPmLAsGE
hwm0qv7zN6WJbZSHoRHAC+2SzsByZWo02wHMZVhYvgdSubD1djrhAjvLeATKXCgKrDoB7HsjNiWC
Is87pYwRKv8CqGdMiSuTlQU10EZNerjlMHPTygJ/evisvLmm4gqyA0Dlc3CJMZZmjWLFMZ2seKkA
UlX7n1dy/MIKP1UYrs80goGbHnywV3f+a0qdjNWhRPdYhd0Tb8LKegk3QVOPZiarF9j22HCIQW0c
8sSd7YpNqIJF46I7b4hBmkwx17SP2izW1Zr9W7ib9gfAaIu1rOSKddHV2koCe5JQ5WibSY3a+H7U
xVU4qnufaIyRJtQx5FfL01MCrsoLBvpdmfWzcKHHcyRmCJxpRvn3Px8ptaf4I6X79E/nTImx1nB/
ZHoZ/W9OahEdSGTxzAu5UyP+fH9fPmKomsYWiaz5RDI16X5gJW7+Ok3xqAR9rRi8wjXjFR1baP+1
5zLW8WabIWu3LWmZEZv5UdVxywFI+92Yi4U19LIHDGbgAlDS1q5SPTxUn/nTFVO54FTeWlXx0Tym
zC/q1G68MZ8TcIIttUSH55grA7LV2z32JAcJxJ0WE3wZH8Z+7MRZ9j6pxa+zpQH/bse0S9FUVe6c
8ELlAZ6GVLrh+CLdah59H+TTI+aATdszSqeybh1O08gU1pRkOYqbjhwWoCN3BFdzv5wPzCtW1Rkb
4GwWfjry8Kd7h2dYVq/3UgWULsz/4daBZg5vG/Q/BIeZinh0ciMu9fSBhQ4IxrDzfwFz8gJb+sOY
aZUb0Bwxw9aTavgjN+rpMsN0gAJbNlPja08tj81MRn4d9SpxrZ3d6r86PMXW9ij+q5fZiSCv+mUz
riG1uKTSSgf0bHnXK/VYmLrGd6yg+IhwyIdAXvmm8Gv8icx3si6xk/9OPgNHs3rwEiJgFjq6RUJ1
HBSCmoKUcB16R10nRnaTBakUk+AOmihSGQyC/817E2EN+PfOd8eFF36bHgrz0UYMOaJczw7rqqhp
nA2/0lYjgJIkLWtShAh/9IUZcFjk1plvoxtGNDAPJ6NAB3C/5CAW7BrT6cJ4Ds0HSsFPNfAaTHO0
wYLs0qPbOCVSY6dsgJP7dcCYGGQQTBHfYmsfIwA7k1CB2/+RsymmcxsiG6sr4+5z+fjOW35UEFfV
fm1GT6TFDHmsbJL5T81n0ZBfC3vTwaazVfGcNJyatGzf15amirJ8tdfAkbuIspUl3ywFtIqZZtVW
9iB2lY9lBsZdVBiSkOP8XqUt9/72MfXTcW633UurYqNw4IJ6blP94qdPGfPff2NmDvv9vdFdpjKk
F/6HDm0sk0ac23m7zpWve2EfrGkPMCKNOb6Qq/QSBwMEH71DGYp4Ozm8IcnS/pmq8qn+HavLQoGg
aaVm3bAMX2wWgmQKXvU9WxSIDBosFWy+BJKa9WXm14bJF3HyqS9GcXpNc+QyFPi4LbvSEpPe1p0I
z+zgIbLptYqW+3Mc7Avx+vj8xlSP0FyAVEQqn6QfOqhNH7d7dmO7qGHJl+uAyPe0j4RzjOsm6XGa
WLdAfPhaI3eCDXsdXNZ6exKNwQH6ZvcjhL6i2CkkiiufYioZf2DaRlU+Psfc/ZdIXoUNq1XbyX17
MYxc+Jz7xpQ1YTCYKND9UlWYCnO6KpGytEfvNw5Wu9tPvq+qPmcOEaRCvSpLA/ftfwx6ZDHUXe77
DMgEGh0Wz1vcTRsVE/CbzxktDnTds2DXdMKvcun/4S60p4ohYY4fe750kO0XV/YKPCYi4nZsqogc
n/FMzSliqkTRp7WQlgdTibZs00nKSQDOESPLav7XHIUdq6kYXf0T72BOvKkURVXl2aKxfZ6I7iMV
/0Gr058qW3Rup0BHuFok2lrAKNtHDw1MtCWLOywA0U8WTK9SXxdIHvs4QFwxGUOkX0TFgPwNwjzn
yhPPtr8Uxqu2es1NIQpOXxSQhRorrpRuxshi7T8fP8AfFOM0hX+GGfGBnGRWQv3rnVEpzmlRyfZz
dd/H89SlcfdoePSDu8vJXv4VEOgWTm4StQOsgC2aoh7KLQQiXZer+LKyW1ac8xqzh4h0DKvXA5HQ
/p0DAfF5gwGXxBNkK8QfOlY6PyJsvOEYB+gMvgPM2mDhyxuEzJXRqUTKh82tRlOfLR22/7teP5HT
VLchBP8Lo2giFzZTHtsCfrABFMP2dKr0x5GvyeCch/M3BzH5zAJRc67uACIm9FiAR94nEClWwlHi
LYY2qwf30n0iyKvt2mIYkl10M+DY7QfiLiCIHb22BR/UpaMdApv0XI+sjR/mQiVBC7ViwIJC4Cey
1A0+45/jmrLKxCwdfKdrDcO5zY3zugMIakspPYHTRB5Hv4NPwl9chdarYFPyXo4uxPSSdSXsmHjV
WAnK4shCCRB7zBnXnLeFoPank+A5bX/7coiO7ulMHRZvS6gTTNjiGbxbC7TCvQhQIbNU1FqoyCb/
fPXvHpaWxa4vmqvQuu6OSPbX/NBa/5xEV9klKEBTWGd0Hk7xD9ed31WTgQCDonSxUgjg1usld8z0
xd2H1QxiyUMGQd24SeqLthj+q0YdSHHcwT9Um7TQ0iAjPOlWzZrwJsJ2uv7RZyQJ5/9d15H7GxPm
ENdhpPDEk12/Evbe5+UdenKC6qli20cY0Q7g3k1Xp6MUdThCqdlD7LmEkYYidRrGSWcojXT7fYLl
WX5mCtC7DZ8aWVAXEAOY/yp8DRhLoJFPGsuRFk0pMBFhYQQvg5zt/fqozoiRiGfLUsTcZ6XIWIQ3
o/mmzxGwFv9DuV0SRzHp5tf7mkCeAYPNiLKDi5R0cGitaqkBGp1rGNhKFve9fWd47qSq/uuoofyM
iA3Ayn0TKPuKk77i8H4gXzQH2tpaTK4D8e2KXpncktcDOoB0d1OX0CiFxkPFmnXOn3uF+ZO4kV38
Gi3N8T8zRbhgJbWmfT5yihqQHBbpMXath5EEHpuP1nJ5Ll4bmpbPOH/jTV7oA5fe4tJZkDMcRvUr
iHFYaIHHaAwEwcIECqgpGJvrsjnggBpb0289VVjeS7TkazMQV0W0V/+sNV+NkeqJzElgtrsDI6ua
rmAvBRpzYzrsvjfrxi+LYn5cqqJwsWE8bA6G3P+PW6detuylzDhNO+16ZV98CFLvolxcb4PnfTK2
UuRH9skdohv7F3QAoqZGW4h0q34fEXCUDHJuVmgXlIZPr/SB6QohZq96r15KDW3+k29bqufuw9KH
vx4Wwj8OypGidlbjtuGU2J7mX/t2xoEl3rbFp/gi/C9OdH+vawdfmgkgAV8wqwfkarlPpkg9kSZa
IwXF/EQWIK9mXReF0L5aqwS8W6yi0DIZD7Iz5gBRc2nVslk7DhLbYsWB5FyF4iRvlT38uIytTN21
k8CTyxryH+3/5Mnga2J01NAfeKfHk7N1+ChlguOcANwZnPL9aj6wr5lIb4r5e1VxR8eOAhdZjPG/
Lt/jLnY6WCvLb5x3n65l9G4b25ozF3TTbIl97xdHos4H8ndh8lhBwOgAEgiDxpzbPEhs6iCYXPYB
3KqouCa6ejPU3GKobX9qHSQxqMjM2ryJXGv0igHWsr/EapEzIcAO5/wBiQor1gkw0O37Y8G9UBhu
dT+hrDOmRazSWjg35trm36U0CplFot6fHSF9/CUDpyvoBsLKvNqjBqyAeLyEASL5fa6SAfM6xyUZ
kyRP2FPThAqFh2X2F74oGzSW+9z8iNsKeJCG6esbPXyMhbfJu0C+b6FDx9htkqWKQ/dvEFI1q7w2
q0N2c8isJfsfpqSYb7kqRcKID6Q7MDlrxCCwvN8gz/lW85XUEI2g+a8C6j3x7GM+4L7vohRmVQMD
mEIz3drauR66t1pe+H/T0AwFGtpEzJ24f0AxvwsZcJHu9wumSvasVlKz6mZYOVaRwu19epjJRufj
n3B9MKV1R48Flw0wfu7HyXmX5yB52ueLAUZophUPAKWSFw54f4RUPMf8syC+3ldHJxNKCxfSje/0
0nF6Q4jecbW2eHNxSqY9O5kgeNF3Tjnqnn2qPi9dnXzzvb6GTYccpro+xd7NQFxcE0Dy1532O0ZX
8ZbpBV4/yZ3inwNApl0HWHe6y/TsIL5S6jTMwxeHtGb9ZuIjrAPjfoVh6wqjqBBtFl8MiGGC0KYr
t1VfYGPPvi2U6fi3KgMN3xjJrHxQdd8Kv1tJ5DyXiVkNCfgSfgxc8T4HbouHnMl8/kr1G2ZVTvh6
2kqM4kCJ6D3ZHdGXQXQKKv9i3g8hIjHpC9BjoRmbQTSdC3HNpxcLf1Mnmmuh1dBMOMupubKmqqaQ
Pm6vfGh1LJ6i+Lx2ysfBLC74gLAKPYVBdlAMigJENRs+KTV45ncWF0sAhU3Bloc3RCvU+n6jS5CQ
ShKJ2A3oLK1PW17q8PwvoG+yBVJTxL8/sfgoXch0hbp0asIAzBBnaV27x397xczTBLShQmT4EWMO
H3kG+2zk4QdmF8lfYMOISgMiXgmO27HjPgF1TC8itKB3k8aoPrqBqbsRY1nxoztBiKrISfLo5jzS
ZTMp8L0Xzc568S8BOthpzsL22muA/GBJAKa7aj7BBlWeSKObIu7K0GTdmuXhI/gk9pxQtzsZCdHQ
ib4GFxntzrVuHkY9d8byMaT8+wJux1oXxQFVO6ThG54bZKPOwizoICYclSfqpmaqZKJnPOD0N7Q/
G8GxKigIxxi366mYK0N90MxreEBdJP9AEbeW2ZW171d5scbEfOH8PCocbYn7h/LdgJcjerxjl5XG
f/8E/mmjFf5+EPZGu8YufFW0AHp+kbgOUrSt5MeHNaFl2y7sZG09iiztpx4H2QqOP+oqo+rxeQH1
Le9YhmckVboyPpLbx4sHhdKdCLmQWVZipx+3UAI/b8Pvnisc6/WBwHNto/moxRoWB+M8Qnx18tro
Mh3y7elG5SxnbH3RCA2A2ZuktjbGxl8c5T8LQZ0dsPwXq6iDYGGRRRBm9HIY0VqeXy29mNBMyI8l
AvMgtFkpqAbv5z5PsRQPecOLPYhWG7ZbLseJRRHoqqFBT4fKUcnMWaAZSWXiezqd/dCCdgKVtpQ1
728zqOFeTVopPDTk+wqlfCeLw0CBVKO4gkAZ+HKXqwXBphdcpnAjpSCBB6K8kth5rFO/KmXmlLGE
6/drcrdWHUwHcFNOqO9nHRwDeUfkhFHHc8ykRf1B4xq/F9XoM+biXC0ddxBEdratILyyN+sC0evm
N/kkjx0Hb+e4pQHZvmcXBJuwL8omnFNWZU+jLVM6I570vfOT5CEjCByQAkdAturNXBpLdiSJHB1x
AuM2CLOafZXYyUPOheFWY5or89ID595crvWKdtDZcmkxEIrZo0lWWp44SefNu6WfjIxN2OeZEE7y
OqtZmsZr28zx91I5Oe+t09iJnmf1VxCbKwLiXg+ANZ5YEHu3pQssAkMpqvtTyer/m6S4OYNXYZh0
hzhZc9lNtKTjZpDyF8n2GhpRSZ1o/9h5WRMftTpeOi0ChS2tFNFegt8c5pJ6uOSrn0fyLGoCFnWC
Xq2JXrS0YKXA3Z6HkZTqSVy9NM5BZ50qoIxJVEDMcCoaXzs9ep2H7bAqy+OwY0q8dGY/zFfxdRgu
8VsI4wdv0SImvXxh1D9XjBQSkInTklqJjd7WGgWuDHgmUcFikpZnXI5QisRDzpoc1wDVYi1/kxAd
DZAXgJysiaR8WZpVI/pse7TYhi++Cuq61f0ri2T8fD6gPVhskBHHmNXMHaCRCJuRVPHMfaiCrl94
FEcUkHr/uqL92tpYZI6nywTmlc+gbHewatU1nmX0wBa9AqPngXwtmBF/T2ODt62XDJHdIfTaiSEa
Eo18HuEeeRkNKF8XJpSS+wupCtNXDwnbyoPeMJVQ2dgQKo4DyYbY9Gui510P3HsjKr1g08twzIvz
08vuWCgGVOC/zCSG3DjkXCQ/pqoZX2q4ryhuILhrG7feJvXVWt4C/sVRxqdRxg78OoWWa4tkTnf5
18WoOnj9tNh68l1enIVdX9UN2O8vHepSe3YPZ95xVW4NziyqNrzFcIsnY7wJj/xJQQNY+cF7t/Ct
7WjLEQzmCCXoV+WEzBsWl6ikMRYkgcO4GV6F9R+FGjtGopZ3C0Jc9jPZlwIRi6jbVuRQ7DE8vzdm
WuDhr9rTc7XuisBtvxB+8f7gaef1iWgPpeP/IFTxVL2rachEGipk8F2zKYn4gNEcjCCu7G1MtwUh
EMDfO9p5AxOCKeYxNrbedRQHx8Y7qFlH3lyKjmyxj9UwDHSSu+wk675di8hkxN+FP3oaBSKLfwMX
VoxpUC19/CNuU6Br5TaUWMuiKnGrBRo3rJIsRz/0sbpWwK/wjee2bY4cXNrCCAAK8dmcPHNfM/Vu
6iaA6/Ddg7LGIrcrbDv/wtL9zCNmaxuEOKpcFTENDZ9trFTv9g3wmK+tJXbnDIUFN3I37eU7+2IZ
lueV6uGjWUbxEgvyIhW6UlpcDxzYivdZCjMw4Z2VwVDJ7HamMPnPvfS3u5opFZrrQXJ2LeZKQiQ4
NvGVW28NBp1REiYji6xZftYWWTNUObFeixVx2mPLtULndGXvBNn3bxn1wUylutxnLNWkL9hp75pq
expzuMZzuQlnmilKKsqkbzC924vbmxL8NGO1GYhi1ttvKYtGy4yxgGGqWCiD25Q6FtGmckyGzPBA
ePnClpGFgATxYdrjXVeVb4XaGbaV6vjO0bA4MQfCRe/72amJtnghJE4ur4qzYNL63jNRMUUk38P6
s5LPJbdSJK0gONaXhmg7UJEZt82mBfR0pFtF0Qozgg1KL05uQPm9Ea9wzNPTcjxAdumMHpd+LCyH
2D2Dmda2tyByOFh0+ZeAXWN+bU+V5pLpWIRqHlinHd9S86eM5CoOAz0CJpbRvFcfk5MzwggTOFUM
0sQO3XVEiayEhy9JfgkSu1tC6u6sZEqCNGixB9Yv5aHIgleQn9tM2kp7SUiUtlAcmOCKWIY1JvIs
d1/nIW28d4TEuW1URIHAufd9InEdZ+dbKZIUlBIWYh4BkNGu8sGlvCYVLt6Ajbn+xn9pBv2Vt3Gj
4LEKi7BAyGFChtS7gC2w/KdmMyvSZFz9/WBxMXZM87GxQQidi8qxtMpW8E4/17In3MJbn6izhoeE
9OX0EGOQxykmRyDnQZ7BdC7/b2XdzSI25j+NApIE2jws7TzLP8ncK31nbpU+gfgA15cdUgnxhdNE
hNqIRMpPPAtmQewnADIE6xmVocJ9GaWyJ9uHmw6dq7UsMZ3dFszZOdnuUHo8FWDfz7QR/bziKbaa
aA3R+edtRJ+i0Qccm0ipWIqjechQ8nbW3G3I2ubCjD/Opla/WRYXswUGdjwNnrRpFXqpPDLUBjde
d2F009L/CNN3EqGZLLNGNLAkTt1Y8aTNE7unPVhPJnu/Gltf19TuIEuK9Ls3YUxX4lr88MpkTsMI
LM3lYezYe34VVEKSx5f4SPs4Um3TCYKt4me3ZNrDdQLHJpTVUczFA9InFRuSpdck6lNtcmNrkMO9
TaZWVFMPWIaLhATRrWv9vPnFjOYoh0FvmVJmAIJPQ1+nAWNPVeQ3qkVxpjVAHSAv39B+g6Urd3fw
hx+kD/mZdy0lOkbhDhFcWDpX3i9eLUleVLKZhQD+qfqgZTzDH2BkXrWqOlajpnDfBFPSBITbqu09
UmcPWow/bv4G+6cVUM8GfgkWpnjDwYlTWG9QregiWL0O07uShYDJSCKxxfY2xiQYyU1LFlTiIaz1
TEe5jicwmX/KdvjPI41/CB/j46lZprVWsJSVsoxIqbJAEWNtGFHdmnlahlqfQobMgQ4T5HSgyBsO
lBAg9AeOnNdzHeTuVO55d+Si/Wfqssx16ICFz8pL4EYMGKcjtDADenybQn2TU55PvNlrxi/LccaU
B1Nz1UfkQP7x+s5FkoGQtOYKG5Uqk/1bQJyzSsK+UIApwKJvFKP/hHpS0MCoMDNp0MnFYFwdFOYd
lKsnsFflD9JFUrnU7oD/GL4t8ROVy/F4RZrerCLTNqMM8LzRgHzz9tqSN3d24a2c3qs6aGz2FapH
RRxOha88jXOH/zzQ4WRRQ4DLCcwlljgqUuqAk7/3FViDQs4WSCfW6g1lkYwklXp89KRicstc4oYr
52KzMAM/utVxSBALP5g7m9sirBUAawR0Gwp+Y0FFljq/qxtMTsniTjPJxpbnzJyK3MJK2FRQghhh
hZmX7Ndpmi37fBs2AvWX/hDVM0pyXxFW5uN8EYfI2xXRlkjR7p89wahVydohOoE172F90WPtXvwE
8AQuvFjQdc9ozSERHM/udbmh3rhPKDB/0xqg097daSBNNckXxDnV817ui/Wihk07J17wuDiuHlOa
Lpr3qy4H4zvJgBjtAnDqEAou6tMwrbxx+fo3MuATrD0eX1LPrIkzoaaAiOFoavTkuWpwSZUP2cq0
uHvERrBYZhAEpQXoOZ4iQknQozjwPoJJoETZ69cYHK7npfPYFsmq7FzMAs3s+UA138gP9mipCm3/
INOPQABrFFkdIpa8Sp3rRh3iVdLqLTEbQmfLZBSVtqN2UDU9zMHHkFZRm57kg8IR/nzjFB5yO9GO
YfS8NV7GNB4DP9PI74UQzE6uFv8HzqPT355rbL8z4BjiCaznvBCDMrVmUy9Qtl++Bkgm8b/iOjTC
kHjA4DCy+e2n0SNcgU3QkrO/9/g+NqisVBD0AUVsXWuKPsYhOZvsQoPrPQqwL4F2pL6EOT9LkBbY
MRyiv8+GH/F0dolMzX425IWcpPFKZ+KXo8aYkYtVVQ36FJMEOXHMoE9d58zwV4klKo7UJSKMDaz9
tHoYyyT9F5UuWXwGvW+fGR0zq7RHrpuHfM2o65il5bS10WPnNX+Wi8qX0uQ26Ut/CdEmLBSi+3Kh
LITmVbrt5vmPNNn8iwWhNXp7xrKS2V3eAKBV+X/QUVhZ5ZDoVBXxlbL7QWQyaTd0goNQJ955mjsI
UiyagQ89FpQEJChv9hPUT1T3dtPWoc3Twylz4ChGvno6K9v/XOkfItWlEtIC0Z68CowLir5VZgrE
ZaOzVY0WLm8iozazrGDY1ob8KZJd5uyIAzHAqz0GVfM6UXWfwldAWUHN8Xjso4ThQ+F6eR/WZi7q
8aNxZJMa+3bgDL47dCXwvUu/tkFvJIUn3VVQx04CsRQhaz/49yP3ki7xiafW4Dpg24xOJOu6r03J
CihEUyBOk2NLGkXukm78SyfV6UqbExhg2eAjuPxBoFbOmrEkKF3FZ5AjaJgumoLmAv3L6gwUaVns
JfgSw1+mahprTHGbvTznpwGuW68igaqbN+hzR2Yko/VfSW3zzmDYcxpCyNfjDCIwc+eeyHwzCE4Y
FGWm9KE+DQ7Oo7HupojKjNVqXdquY8Srb5agw8dnjLXdJUUdOuDBZ9gmepJMYWXi49Idb0kpE5P0
eCwshRQOJonhbjm4X/AgnCkBKwhcE1NrqBNmd9YdJ1TwUAYxjk/9rmBBxYAdB4j3miOKjkGm5nKj
iu979HWhHdaUJBXU1WdVVBOy+gx380AcuUwQ9XXKA0WLDQYKnioY+Zl57SLvkpbCT1TY8k9uvGR6
bGaNvg1O001cuUtaq0Ft+aNMv+9x6b6Pmakeeegf78ZTnYK/qactShMGcc3wOlzLBEqdLiLaAVd7
DoNXLmRaUuX2iFr7jll3a13Ltl3j+xicdcScNw+c6Njehg/3UzKzV+46TCNNn+dIrfouPj1479cn
pGcyGAfZrSNJYlc6B+6PRF8lAb4iLi7Y1sk6P1ju+3WRG5r4LPd+IQ+iUDmYrdYFOdoYeAIDE5yJ
ZYCoOsE3/vDGOt8cyz5leDzy24VtXN40N2IH/l5H0Bqgr0Ng6YcLp0UcLjWVR2xt2B+ageMKHgbv
EkymojUxk2ejQ0s93994dhyc6pCOp0GcULwqgZuKWEUZa09wiAX0RswV9NOCN4yWYdlp7uVAjtQ9
9PJE0oCvhhHEBDqvjs05Rytj5UA2l9gOFV3/4gabegEDQkshuL8H4XZD5V0g8YvQnluy+VA9It3g
ZShhLKyxQayLjZmYOCsEK6G5eke7/W2CquIHRNwcRmqNo2Y9JeKoAy6dSSGthAnkffPtkdnt1Y0y
rO2zsthyoxDixRLpOegSFalspHoWQ/Ux2T9ajHbmKeVl+dmpsBM7I+kgy7YRyZHjJOsC2tEPLyFr
NJnEKc7sejX7xgWy1sZ/jGSlH5ceyZjQkarp9C7HWrwp7KzLiIjH4F+3iOcI9QWDyNdtHvtKJY/J
SdBgUPbB5O/VVRz/ITPR4AjcPk7BZW800wpVAOwdTRVnJOINeo6lRHHv85ovstErSIVi0G8HE8UC
hziJlJY+tOCGnVd+K6vqzQNRUx2muaR3ZiMo1xxNU7ZnuXU4JVk2MbcJhvOOBGdmwTQWSVabIGGq
9TxfrEz6P8XsXoW25BKNJh+8zT07YeMlm/FXfQtioB9IjEa7V1bvvJ6ZoyoODlYT3NrqZODUqGIc
T1xsZNc+6PXDtxV9O/agm0viFdBHpcpCaF7YlcuD+KFQWQgOAR+RMnfM+Ad+OzkgiR+JTJZGzWbL
Fn03ZmnNLXzAZfIyiTX1Pb+5gH8ZS8ezo9bDqjftROJuOxCmqHFxsGt8rWTgVVNesoakAjkqouLP
SvZOco9QTsTfBDMyciheUL9D2M0OHvcDGMjy7f/2ve6i4CN55hPwMov5gwcAdivZCRHMbDG/x6wD
a5Lz+NQR5tpt0TF8N+DHLQu6bxkDezNtczBZ7MIkj6FtYkWg7C362s4iJYp1m3Kql3Om+vO44Yca
99IpvqQPTYF1hGOaWj/BIQMl2EQjuSBjOibhlZhxheecCyE/til+odQ1M6HbzayUDiNuAXathvfX
YSN1SCJrtW1vgYYVtZY1dTEZrK+jD3DNmbDrnP02YEzHKVbuLahKfkfZk+Qky3uErOSCJNaObNjX
vfzDz89xj9IFeapR3o8+M98VXFeZtaQuY0+8HyCDQM3tpO7ECj2HskFQGodF543jYmaLZScDXuAD
a//FUF8OXtiNlj2LWdiJzWTUvUeJPGWPHNkQ/vpLiZuNWxJFdRN6OYSZkm8tRG4/SDp8T3FZkYTm
m8Nqlws6x113Uj1ApePd73gIhtHFxxWef54xeWUSih+0DAxIL8nxEKqG1IQPS+rOK6Tsyv/LVj+8
MMRm//r/y04IBiBc9UMFH+U4Gy+8i43BfL98O7UI8Uxy+6K8BGbUIk7bCWTINgLGrWeISARHtDma
kL8k5PWNo7mbi5vix8V4bEhe6HkBjKjsMJ5nsByUxMSjLKHIKkVjBTDFWGSQscdJbcVKJQNVyAR5
G0RbsCvMpjb5EI6OQIJy+bLfdBIpu1FQaBmdXnm79mdIOpD9+8yIywHCkexZyvGxifuleQHcUNQn
HKwfnGQJ1Wbh7ggFQbN5BnHZpnIl17EGEgLxpV7kLUIOnUS0g/nNOtqr68eNz23lqFW46n6g/+D8
W5BAYb+laZfQFUWtIe5Btuc44CvrHLAHyv8GtesIzg7JKS+MYyyLOd5yr/C5x1eZXgmpis/xAM5c
y5p5artlb/9Hs8Fs2sSQtXupGvfgg+VuoxGBhvO/S7/VpQZhjXO0hr0KWAsNSY71mOZzG+gq3bbX
69Z3vZZY8HSswA02rJYc5563K+jfVV2/fKgXRZAaKyT3a7We867hbJu3HFyaHD9vr+iTTu4NidHJ
46DEYS1oluQ2zg7Xx5g50HQbNDHBiU4O+G2epg7XOn968QkkOBLVLs3sEIeNX/Iao9gwslEArM67
r5DEB+SGJxVZ1sdkMyctJCaEBFbYiXzi/Q9+EbHz0Bo0GXI2VQ4PUgDdWszbIZZT5efwim3CXfgZ
3BmnJztZzzyl7ZyuA2s6ctVeyCmNEXIKjAJFKPweL1guLXJLU4nz5+2RazkiK3O9RFFpBHPVsC9L
f7WCGXFzjUSk/J5hTX/7W5Gg7JGg8QgnOn/kIh/2CSIWrg4vAxKp81BTSwORVn5mt1f8X0KG0KH0
5KtFwAKpFKtnzlJzsVMO8Z+3eJyoDafDymnPCZlrxnASANVwfce75V46ZXOAK+3PCiRNZu9xup4M
GS5IZPMBV7sVGg64quVzXzIMArzLjdMZadwZBGBHBB/1PTDrtYElnN00XrnUVZfXvabnYwAVEEIa
N47Q8lDIwaUFqE3cK/LDYFp23YvsOFxVO+ZsDZBTDobXcJqQETVZEkRmB2KxGl5LV7wl4U6k+53W
Afa88cBk5KFxOJUubdTiLDQOWdULUz7fMR00J+4+FwFaP6Nq7eMyKy9hW1OzGgvXC2pNIMuYMGz5
SCttchS/rTLK9BDiKB/SI4/Gvs357qOv3a6z852E1sRj6jXe/olITO1tZUOzVoa+LLDxkh+DV+IP
nm0FvFvSs2jWtziquNui2jPCLAwUiRmFGEZWI4l1DW6EkIsbPijiLMaJw/YdKIaF0OwzmvOri6DH
o5LUZzCoP0l6UW3O0mIwKCbc4uKk/1UrT4YkwL/SiVuhyi5/epjlcbZHI67PxyrY5omMKp15/RwE
f+250bFzHQojMPfFQo1KW9zIUU21+Kt5tTo6xgTHYhrsc6tBgPn4RaDO/tESUsr09/XcDQPxt3fY
EMq3fiOnjMhTpvpT9c2p5gCuAEZ9HN/GjtaiRjNMMHE0CGtnyKajBN8JygWTvZyp9oB8J+GUQw9H
rBLqSf2PY3apt2wqUx3UvSYPU8/hivUo69j15NtHPnalzyxExu/ObwAeuDNrOV4+uD1B0uRxC4cd
YBm0tYOsJl11vV7uXJWUC43T781dxg2A+iPA02lFhTP01kaMXQFkaPlaFLZ6R8AeTg2RmodBU13o
yOrLDkdDRw3GnEGWT9UaK53ohBbEpM0Nl0CpZtSBU0nIt+WBps/jl64LydR/4f7VRwkQ6StAKuSl
qAISTMTOARs4/kVxhsZdbMMVDQlGH2rMVNSuFMIGs7yqstVTa1HyDEHzroZJajepTvkboiH/EupW
aI3bVjgGkYr5pIIeZRqKetGzHg5pzYECdKmdIwGc9HLeO3UyXJVXB4mM32CdKs2xZUbiQVnDkLm1
jYAWNaVtgk+jpJQ9kQKMrZK2BIHKXKk3OIVk2rL28+/9hcJ4clkFvXn9xw4Kgn79GpMa2EzwKdhZ
tHzfOzLAOHIVx/k9wKi1rrjJl9FHygPH6E/VvfZ0ZEn/yj8rBlAUzN4xkNPL9FrmniPP7UePwXsu
UWOzpAwNL4bzQqgeLjVLo+sjrcIEOn87UbDWjeRwxLshFTvCEr46IVoC11IVBmrY0XnZY+qCQFfM
rX0XNu1JZeHj3gZKEDruLhatjVxLHBrhduZu8vyKeXxScZkvukoqI3ijLQ4/vfCEP84hZNnBWXOn
n+Fm4UOJiNfM6v4llaKuXyD/IrzWmLj4HjjTABSeT7a2VH/bRuPMJwLpAlfgH2aYjeeAPMwicARX
VDNYUYd93iVyCKF9H5NyO6W8L0KtliAT5Ad0FpYqgP7q0ytypPUKeL0wSYegAGPzcoISOV/l1rfo
2HFK5x0sEbOsEs1cDf/iGHIS6/HnHrIuh0TiVpcAO6SlyJY4cOBkeaSRpWiWB1uGPujgXVmyZzNT
QWN0bns8DSThF6p1KdYo/ObAjQebzx9Ii44zhAIwBvF9tLYC4gqYa0poa31w980o2EkiWuON4XeU
U/U83V1vjUj9/+0gPUFi0FsYSC65HjsQvLnE8YAc/gPs7ZiXkCctbqWu949YlFtXGdmPFIY5xlwa
zgoai14Qa/+glNQ8Dqy1BTtCZYXFkTEGaYP1d+pdEU/Ph2hi/GurgnTZboVNJ1ETEF4x6vFJE7zb
sc1sQ5FQEQ3+2Z/8AojJhyQtLnFoc3re18CXT4A09syQ6FSJeOIZVEezgdhLWd/NwZqxdyOfzaRV
ZTy6FtR6v+uuzPNBmvSaTKnGnbrdLq+AXgR3qDN6AHyVMMC57FtWLfIirQgI13PQ7A4pssulJQM/
yQCJbhw/VlBLJUwMaErTMvmCBDz309X9iKRJhx0GG8rLPTMCANu1c31bf8ay3Oh1yzCv4YjVmQLW
W+9zojZgT/X2V4y+f3rdtXueI+ADrZBKFCa/vYmu0H781oAcGSUwuTyKeW9mnOn5KVjl37mJeTEa
SfDQXP1LRDkk5ILtTP/hMtoSt7ItHvbrEBUg1k5UnXJmNBWUJu9R6GcnZnZcenwi9xUXGeV22Lgv
YOyDQzp4YMWGdI6U/Xmn4O102Bj+O7QrgXRNbAhwOsNikjbuSnLAndE9HH/6bs8c5QDco0vnjHo2
2FQBIZGhDkGpEgcaZZnsqGEcQesAm2f8P3HHVdMiXZGkU64GCJvUPJ6x1ij35oqb2SzJEjmn3Nup
Xke6LWeolp4NUDCOnBW8DvvewzhFeCDZJhA/L8+S3zVr7FPvzhnSWmYyiOePjd+8jUUjpFC0AgTv
sQp5tmaY5w0YSIo26op1Q+aN8v51jRaG2fA+WWTbB8GAo8ryVJ1bIKnDrCEdD4BvFN9actgUHa6o
yl5XY08lJSUS6rzLHdDxh97w/XNfdpKJ2+yZjfxqPS8oTlPXLp2D5nEkBEg5x/MXg4nhNz7S/aCI
GAfvDAOSkBCzEiVR+GJxFID1iOs9eaAbwRoxZxQK27DogCYl7WmMLN2SRJwKfQ22O1qHjBJP0mh8
fZLiOXzysnzXRAFYVdwDxDAqCI54wkvYXsgttZephQsskL37uL8n9z94VVYiyov+3DfhI5sUBpbl
nNBffKKsM4OYD+bHHy36/L3Eg+akhQUJXZmNfUJaN9/zSws/qRHW83/gxaGe5+AJ0SBngdW78TgV
NyEk6nQmbFCJp27h3/hMenfHNHDHjJ9AinzHy+nSvZ5qQeaVf6Wqf3O+zZgI3ucwAwtozlYDR21i
6zywpKPAYaH4jGDxViEAYZNwTdC8YjA6+21Sda9Q5TngFXJfSXmuuAwOqKVKNWUhJ8N1CM47Y3xh
YWKQIhWALSnJPjqcsQh0Aq36txwX4QTtNmBGFHPJOB9b/fFLVegKtnYvn32WBJ+oTDEqPbHBRlvT
tRWQR3CrLrMh4szXJuxM3eE7a5Pu0T5a45+P+SofOPsCYgtKo7bJq/j6H59JjNyNLbzeiawdQx4W
P7Sao3IqkIsI1lSQqTO4xvVPT3tspvDgUH1X72Anu+AKeGw2TTHaqplvNXVbkr1+wwU4GauvKaq3
AFSSrX3FDNVaTvXECSnTG3evlVf+kxq/EHOUmKSD0vqe1SLs3kkImNEIagcQKrmbcBsB++fVeygj
UqyljFldpcUjOtkhpyP41pHcTDU1K6N8qHJvFqycTRl5SWJgQkUsHEdUzO+p/WQfDwlDeKcWKHS6
L8SyRn3E8TS1ALzadvoyHRlRSM/ZTMkOBCVtZrUR748aZC4HEbP5CXs3LhfMqqc+w1WqLfnfzbTF
dEEvyJW/1ywyx/nuPbi3G2W82s7o2GXDsof1I3nve8Mgm4iYJ0ywPl+cjoi+a+AuDSHD7ZejTdg2
1xXa8vP/mi6ssEma6SanO0H8rEQwMuKJGO94YO5MgHs+lBCXe5CPFG7IaE4ZhT0nQDiUzzx6ZujB
vyN4Rbjsav8EBq3hyvPIWNTY2A8ULEvtOmZOa0MCK2VlsMk3tmn6dBhrYCjzsGzd3B6iK5xwHwp2
cSnyika81zUXpa0yYa8RkL29U5+SJ/2ln4RrIT1O0tVn0fcUt1rWOjkWKeU90dhj72pZEec1Q4md
2PE0rakLOCN52TKCs7NdVrPAMZFZLL3hHTOy71wv5Avja2rhSsYZS+h9CLCwp4i62clrNtj/Hju+
/dsCKBPNs1gFw5H/kCBs7ooqE3OjAHDPzdgLiyX9NlDDlyF8XkOOMn5Dbe4q5x9GsfyiTcF9JM97
fCxdV8LMMTFuevGBu6lVmy6nRHd+tY5aDZp1Jl2uLKq1Y2/R6noiw77COObHFQ+A5UyIkKByFdLc
hmEl1VkE5W4a90eWNZslgIkcpUbj/1ByJNwokGUA3E5Xk5ycN87NZwRmRcJi/Q9R0oBFRJ0ykg9P
OV6sGBcofiYW6Ta5evocrJITSZJB/pzJqmM/h+dlJjSaAAO1pJiIAzDxULMHqSdQ03pd2rTnX9b4
hhfqMfm8WmrvZIVraRbfLKX5WdTVmr85V6LhpbZFfv4kXpFVm3TQpfhIKqRFWeSSar+qAR+YGIWe
eDC5QVkL0vgncwMxguXyZHu+h8A2ckVNy7ji4z5cVRI/04KtaRTTdA3sR1Cynk+ZjdDOKna0NfiT
dt5sdLRmbVMhmnrxotzmF+N5+S10Vjd8hojvSOv7lgXXa1zIh7L99Hr8cKQmVJf+/r0Gir7Ip5or
Cvq1jrnGjxKTegmdVDM4V+de+W070wbhQ8Gh+GK8QF1hOYznKFHpZhDN0xTz4YsW0C9i2coo79ZR
6NDODoD/KNvRaSTX0sZA9SLuynxEETG0RfQNoAlHZCcN0B9MeQK1WagqSlgp8/nChuWZx0KiCCHH
5g2AKawoVOUFQVbOMM7Bssbqk6zPXYmCrZmC3PEYLl/+C6d6tZe+AWbDMMo6xVd+ERdECdCNQypl
EpcC9N2PQ7IBgYLkm8e/Y5bjWPvjgSOPeg5mi1kqPjfqMgIdP7V0bmNhjWZh52Lx08MAqd+6wI6G
yk6DxgadrByhEtgbhUByhvOeolUQhwfmchcHeo0oRYpbYgZ9iRfXHlI48bS+emwO8OZl92cLm3rG
BsNMLX86fUELAAqcDT3+8ljJOTyzii9VwXpyv06CY6xUO3c0c3SOhi03R08QyTteiq/ygOpYW7+Z
kEIs7Ii8Xqcx9CwkGf3ZSL+hLcu4oQoa0lPK1JeUvVlkYX3eOhytjX7rtBO8cK5Do+ICMwmbx7jj
yrJLxUuoABe23hiwW9KETDC2zb78Z/doEf2+vxI0c4hvpuEecOTxjFIHYx2uBS7ZqeCH2Qk7IGeU
Kws7UBwbUjx1762q4kR02OwSuXZGaIHqGtzVl+C+zm6DCkYlM26oGxx3QCgNsy/7aoJeH6w9r0Ox
A92GhdnCrOgZKInoqDAJFOUoejw3v1HcI+jJRZCQl+HdzoOKsbEqg7J8UwG5qscWa1O6+Qt0gWnf
fl4LS14IjlnoKaR0KGQtopDhD0z0j5swVNiD8ehyBwnHMr2fQw0KYhd6ezDepbplwN1A2gxFOe3t
SvbfAtF/cvsjP4UC2TKwWJtgP5pmwHYhWCD/LBJ5ajcCtinwNrf9Iq5aWuCkZkVruBu0PZrWT+nV
5hQX4D7J8QngELAHuAZVjBQRgylKaHCJa2Xc7sb4ra4wli3FBbZ1wMuItwANlz8NDp6GTQxXeEya
rmOu53krba6MmNDaCKnNMYusirbzZjUsw6EyswGBsJEUt/ibtj6ORmObDI+lj0WrXbJeANrLGhRw
ob6IinLw3DO81gJJaPUrA0u6WISs6a8ys3rx0LHkT9Rwh0vKfEVf8c2uJvTAOrCD7PKW8nHuCY0f
dPQLxJHAi/IujIR3XeGbtCLSF/eLOMkKUz2OmsSWfVJmuQNynS6LdGMq2Cp7cJIu3vvjO6bx8w73
mZCK8nE+UoSj1Jk4qQUKUHVRIndl8hokwQOHueDFfo+vE7ed67JQdpqhF5u5xGj/rRd/qu2m5kDc
PhLKjbi65hxvFBheo7drszpLedAZnBNUMK4+5pp3MQGgNLvdjrxDud/V72khB/6w+WPpIo1ckUM4
FaiNnsmZ2mLjMzH2YW5O4TFPsEWWSWrnyVxkjlnr2e3yY9YVdwYwNYp9vQwMK+O3gEY14d4QLroC
5saeMuw2q9ii6vF2/z3gyZJLPP9d15x9Uktp+3T+Ch+Gc0ZoBU4r/HaR/M6B+CB4HJ2EJsUe0TQM
JefLocvXaWSBNzyaL034KRacsMOcOFPr7sRVYFv3lv8afxGA6Urv1/2+JvdHF5FBpTxHwz33xQIN
GO1L2DOLQC6ze/v7qhp8+smdvb2gWR0EHFxs7Ukv7jQ2U6P4yPtAo7WnRZugVX9aJuW0NcUCb3Tp
YRLyAZN/V4orNXOOc9YgVZw8Wpv226aLtakFe5DAMehYuqnnCgkOurKMVF7hzT4sqkKafqAdYN/q
SXw2jEIFWcdNW48gsBLPteThCDDXimQgyOUQDtmSTPNAwTwQzhRWdMjsZAtr8TC4ixriCnpS/M3r
t3MrkkjG/iKZHfzcCT+Kz1Uyb4VS69EzTAVTvJqserzAet6e/glxfxw1yowjJQmF+9inOiXeZFlF
haROABWhflyhlY6iFiY+mkkh6FjyL/pvtz7gymvdspmlQ82twZsWsvT9ol4reYlJym8hW+Th2MJS
nNzVNHd7s9Hoy5sg6EnLgp0H7rCk/x9+8Iqx7g2RxFz8aLOJkXFynWMKudqCOtJlKZ6nh9WUu1BS
swyShAM8lwmpfZT0Ura2DWtAs+xER8TVFpJKGn2jpq1OewO6xYtIzUKvbBmG1hmRDWrVPd0j8hbg
uh4E+InJrqVzyf1lqM1ftzwour7710ZgzjmP6kiVA7JwEBu7eXalNO0DZ2LEiYheCMOWDLeaPNPl
0N9byxwepVac5tWIIBoVsdf4rlVkQRhAPVEikhYPzhIZeEg0aVIqu4ALX1rQwoCtf6HJHqqjroJ7
ATH0RINSrvl+9rmwwiR2VCUpChP6hu8X3GAJKtL+RUBj921Q76eRR8+xgwb6UUTFwBTS8BUZwnH0
wJEWVmNu7/+t76FRhEErPkgeZl9cjLMYZYmzPTzdq/2UrHuAephVPyN+iN1XemyBT6XwZfbVNqV6
3S4hON2YDyjniJA02EhFdKNsbKo8FXn0eB9Ez4lV1aiU7owXKHlCqFupD4i8iyXyJzIV1lFjX9N/
L+4eCPbZyIHQELR77pwS8kY3rM4fCdQp7Faqwe25OqjiS+/CmNovFKT7BDDsQ5QAyzLzf/AQnNNH
RvdiLT1o/p3kj47qPVbynwj20kz04A0JgvQKsr7B/z1ROXcB50RldQ8zi7VsZ0h0KpABsAVy4GmE
S8MeJ9xztniRKSkzKtvHsN4AB5yJ7Zwcq8pzUfQZbsz1W9LSA08WaDPkNWYGiBc3ZiQPlho447ZW
zlnS5FZfVOYjtwPHALISr6sWQbQnPCT8UYmZ8G1HfiACFNPpsKDnhKY2k9CwmJj8JFCZAeV00uZ0
8gL4vZj53J0WA76xIidyEqv/4tHiS9bnLpww7UVjM9eTj/rwFFoMX+x9lK0XiAsJdw1xYZwXjJ4f
s7+nbCuFh61edvlUZeWHSeSKtTccFt8Pq9HQrcAxJFKgVXQR9oL4YSxD86kfzw8OBAsQicZW33/7
bRVlP+bwYaQTf8ONvL1CmIwEuomU7l1m02O1REaEpH3v/7GJsHFbRQSPdi62LbyWjiYRlaA9w5+x
CsBgMtADlzVCVNHxWmJ1alwn74GgCdr8d7YQ+WElffPz5NvJX6spqv6oqAXiwE6yERJ0IOmA0bwS
8BwaQbBfIC7/6+khEGQ3eO5eq7BbMfE7tLb2tSHPIcWMs3/OMAHqnPXGMrGkZPyaPmO2yTluieql
YU/HK9fVR6yEvw7IJIL1dET2N4YKgf7Lnr/N7Y1xEyNZJ7i2Fx1JPzbPZjt2P1MGZ1s9FddVT4Qi
2kv6fnqFQKNgd0y8+ZXuUc0TS05A1ELJjuBBXk7xPRiNLpdF7kt2sPwIasa3ETPCnHondZnbBkeF
zhlk0MmohsRix/AJyZeis3f7xiy7x32x0DynIsEJCH3oxOa02JIHlf3wI+uXNiX2s7atzaPT/6xP
+4hRQSM1JGk2RBlvaOX5NXpC1NpS2PeeSvCCNvIgIDcirngcmXejA1EL0mnPgQHwF5GWP93IpHYj
Fimxc5FoYPEXDSmclyC/sX40Xp7iTnTkaal9+7Vl9c+9DmOE0541e3RxFOX+WZcOPPj4WPGZiGWH
0t8knbcsLGr2wbfXR3NYs/OZLlW3MUDvWTHYi+9tbg8oBzdjfusom2X+1Ndl3+PDuRPsiWW2+QbL
r1lAI/VMevqPjlBxac1gSMY/SWov5SjUWloFA2cvE6zHV1guRw+vJjpl9iXlOD2wy28/2kufayoX
fMtrtgDIClwFZJDOYvWdR8bdXraeH9nVVpaIEQZJYxHmXp8N+L81LkQJg/FzOIfohUPHrwKm4tsz
M3ESJJtyPhJeBaEbU4czhqzDkLmGtCNixxG83yfF5qFl2hif1U90JwbKD1jq6WdbT13Rv4hekByR
6F7ydijRpuqFeWBHU7R5fF0yGcACtW18BkYIPGwRCBZpMfzkdAXucl9ljp4KOGsG4LshC8kKXMxI
5EtLjYDiUARDqFn6Dhjld2JY1R6+J1MGYPzo/EXe7naSuMiIWh7x9SWTcWCVsXBb3Dtk24fuSJIO
KiUoCET4D9yBgC/ec8xkZGasNXqwPxEbJMJUJP9Du8uW2VqR/AVkdbebpM6i9YNsEfUqI5eBX3N/
4MPglaDCIStAlliyqaCz5k4UOh4VRU+bhEU3AhcKHm8YjdbWodoOX7wz2moq9IkKN7x4YzDTzrkZ
zpKR1zDi9Lyv2B9w2Iwxvi8REBUbcy2lOPJHR3dTeajuK4JfhW65A4Nz9JVKzceLlYx+1G7JHK2E
vJCmNQ9wvf1/XMQpzLBUu+Xzf2OrO3NlavRVecssYB5Sr7OY3gsIhGZbVfU0sDFqqVu/GoKeCcSB
pVTKxda/Gqw+JrK+RVGqG6+KiR/IYPSDEm3K0naoWIduJPcjgFoClfDEnfkjmxrcU5YM7FVvRJyy
bnjDt284WALGdkNgMaYf21o0ZX7ImGaOggQLbrpAHq4WAuH/Dyr9ahU/9L0S3J3Io5MwYYPjM8dZ
bXNqOmVSVuzRsam84etZRrWgq5/C+zM9EO0Q57dDDXj2PiHn528uihcXJ58pn5flssk3BDXJXQg8
tQc3oha/hJWcZL3o4R1d/DH8ZTW9bWb8CE2gj2Q1Bhnj+O/cVGaHjkdGbp/cSe0NiFeJIikbVgo3
y0Hjum4IXESwcn40lFPh0EpKsk1vqTPjCAEood4TfSg9BIiIeSLLXPoUaLJVluxWQkFCA/gRRgzP
FafPXndlcfdBzNxKSTBCodyslAGPdNNOGslvFUkG9AxPjePFceaHmdqzrB1PmHwxHoV7Yy+94bR0
Q/Trze5FjQk3GGtSw3NNCz6FpSSnO4v2nh9iIqtIs6zkRkaci18sOZcxxxmlfKQe0k9zROdueQny
UO782cmFeDGIXQ1UbjIa3At8JtBF2ptheqKRcTKjdM9eFaw+/oAYZJsHdSWusjHT73C5EHkaeS1P
nY0DD+sSqjsr2jfhoOWTECX3VC7U6EkZ8Qjamb+CgX/DjuRmAMcWk5wDa7oGwuH94v0dNgjjkb/D
PGMDMY8DnMA1lSbEEf/U9uXPa/IDh7jGKw7qClfrk/uyzkVb8Ao78TebwpPeO8/Fv//q6ldWMe0I
5BTGv5+qT8yXBmJo8Tbeh3twng7Ryqfzwvx2x9yc5jniw9PksTyogOoc8u2fqhSD2g9w4qFWPuPI
5014Lrdt+VzpkXdpptE3HivYi7aHVYYIfF2ixX+cCBlNF1l3P7eqWTedMjMPQDMFPMhjQaXCZSGu
vfJQkQaOEophiPFMbkE/Aw1egXfBkB3/jYBXp6FQZtTNt4kTFCzsLj75u/Q8jNfEtxRjO9tLAhDF
mArHwlHbxsEL8TBgCmR7c1+3gL/IPJkmnY/0U9bUDKrRBQLuQuHVa0Tdow5bnqoliY2bZpya8dok
Q4FK09L6TO8VUf5pdTsTkUtgqOHSzBggzLTTJdUOgS3Oi3Kh3HlWXFXlv69OJ7mXGGgJHvMjO9JY
9cHQr3n+468+FdDA6PsEBmePAiyc4PPbTxhLNrIRUuNah5NPFWO1ODkDX0bk86HOg5aFUZpwVTut
8zvYT/u43x5Tpyc7oXqrsm3uEZUhB/s9O5VXdWekBTbG6TUQoKfN+2OBGpXK1um1vPgHpqaQdmDg
DD7OAd1R8I/chW2czBJjfsztJiJj6Ogo11kAhKUSlttEloyo9/E4QW8UjNl2ny7TsC4+Yac+i9+b
uS5gKnZCIHM431bGgZcu0CjUGqTbd/0DPQcaNmNopOl/eb2oRt20jOhJO8dBcxCqt4skY9LPhvDq
hRiVoJqskIiX1MUbTetIHgOF2VaCYoDeGqWziQuMoiqKovmTAtzfGtkx+2KN9ajrwvS4YKhWu+JO
5fLUmBzL1OSM+hgDB6IyOKU71VPuP3cMeKhiRpW6hA70CGPV/lnv8f7nQQD0Zj9oEt/hFZAtidg0
SYdnGaHLFkX0LpCxf6VyAKMRaDwmWZiFEybU1LIkoVDIwLi+5FBS4PsAzrDdca/rFrvJH5UTzanI
T3+97KTO3IGNEqZZvL76oQmNBeQcJ1l/4NOm650Z+XRZUZrFyc1w/Mfb9ZARCSg7UNPB/f9HZpD3
R/H+UH1q3AoH05+B9mTSMMbey4YAyEhe1ElIvzwZJxjS22tIoPnSrw+h/BijOr0Ftilv0XJtBzoC
xxNE9heT6xRtwXyDkdrqs8N5Jywgl0WRGBzfYuquBSmS7cwFoY7pxxf/fmp2t6I71p8wEZ1PFhNY
JJlYahJKe2eU+Fvf+0BMMxtboAPitIW8KChd8yuzC9dHEGGOETGbKW5hfkN6B8Czkm7NinvAZ4hr
HRy1u6pTxulDSqtCDVvJqsxfV0d9TKO0QDRptUf1CB28kfy7rtT7GWMF2FX/J3BvsMA17zOArUXZ
eDsgY3/IK0w65BFfqu/G38Z4QIOaK6hiTuekH88G3E5EMtdfEBRBWZjymMmxEQoYA7T9Ep9+qsLT
3kg/KC9vx0B7DDtbGF+Oih9u8ZhQXKyeWjSgokZH/qT3c5Th9aqe6eDlbXh/3p/uodVwGSEA0Ymv
qeUyFUsSYVEifnV+zN0YFQRAkqY6+xTKyL5UMiC+gew1r6x7NgPX20TxtHYfnTIeXtc/E1zxBlDE
Q5vBoCr2uvyVAZqiq1hGg7hPxegUICi4Wr+1JX6U/YKjwEotbZg1LVPdY/6BIYJIiSZ7qtqQUqxU
AX4vgCWpQy/Ocy4icyZZfBnu466yjLqnsE06cN0xgw/jfbp0VbrGd1eUi8YnPOcsMsLzxmBdSD8t
R0vWXOafPQhaFLkemuCRxLkTdkMrTHY0pDO65S46mHSzE2MVdlu6uRniLpqMjhm3YvJHI7KKFbLG
qMsA+ygk1qwnOtkJVnhFCvjjby0zjlPA/+gt1EWzplQJmqebroDTyPxjnWQIXfn4YFvzalRTPL8e
zT2hs3k/l5n4Wv06PVNzh9/0+5UwXI4cGiaKE88xcR0esQZxgJ9USMtK7SU5lh+9a+k5ZWA+9Ez/
YXjPUPTuBos2SvKKlR4hvm8qa15Y/R3s76UYcMVHLFEMS4srQjPVnTjLmfQsgRW00S7odObwOr2Y
xCTxStqFXvCwzrXl9WUuvsCvL8R5nFX4iIWe54UXXrvenPQymkVQu5SCPh+mCRjv0ntKZrGUOfxL
TgZwZiP4H1uNa5TrrOkp66g2LsB4rvDjrj3qMMpaOVa+jSbkBurVpyZ6uuugvBABIaXgyU+S1wvH
02CTPN9ZNrsGqlR0Fr2JuSmuVhOnSJuIpCbka7SitnI1eXdWMgnOp+/RfsV7/4yo6IL/VVx9KfYo
BAXAdNse/2jRWXiAGCvdcW5f9K3Kzxg+T7P3lfA0x0IdIXvY6lWjjQMHTKDOCn/uVYzhBgC0XSF+
PQd9EHDoKl9lDopX0WzDBUbokLuzfXm29MesKUvsdv/XTQSVWD0+ZDaFniTAgSeB69N0ZBxiJCAp
teOh1UF+vf/duHkrYDpV6m1RDCFkqNI9PPJqFlm91yv+V7WejkLjaA5cRuak+za9W3tmXdXVCEGK
1RSfQJMP2x/d1fQmIV016UYZ4s5uSTKAcSpixiMrkRBAJeZwaVqHFCzpXossx3gX7Pl0a9G4rqts
bSExrqwR997UYEfXYaUINi/YrqLOz82tGibar3j2BSPLrcisYyHWLRSDrgr7SPtMPNr5NH1whf2Z
kZfvSWUniB4DTBE5Sa9MGUSx4bgZJUJAUm6rDImI5Q+yzuP2mNJSEcIYZLQkA77gUjqadp4ZqtzH
k1cSSGJkKFFg33BwpcztSiMIT5uq/e7buzxNPGrueMhPZPZQ2s9RFOygZFY0u4OTXbVOfnWNFz1D
sKuVAM0zz1cYGGFW0x7TYApB2eIEgpEOTFDJnr15LKgjJBY54YlT/JwvdeLuxCAvtG8tw1xTC4nJ
raRktoYJ4QJNA4/Sp8YsVd3ip2smMSUdnktuX//8t+yflyHEoo2d5sOZSEhlhPX4Szhpes9jhU1R
BkGXOuvD8YOjsf+073VTrvTVpBgFkkIAl9S2VBgGyoqtbf5wCpHeU4rFC+NyEIr3isuIz8faYDe8
v8krk9HNZHYsEsNDxOkzvtIHcRZoB5KiUIx53YAw9wsHLpY48kDqslLD6HMJD2IR2/2VuEilDHLZ
QuvAPYVIICt0ruaTYYkcZjpHPv4UmWjMkS0u9GEVo8gAaKEqS9iwNijrElI8qjwjmpiZgejXFViI
lsxFLCvH8xnSMySKgwVL2eFgLMF1WSwdfkPkc8V7GcB1JZlJXDv52QpRjQEw5Lv8oPvTRO5mgLTN
Oy0XUMi3BVCmVeT6ufafIZCTdgR/9PgsDABWyYVMh5fyAySOrFOFJkbJaMWp6mFyZdfWJBcbH8/O
aBcs6AEnipbfufn+uAiu1LS9ad8d6iPvSlgWL/eHXEnd12Bysx2idFXOlJZTjdbhWdYhA5C3mOj/
YH4FeFaUmcHkuztt32eOFGk1f2+Bdor+DJVyq2RwJFyu1RfXbqbvs9OMJHeBSn96i7AK894ZECWB
xygMY9E36bkE610zRFUON59240XOANmwvnSnKJP/drFAjBEeSyqCgTLAP6extwgDPgZb4NXZMG+B
hd/Fu5nqjdquT956DKqMy8VQ9XOvzsj9ocD1pMXp9sEDjcgoFhQJN1CAmbCSKBgkEDj7aS0TTouz
sJjGzzS6OKuYHmJKiFEFrVYN9KsQefhMWDRuxUzIc0+oDpJXu0bW4aZDArylnXanWxIpL+n8wiXq
HgJNxhXvZuuevpVGBzrAe+QUJ9EUvc/pJGHTkJxdRpe1L5nF6Y87gwDxFGDNHjvHAXT/vRTSHYJD
Mo9DpEyCq0sjKDEQXVYFPjQZ9QTXujqFhQFuq17dQxm00JFpDc9tfCuOPIhpI7lOWkTfTodfJqnq
hzt3pnjAy2cm5jxZYo4R9UOQcodlSwr8j8z9BJCWr+bpNFTbaYlWRuUgy7cjKa+7EeXliweNmUVu
I+oPHpXr7+LtbnMTfShQgG0XuIdVfP8xydI99tyvGP/1Gggrzy+bvrPZwXWKaLyGmg0nSJ7YekqK
b3amVzokgXiAWMh5SG50Yo1v9paAoMMB/g6P2ZkMwdXUzIlgAqDbBSL3SDuoGqJx1+eYVsecXgep
61RT60O4/PxV3xalxzAxU95Si1dZlMvs2jLQYaYiOXQeqRtKG2Jr/2xXHR2I7higXaTZWhU8sua9
/2bRoZGiViIXbnSMXL7l2TSrshjr5ApSwiV9qEY7k+Hxw+o75W80bZ4qlTtcbSRx/lt0NmVEVvTb
vy9XOEaD73xrNQB6RJrOAPH7nh1WqYaxaUq7y4uKEUYhoojg+kfW2PaDGnvq8sE9v6Q8SbDFMBOV
BNzpFBiFcbtpMrSZE/OREjmSVGUAJdQYHj7frYJ1EFkfNk0eyevRst41zMB895L5SYv+tQwXZ/ng
vA2hVmZUzGHNobCoV8keqBM22ozmSufhPBrwvKCST4a3UvH6CNSz/pL3mVom2FtnGShOlD4kzMQY
CGuYwVSLAeKCnyq+YLUesXbZ/tSh3a8PpusMZ2wyPdmxv+qOnbP/HwfDAASwpHWFgFrliTxjU7Lj
RiYZ0hZ3s1dXghZpLb4UW62X1RpBBzPfaZSts4muO8u6BQx/Mb2jfgtrOykKoK0Y2NnvmS+Yb2Vv
Cggi5OkEcjDM5aaJOdNixX3Rt1PdXDHDCx3QMcc/i+hZ1GKukyAA6CT89E73kun0njAIGMogxuaB
Pb1/y+oCTIMTyzz2vUV9RNxkxBoMHbTSpT/I9xiXjvO/Lh4haPS2GMZydQwsW0cdjVW1mpWHFSAv
/jQoOrXBn7zVuqiOzR8//fDGIspwm8LbdY2UfZOCul2RNZ+DtXelk7uvovKuedHmd4sGjN7cAWCh
SuR82M/NTysYi7UrzJs5n77UBazU4elsmfkDgXvGpa7S/Oa0GE9uDdoWCfInq8sJLCisvjHKHUqf
hL/VLQCXIXI7OYS9bL6K3+XHzMmYSOh734JKgJOoQwKJvGbnMA4+XCDGzVMvonhG8t6gtGSw9v1g
h5l7U3SDxQvgb7h/ASn5yrKRvjmPssMhy/6wAA+wcYJmhjTpTdCft0mW7/riUpfRQx4Mj1NX76Vm
I0wFnaGKVi1V/IMKM6QI+a+iebJTfOuW3G6MnpBFBxcjt4oLJuXMOieFsxRtweRPqad2fM39Nee3
SHWdrvoqonppDNmhpdR3WWFDc8q8zmroRhqlQuCBvKVrxsxF/nqzoXmRtnvlqlP6BkMow+amzu2h
dHc01ae732c6xZ7OKqq7ufUGdC8QplDH+Mvb5AjQFdsO0RVS19iAn8hwcvT66iCkiccTmSxFLGjE
6qmMDGQDGKYoR2XzRNTJIwF/TTO8ei3s7OR0q5+dNFYcWSrV6YcquffIQRKr4CabjIv9dtpuQwop
cmZMXpUPOy3rNGrINNLJtD3QbIIWOHSyZAGaBG2vFetEKg5uglZVM80ziOQlhEFNOfLI7w4H1Edt
k/Uqn3tWETKPHkK4s4DeE7Lqll5LQJ7SVfnDzQ8PCv50u2LSdZmA3jnWPatKqnir70dPPjvhtVfO
tadgooQb70jTMDM2eIx6PfePM3HmhB2C6LF3Dfh2k25XoVVW0h9GNgcdPZPNURAN9HySiGiigVC+
KBkKrX/DoFZIDbBeIkeImMFjKcX9nJEb8R3v5Xx8GTPDesJB5ZdRG9oVGUfhnt5YFwdJtck69h5C
mkVhdkNtxXMyvBV4wE5l76/jAdjDtIuKBBXS/Q6JXym1DzwMiSaK/+hZKAB9s0ec3UYi02dlUToN
8NLaW15AFchEpmANy4xJUVzir7K+/hyc/pSLwUcdI3Hq2pu5BncQid2dbrdg4mfCmHqMyAbx8dzF
Enx2ZGUeZe2pVpUDD0SEbCQZZZzmtZz7b6AZAXriy5lnyyiCwb4+sfeI+Da78tFIhi+9bmsvpB/F
EAXSVqhCvDu1SQjaYGHOznJ78pEXL6WAU01RjThEn1LLyvrdhrlYmU+bVpR1zAr+jP/8vOjFBnah
I23/SrnxQ3LfSIzZgIdBJBDsheCI8ltMrSTVHYwtk6qkuvtEy2xq8BRZG/t5ldQkIjM86V5cqAGp
aM0FP9+oG55c0BMOb+1pBcvuNnlwsKISGkV8dP8DM46vTkz5FGqU6R9Hf72d7QpvCAJQuEFmsDha
Ky24s4vsrh5tPm5M1Q2COegq4VxKM/O9r2kbOQWqq5URmMwTSkyTSk0AjMnElN8QBjdGtipmow3b
T9xiugWqquHBBiyPp+gF4lCr/eMe3J0uU3zdoOekMmO1EuA4oT7dkU6M0cqZgX8OrEN/IGWNEUs6
V8kJyKY4x8Ocuou8sDhsChsKK2okckcIakqeD5mbiIzJUAGfUv0gaVjruWAvED2G5NpaSCZtkS9M
0EyTxeDI1SKb9Vf9TtLHw/iKix0LKMe3igDIomYL1z26hUTHuXps6/MmyRn4IcCSGX7irG7tg+Tm
2cLpMYEV2wBQi8d9Vkzh3S10XPUtSNyC9lFV0kLANlPg2SrtNlKMOg9VKlogosFoQb6WkmhmAaPa
vuWcvOm9745RkgFEbfHXqn3Gz/esTPaHj3hL4dDraswmanmEjOaA3FvCGr1zwDcU0c71I4uNx62f
KWrxJdEdqX7kyQ3jAgjjBHeC9ffi2iKZR0wUkjphYjAdFDeZqNnA7aJ5WeBtkgNz5RcDWXAqqO6n
9XgUFw6DNvg8hI58ML7YVZxSMexOGMLLQLh6BVbazG5c1y3vMXSPOWaSkazLtQkFfE7U+iKMnKhK
S3ZlwZAIYhYK45ApHJh33u2v3Zf0RCDQRJdcEzw8dwS0wIfXBVUbmSHYzviyIz+QRXeuhywd5Qdm
rcIIbXGsEEZbhWDeFAAPHeIZpfp8LeW+KbMX85qM+eqytt0tPVCm914Shwo74pYpW0fi9PdssvuC
/V05LG0fuNOfNbOzws4+3rcH1quo7g6nU+L65eFuhfoqs0BQVoGAYxwVrNy7DsGWPGWbsZf0jecE
z9TcICeNtMBcveI7SMxpagZeuGmYBe0WNEr1EM5JYlmyMPttp0WixzeYx9djoADXReH0tF9fLE5Y
PcgLUs4DRn2Cx2ID3/GkOuBl9XceXR2cdPKGWIMCpatHM/w8dwXUJC6LSamgCZ1b85/d7c0J9l95
copzpd6IqxLW7Ug3AmVlbmCzk0y36eXikMTIWGUB+fx5PxvMdSw8KgdatuSNu7cQtoAqCvI6ZgNa
DCGXQlMH6nCHg7LJNdvVJphYB/flRXIQupJbgp4I05hUywSfkP98YXJWuU8Ui3SmTbwksxAodApO
94Uu4k6EuVit8Bu+mPfFRg1b1v9eG80Pyecnzt0jcTQhMXinNxrfO5NQu2A5IYGFoBjVs+o7ayXG
QRINP7ATYaTJuCmESc82eBYOfBusmM8j1nUJcQ4s5AGVplsJQR3Ahzo7HLa7YBvwT/rZb1TZ5+Hr
dznqJ8Md3hrUG0SIWEwHvBVIaJK4FghhG8SdUi2d7XyQbh4bh1QxHM/GO8UaDNcsbKblifCQ+N6y
cKkdCYc3ftJnTATVOyS0YqByTdM014oJxQkgJVzAKgjoTHN+ub/CzeD99UrhXkvB64W2LYNbcIii
TLTgaEA8cNOUohP5rhYammkglvuWJprczdepvjJKIHIWjHgFwqyBBf1ir3VVf2YtUU3YqmipvdV9
vqe4PDy3O1jF8MP+7N+HSl8c3JhUKU67uAAJ9ec3SJ+F31yL3wUHSxTG3SELzUs39zPy4XFH2lfC
I8vgO82rsTUcC4PoYc4UfrUf8D/pGV5OMtLKQGIqB7g3kTNMVa+tL3voI+4kkyVr/DlLKbOkePo7
OnDHgcueW5d8G7sNy9SpUvU1mgF9tdzLyCQLfZ32CBUjH/07H1t0kH9pDj4OMSm/3NSOPyXBmJwW
JkyMyZfYcyWWMuX96JfBfMJiOkoVROu4FZgYvim+xdr51zhcgZ66mfkz50tmRNsK2fms7FhpbVxP
YrqVxORD0eLSp5Jf8JrU2Yp2CVGKUziTnbLaPh0iWrfAWubYrAEKMzjSUw6bm36UFcHSzNoLf0Z5
wexpNg03Sozh/Smi0GPTmwENshT093lqHCYddMOSgnnH92hNZfwYnhKXYwjgfqUBF2euItlnIAVg
yti8n4cFscixcxjmGVm2GXKKOYWi1YZYizEQkoO0P8aqmswrkMjXd99g6Zl2b3DoKsUdMUqM8l1B
mSENC9jMt2/09IackxjFXortmnXjM5TVTkT0W7nndC27lWidniNQlEUXHkIxMM7sMlnigFlAkcO3
ZCZxNPla2hZmNm5y9dtSLWZ1cUeERklnv2a615U4uL3X5PoMlBsirwqskDLp4L24Iu6XRbUWaodd
3Ex5eFj2MnFj0BSz1t1jB95KE2CxeKi2UVyvkDGt1KMWRwysC2s5G2M9kMqRod0beaKuaSL1rg7X
8dXNMeYJwwBcPfypeImVZMyaqF/stBVPPTkgKqHduyN9pk84nHU+MXo9S7mCMp7LOuVBTZo681Ue
EFOILaZMtXGoR00voCq5WY1NBrDqyQO3YA1NiTlBfhEfWniXDr//wDQxFkU/FgVDdMUcH3TF7D8L
a0S5DL3qSDujF1UjGbz8rX713NpEE4VAWB7A9eBUVE8zE2sdFnOcXUnh5aWec8xUEnc8jsI3IOpr
B0+TA/hl6rZpKJ+xZF18LQwYVmuxPuQwl5oUKGEBOLE+Dix2umcadSt2pWFSKWZc6lLMErk1vn5d
PWK5D5R9auNAC86yZPeoN6Jdt4c9MDbaE6nK/tItJF0C410nWXqQJN4SwvCFZyieU4MAC+jHb5up
TuuxN3+IwdBRq8SBWFVfheHN44yNT89M5j/HApEOCPGlchqOIxbE1CxCh0Z/r28nxSpilMbqTnWj
N6VwqcpJVz70H7sQvNRvmh1SIU0Tdd66urTc81vnCorAk+Oj7qFgEZBq2HDL3WQYp8RWnTviLkmp
Bggq+O2bFv5Hs+oGZWMvVZdipk4lrxunwcJZfKwMpYz5AVIQSbs14a4UnLsv6ewTOfCqCOuoqc4V
CdFsbZ+6VfbMT0kl5xClxvfscGKKS7CbuUvW64F7shvl8ZkSoRHTxPz/eHY6CDXfM/xVnAQkJ8Ih
4x0f5k7ZgMvgZHBCdHZw+5RESlD8184vSnSnnS8X3H68+O1DdMBsdFqZgBpZTyjBrbuP6hAi1ln5
Ww/VL8b/ltG/TjzjK2vosBLlEYGVBamdThr0zkUFTqrtM1dcy6EEwJSslP0PTg8M7sL8p88jD4GV
l/bo46h5XbgP/9IUx2KGZJbmkDv/wL7iqb/TyIsIU1U79e4NrGglERumAW5pd07XIUZjs9uRLNg2
tWY1NnZBgop0T0TbRC229t5aK/DAVAJX8kO86cZTVzmIhWF9T+ryppahLslc/H86Y3TWsOjBuoDU
42JIPlUj2qYE+ZO/OO7u2x3Yp9B9mneBJ+bb6dn8LLItPcr8A29V5SuMVxiCNeGSBgzgCDLN3oSb
9BA10xGaFxna6ah17bYVYFhwRfJSgHpjOBpxkJi5yjE2xfloiS00FGdxiMN9U9mW001gEE1Dx819
94OEEwTizDKeEY5cORI3rCwueI4FzTMzYcpP4t9ojzyPtFVUR38ksdZAF2NsB8Ab+fObxJgJjHZM
CQ6ul8KNcxDZuR0RaQ13V4af9ALc9J0BBvPCHIegvktrLlUJqlOCo+fq4ah9DbqPweCb8qXENJ1l
kGV28dtHoQNIAyy475mKuoCzF96/TZN8lNxE9BhlO4hQCAWdNmOSTa+ibDA+RilW9HYFqfae/YUx
jk7llisYdESJWHx1O5eIHp5iaxOIFa7Nhcs8TNHuK706mwTjrDgxqc2JyLmAHnt02SYacj6vLlDn
x9hxbzhbbCrBr/ckGQ4Amo+7fS8SqHVYLl/Ves4saC16DUtSwpVu81nzoG//K3upB8bO3GV6Ow2Z
z10oAdTZz7WK7qeHPXtrSRQB0vweBkvmVzHDtOen6//MUje3WCdY1tUkMcoTZFN+ZT9extkF6w/9
VKrVwAOf3HvxDs2gmuNpjQU7O5xK4ZeH+V4yFiYC3z5PW66nuN9/lJfFOKFVBs7NKGNt//GT4Uyo
OtQb1/Z/TthbI08QQkz2u8wqw/BN2uxIS/sx8WtjV2g04jt9gITBqC6+1x5+VOGivEsvJBT7O9io
MDRRnfFmfI4e/gcaTxHl6UJx0/rs1sXb3Noo02L5NhMCvnAcDqZouMBc29KYHCfKvUZQ/EiMJQ30
1Uhx+FWpUc0qA1WhY44dKJknAjQi/pnOvBwHIf1+g1hYdkkWVB0P1+cPpreKLThf5/tEH5b8jFec
3T8ILBxgumqsqb6vcb/uWu4/lvIdkIdaAQymnvVztOh91w07BHUYj6JX9iiX+aosN+ek8qC4SeDw
4Dmk62kLgUH7kq0fwmbQ5jkd31SjsHjZiqx+2+9eoDmk8V+6mva/HkZ3zpYMb5Srk7ATe+mITWLW
lDVaNbzY2p6HPZS5oQtA94B+Lo97uPdl6x5RMNZGyu18WhbFARn81iZSYznBtH5GhuwJc5Af5OCZ
PtawbhcUTxdMhRJw5M8aFB57e5CesP6NsHP6fAcO5LDpbiF9QvpE5A1kbRJUy3BvUBreSIc7Sfra
QWNck4O73s+srAuZ3hz/pAyNt1AibUv4pn+FGs76hG+/n81yL4wN563XjEDb2U5QNAK+eoqcPI1l
4ZcHcGWHvu+JlrRbQl0gxQxtOzHPTg6OlyhGYEQfdw21JQipwiRYdE2YfbsIcP/WaR4Ra5nip+VN
HJ9+FoWfDiwEpqvsMdJVnh5xjUFhL1WMnmtfjEKpeol0MgwfNm4Ky78Eqp0wohYMoxfjSnbbENp6
AeB7nTv/ZD+JvGRDYqWDvBJgiqX6+cLW6AeLNHwvDiPq2g2zdnYa/FigS4Ka9HinwpRnA1dGdwBS
uqmu8WCLwdCxCsJEov4sqg9yGKAqahUlfgP2MT52Qx9qSlgOcc0yn07+AoVarVWa6ouFCYTus9om
fevUrvkW4SDg6YzXo5cj3AbhM4OOmADKJfqem23SrHMBNTHWcOdDYKG9KQ5VWFzzRjbGgnsBgprN
PgEZcm3Q/OXSiuKvyjWfs0YNihyyHfb5pjSMK3pvu/scehbVD5vUKNPl3KhPJeSo0vgoaX4dcQcH
8W0k7pVCm9GJWbyOIvp9u1nydmGqo7G4zuU4rfvMudOYAz+yXA1YA7PGxHsqa+yazcrRJ+YMy27t
Vm6p5ftVwi9PcWiSSsd/NA4r568xGUx/DRmzLuKQ3W6V87WOH8oI1UNFFmm69VGGoYoGOOeL+wlV
fcd+UfaugkJKngv1rld2ovz9DO2+klSJAk1nePWuJLol5lz6aNGr6oXl4gwe+6c7zfB6DpRN8edF
SgNnebEMM4G7Jp0ML+MmQ03idYffDw/ZrLl6sinfCtzl7gYlF1BjhpILJowfQ6W4D/0Vs2MTFXhN
pxF5IbSgoQ40v97Vc66dCwV7dt+DFivdB1Q88GkFhkZaK1afyV6UhVRGTw5ylTlWoVChPsdB9ywg
fwZXZFt/tEt+re9XqiLGeU36e6rIARLwfCZN4w8/tOKSoCQnGCYZfDHorM5N4mprfcx2GAW+JGVB
h9dTqRsq8sMtQOTFnkKNYcbx1Bk+HpJnkxywA8RYLW9hZDgKHbD0sJ/IGLF5+Wk/qZ2hU89XU2A8
Z62PH5+VrDyZOQ1s91NNB52DJvIS7qfltdLqeGuCyZbZxRog0Z+JhVTbZBHi1Ieo7OjZscXbuid+
ze6mFILJCJefBI8thtu9i+inYO422iW9rXBfJpQC8/G/3AtWy6zFGsCMy003D0G8zuCDiqsm9nYG
3cfpxxqf0eHGwGBIyl6FghflISPETTzDWdqnjFIFPeSVh+5zhUmEYAC3QV/2GIDZkdzS9Xl4mKfD
2SwMzMZhmO4VbtJ56aE/It6JzWmM0z+enW1pwhAAWpPRbPEOBTdqN8RNfnxTtGaHEQ2N3j2DQ/cv
VsQuJKfHLLWDQZwBnCxJC9Gnrmy4VHD8Raoyj1cJhG9Q89wd01grvPGvPfDhgOj3oHRDfBYnCC82
kMBCl+RJolOPOZhaqoI4WTm5Ay4h/aXhx4gZRCp5H6yEgs82StLqSQyZJXvEokrMEXsQ+wd1P8Xg
TZIi0aBy5M1aNB81AT+pST1sHoKIZ8znCD6BiGj7hRnF1wwFlx2FjEF5iGl+KOt8th1tIH3FbSDY
YSJqsHK1LuXfh3sXOauLyNYMAqwE+8KNY6skl+V+YeRjqIfSrCK1mndQJ8toydXTka1xSbFykDKg
0LSp/Db5VopOKbopxQ7X3fKhd3S/XLRlTMpGqJvQs9/vzgZ95xl3Jh8xuT43hOC4gvxBFxj2jzQP
rRC6hGmR9Gq6NNPCoEVpNMp9YyGYWqFSe3rqmMl7HaHDYVeLKSC9mHceH5uq0JQ/yIdT86muLzPR
jRgW57HRH4IAKgHhBh/Y/nbs8tlkQUrvMVFy9sNFrbQJHp7mcXIf9ZzJnXS6LGZXuW1SndEZ/7HG
xMzP/8wF7j7vZomZPLEA9MSa4NvSuo/8xaY7IvVjpjQNX+XA5jg6kdrrhnwzDrf6dexPXo3QKmBf
5qpOukJS+dZvTT0olji/LxtlFkzTOj0/oKUKLIZr3TlN7O0mef6vUk8k4oviVb8kWKeD+1XZYV76
V2b0ctz2nTGqNo1M7LMlD47JT3uZkR/XppD1e+bbFhEjttK07sMGkRvszzep2PZMUsDXJMx5MShK
DlGimIRd2DgubbbihaL9DFCTLh/uIqbNIsc8o+8gHNoOjl/z9DWE8wBHZttnHx9tDhQVIY3JYP7U
81Jp9ucDKyGMJOUkGV7S8kwEv5BFG6zAHacID8Zg7YrBcChTM6FtHmj5XrsW9vjRYqD4wWpVKTkn
r2q4uy9Aa/4Zcy6nb2rU46EPdCiPuK52ES9O6W7RE5M/8IjJIc+jLMJGf1FXv7DwokAnQE3+xOot
tlKeSGa/1PstcIPUxZK4tRDLfxTOLI+toC4CDN1ukM0barklnlGZmK0JLj98kMkqz135sK9Q4qxA
vBneVlTWTDJiPnHM4jU1cvxzbLYr1nlDitwErvVReXgrpvLsJR+1GDyuL+Evyk3qOGRjVKdKbEBw
PoX1GGnEIOAry6ziWm6tI1WeyOcI/VQJtMBuerwDQxlbx+ZvKB20bX07hCUQugQ/FUFEsCtzD2bY
nbHnJYgc9YDUG3S8pU8k9dt7N299NSXeIWzc934TScP1x6Dot2LvBQ9OqTDnUfZ0ERVdCwtuo5mZ
Sq9klZMigBe3P1J6izdCUpiPgP4zOJ2DQlr+1LFY7RcN1Ydh/pQyVkNQuuv0fwkdH/r7WVGuNKE/
xO2jsx+uy2iFWTibuWAOQaAFvjaYH3QQEytEC9GH4RDR5fglpytfoAJDiXbQ/+yT/vCu4BJqjTZ6
L3ArilT0+aIlqPkLwqMKI2UF3B8EhS2WPLFtdVrr2xI9W9ExM7IwbeXxqlgGkzikfs+7vMKzTIUI
DTLVQIEIgBfhpuySTjJ4f4GEfiPFlfACYD1nofr3+vpuHmG2AHFL8aTSV/dYKLV0tpSG+UPVsS5B
kC/L4RDW5Cy0x4NxxyeYyvHiq+DNmE6dH5noe/Rr/9T/acsPfZve0yICJHusemnIOeSTvKPu++eC
xRsDpCq/PJKTN/m8IH++beOd40I74sLLSKdJoas3RO4qPcs+E0Yd8Xn2rCvBMzVE64qrMKfbEDCA
qJld5VKVIB8vhnnqnjVsKLYzoPDlrywtRT/IGejRbMI4dtGSJBBzWCdd2bTyOFrfbqWZ5zV2d+6Y
t2Zw0FRfS7n+1xR//ZCU6Md3wf16ceXwNVA/gtVLllpvM5dAlInNynwD+YneWop6XprU0LKA75ld
Xyh0kA5Nb2IzfqFtyleTWIuNzwEa4uqJWFjNAnaGOiykVoTRiVHR0VtxkiPxVc6OPR5cTJHsuBhK
Ymg876wtGLwmVMAwU0yzytAuWsEcXq5/L/lYQTCXi230Q6n6ooPsEfHXizhdp3vCc3LnRjyIl6iq
zMKQD5HqAzSeIz0P6ACqaTpTmoAxSVUvH/nMG9uajhNmqxWrEG/fn4C3/l8sagOgX/oey7I9wicM
LMuEeOXVboIdQ909WQ4hAzFRaKON+rOljOFWIJ4WQ+zOXjhkdos7CyfZYKWGRjc3Qd9LkovgQnZK
gCB6S58Bfu+8I4r4oFfuPDWwn5qpDkN2hTFXPEXtpiTx+y5qFFVlpG0XgfEmcPYTY02xNaBQi3mt
z9qP1S69M5U8Q7tiKXoxjJ+/+YP9COhP2cCv6reRCj8fHisp87fgmbyidtXTulNom7MdLvkplLm0
9J5WXSKNkok7pthvp+5YHgF5Fp1DjMjUATNMc43+Tkd3GUT8Yl+U91/zZijXlu1ImeeRQJWQWBw8
VgpR7HmgKauJOBvtcSwkQFVtDs5yKkThlBe1hBUpdm7c5qURo62Fm9TlL/ICZsaJcMXEdko2ogaJ
cd8WhPrwc2i9PozghOKgGx4cz3IEAHNrHJrP6BoY9UooGEZGwo2I/RZCg87FArxCXdqR4ycyr5+q
hJdJLkAkeVBhwtnLtnPMkU0wYdJV8g6okXoe/UW3B3rVMs0bToft1fPqP8TrTsiiCpIvkuKrJJ6B
seOGeRd9dYWms45SJPFIf86eXYnj6FhGhr8MCEOch2HIUl3qmxYKDZGxgFHQvp/B3lmY9+UL/zPC
UBJwvm5pXVdEJpw2Xm44Tj3bk45rHcWbaeYD8AUSUhz4MBovERMIPpPjciH4YjTcwSmX8H/pcnLv
Zz52UkUkKmmF/GWhUup7bObM0Ca+JfLDJd3eBxVRPvX84yJmNz7iHHLFSEWfHxo7cPQkH3pw8/jc
gh13sM4dAKxPLaLeAoD5u1bwFGqvu5WIukzTzEY1hCNIT1/O5oe2sR2Woto10lJnc0nMWx08ADvl
IUAaNxdAcnTzmAfociJ+7gW4jXDJ/KKKm8HXrelRfK+PI/SLGjVgyH0eoqdK5vbMzJi35itSZDL8
ZzcaydLzrzUCG/M5njWRwUIFenByLjzmus6CLboo1EtzkuZDm85LCMPElXq5OY6y2J6J8FXMNQug
J78Ia6aRPDbpJI2Vbu3ayW7r0jC0KkD5SWcMvll0S/+6tZlgmU7ttQ3gBRlrH7Cah91T5PAsyS5v
I66M/aJ3QS20a116id8wUkTYnbN+RBWYMiaM9T7qi24Pe7kDaUSz6wK395LBdCxB1xEnHXJUEygL
zyYpZLyWlaC6HIL8h3N7nOvfCSTnuxVzuz97d+61d0gJrlIeCqnZiBWFn9xeFAu/rC4EV5J2cB4y
8f+PcLYMtmYFiCtww3CU59Lt2BvY3W2ZV8Uh3pUM/bFvOHtFB2yd4OFLYHcyO/ZItwrOBkhjP/iW
3pA9UlcsnW12KiByknX8+tcuRJ734xb/PRnbB6uR+eXvnFeBHaAg3AGkiEWV+/E6YfRm6FzVgBwS
JTOPmSLD9TWySFhmEZOBnCoP4DKOFfSudZ2R/6RlzNRGBlpsBMM097sQsGbbVJ1kGYvMN5AShCX7
M4luFPHGD5XNOdwF6En0QBrFENaAfuzHY67grjmJUiNPvhOuvp1jC06ays0PFoFR6tgHZ2MhQfIx
uH96sWAAOas8AJd/XhifsXUUNxHIx9PXgyJuu930Jpfhdak7lwJ4P3ms+UJuEEZBYtEqhL0QUX+K
iGoimDAoV5G5TD2UOyy/OYNz94RbbXM2EkTW0RlpnSKNPvGhHkQ7zfH9rCwSP71ZsO6yMT8TLn87
hbfIbZjlul9DlIMwKF15bRn1Y4fuZsD3Kq06V1+pSAjjwdudWARASI71v0xxRr1NXqI3F7aMZHB9
D+Q3m+YBZvmFrgJL4N3hb8nzm/aJwJS/KQqw2a5Ghryz3VpWO95DRIAE42UkNA+PjOdmFJ8YQZSU
hM8UWWKwNZvMGcp2M/iJ825YPXsBhvSzmTfpnHBmq1Y4KYpVS6CXM6zeLwo1X3JkFjMoGx1pbunz
8noz81o7I+kiRnvKRfl0Hpfwrgr5iQCamhaQBoGclvmkQq5zxc3bS3UAgXWfB59eddHxQguQG6HO
m+ZKmTcsLB1vxe7pion+1e6aXS7hSSdYD3o3Ey/CGLU8DuFzLIzzeyDQY328QeUJd4M/kexuXA0p
AtmhSb9ZD8CqE4wt4OT1GmvUQeSC2YzDQkYT0mmKXQx88RWc9mqbDJrRVSwVLoPtiBaFGXtHBLyS
l2d/nbW/rIeMkYzglxqEduM9jjH5J8gsZpIHwXO6UypKN2ulXayufh5cJbDsPjmUL7pfmZJ7Jfpz
kjb9UQNegT4C2XKupIF95A2+wfcZYTWcvSFFOljkpNC3FoMaIfPeN/SOXuRpOl4AM+dwwO6f7U34
ZmpjXwQuGYRwK9H50JFtdl0UQaaIQ+sW9TYfRrBFB7ZA+lmy8X6JnrYBrvkyqab0XZBZedV7jj1a
r/x5pLxA2HSIZv2SA0DR0c+ithsRo98Cusyt86mwjDPgnGO5zTg1ff7KbH8n7JpEQs1GvEJY0fII
DLHqjUSIY/UZyocHr3qm/nlDJpSmosmEd4T0ZOHYBS27N4X+gvMDXerAixSuIAx8a6UW+HOy0OaP
CVIULvYj3BMk0bfJinpjAqAUZ80dWRmDs/a1N2H0ulVf+jYqjfLNbxQ3CpDiL2I4Kqm1vly4yYjN
qsfxhicvlZTVgVXY/1bwbp559b7CT391GH1Fv79xcXjwAM0DuQR7Sd3FSU7hB5+9vTo9Z1vNcwns
6E1+rabM+fZCsuIjAbvjAIiRrB/23jP2fPalVU/TU7PSYSB37RTrQMsAYx4IEmXLPUWIA4NpNPGy
paZM9A+Io+eTqLwxJIBuryDuYij8QIK/uzaH/I+KtCpgg1HTNEX66gccT1yfXD1lzhnGMKLkR0bt
b2untx6VKDYsm/IKC8ajyUJINVVjCOfdYWpeu+uzrC1vVGfT0xKmlLyCpktYB+hMrDUfIOXn9K0w
0pmisrK3OiC2VNg9JO2+xF64k64tK1L+Ua78Twq70qTtGEl+Tobm7Ll3f6tv8FB/c4ClGGcuOElH
X9xkmN6gN1nambzqKW35op/jc6A4IN6YGJa9JBfe5IIhwnmNTAiA6h9YWRswLbNHWpZGHxoVmJ5y
Nn1j2X+asSLY7qadWNXaCw8GDv6cfjcQHv9LkR0Ld9G6vZjIKbSO+8iUQaGWSZCwAGYXPH7WPKIi
ivWD0KsykzGN94Ef53t4b+mXeScK9L5SFRpgPQGwZSKqHcpHjcPBM649vCVf6z/ZGeJN2ezxt/pM
jBGeQSKTDvtIe6fos6X8oCHKdHhexb6xj078cAtDr0zRGqhHKj59YJfFpALAuFbMUbaGUR4htDY1
e0sMAWly7MY87VeP/uw8hxi5BBQXXi718jiYMUBhLYHPePwEjIqNkJMfOqTeYsC8jwYkqf5pfRxk
/Sps3N+WMBMipIzOUzAlbEEvb9e1TepxdFnW4wO/4e7aksvHoXKKXZLOCqyxjmiUjjjdxZn9OcUf
G1KE30mj6d+mwJhydZWxDfBnsOPOmFhYUkdY/5GJmH5qUyOkulQYeFzoJ2CQ46CfKfApojxAWDcb
nGRXO4gcMZ0nVaVV902Vcoj0fGqEEEmVvbn5282fUTGlUvtQPObUH0Vi93Uj6UTmqEsHhzB5ow5l
VmYZdXN7ipOXPVqt8cSENH0Fsgy7DAZCQIxHAQsKxWTtEnFUXBWKI8QuzSzXgueiqt1Hy4DeQrIn
pcjgSn5w6QApU5ywJ7vmqqTrqdo5jwnzVj+m6PugoOdNtuJx6zHXQJN3wgKVC1m6+0ElJtfHG4T1
vJ/EkH8+CLCQTtz2Ig9vG5FH9DjPEF1Aakupcm5SvMK+S0rE1VyvRw0at5NM8n4fjyIU5+Oz0u4L
dyvF8vp8f9twY4+bQeUc5CyWRpPEDhQEB9h6Wiu1HIgaWZoL/bOS8zboywTyJEwVwGo5kmK/RzLN
BgBFylVUPlSUEEwWVBCkCxxAbxjwB6tgQ7rXl2lGqXSuWSrv0XeOdZmhFZM5tjbfcX6v5qZYBrCP
sg7Gy+6WQCQETnWMZJMy8vfVi79RD9fv5E9xFKlTBzwYkVvAEY+9mRkOJbUvCk/WoTEQyUclPns9
uLt4RfUTBvE9JnCarCRbRax6POPhvgXLj6VqIaCI5qN2UB2li5ePfuJeG3W77V+j5TRX39LfY9Lf
sqNkloT5phzr6vcpTY5JcMDY+xzXa8Gd3oVoKcwTOVPVkY6wIdUR7ZocRbzZp5IMQBb7872xih+P
UOseIuykKkSldWzP5e767nqVZHfYWMvTTfA0YoNdT/CBovUDdhwTKxRpnkz4sncGfQHcIoTQk+Xd
k+31ClkAkJyCRb+qUqTA03ASXnvj6Z06JQu7RNbXypk5E1ByMXISzB5RcZ6MLfjxMH1VyCh6xXlY
YwdpFAbKs7DCleGtBbL9LD0qM1xAcIqULH3eIlrSF44/CSTYg93p0s6WSgaPIoL804SN3gZ8cATo
xw5TprKiwZ1oSqWdsfbS8YwCMCEPvVvSGRfECmPphY+HNQcvgJE9qhoCHG+vxytfYFmuHGrGBzQK
uQQZlaAixR9wP+SamIU0V6tMSjHM4F73N+HzywSs02X+qRrWKznBUq8IchFgKcZAwsNkMnSeVkwz
+g+bAri+o2xRJz1MThpiNNkULWnwthc0TAaJ9fCtyx8GIo0tZ/mZ19XZEUux2EZrgoUZVKB/toA9
skIwVHDL4ISveZULPHRtU8btsNicPYkTXPseud6bejuY3f9J85jRCdoYbOw9CUxt8mNVIUn3rnNm
eZveZ8jBFKJXO/zEMZGImh0SY96jaoW+9NegMiWXic1VS0FpPv6c87IElEu7vNYL6pZLwYOp+9TQ
FiVmr3QRYShESf3f3YaW7rMtTvFwH71wvKp6HsyoKmRjlpBUirAPc3s04MM/gv2VmLzxE1NXwtRq
DPOE3WAVF7bFs0QWP59TcNn9DNJsPc0JTNVdNdIJRmimNWH8H0fvwY9SPQWEts5H3BGvpg//A7hX
kEpCA7epq4fesynM+r69ZS/lWbgsqUK85Ki0QOmlhWP5KfZjS7qH5zdeqK+xaqzWvHnMmkScmp7k
aeN37u2ME0W2h6HSaGtlG+j01sJhVa2uDGi2jhC1lqprmZJW3c5G88PPj1PihpbROlGgOTaT24p4
r0t0KMk4hAF1xjj4y/5jZ0h8+SDvj56KSAoaEVHGmxBx6mFJTsCCUGVr2lXfXuBuMkbSg8TV6dMF
J8a60i3IlIQ9ctJPy2+i1i1LfUsE2PD4jlI5CXIwQGnz9tLZ1Ym43oWBI6nFfNJVcOZmx6KKWd4d
HTt2borCWwkb9MAe2QO7wtto7Vx6cBDG2GZr4Ja6etycr246AC4DaBEvNGGXNK00khXgGVGAg68k
nMqdsF4wMjng1I2dAhNH5DDzYxWsn3l7wZcDDtWw+Y1ahtoHW3ZTuhLGillg1/bgAzX6jNqDHYDL
IwMY9sZx6iSkVlN6EkQ1ZHWpzgMZWyccacCxPIji+Sc3VRG7+Rjtq1rXxCXuzPd0h9oY+CjCH7w5
6EG8jR9BcAc33ZWJ2XyzOk/MZi1t0RtOhoQjOEzIGUCfyDX6XJIGlpatkLOBVAMzaFRyZzGYDe/5
RQXx3SQVI3xMo9Vb36uZPRbmVXf8eHABfJD7z6PdKYtbHpNdlicyyN/RgWOJTLO8hL/e/FPrUPG1
vafYMiO1UlPfB1CtmTOeWAcZt/Mpeoi0aLRhN4Z4IAaOw5MAPNH7m1EvF3kazeqyCHBLbTadINKx
sb4EMgs7SOdYfnlqFzdvMqxoRMM20zXJ3S0n8/q7d02ckcoyOUE22esNTBPsLiATRPxJvVD+gkU7
iErj2q4fi1ADq5ClGzuk1LvWbpwVU6tbu5yiwgCgaUvvc8KWhkDvqNkJrRQBpyy+0OgYZOQJaP6o
ouGkCOw/mj1vESWB+QnsfFLr6tH1b49x3bmiqfycxUfBrwg8PU8H2F1MeHvd2wlGrhUnsJgk1vAt
oQ3KBUNw7O10SfhdHKoxb6snPQ812yYasW+reT1EVj+xZlNkuyHpqV7hA7DtLIwYdifd2/dGA3D6
5/mZbuUYryC5Io7aFQsoBbB9LHDLd5k/HOAzFDg1U5wPuU9JsZukZ1MvzjUGG0ZBvwDppPqytTQM
OxrVtc8c9IW4HQq0E10YHrNAv1uEPw/ewrydi1bUCbHYFqWbc0DRZZFKmamV3IBQWXd855vL2Ztk
33m3mucfAY5BSA+ojfqLJH9coCZuVwU87XSrPUpVlP76o5VN3nYkUajElTaE2Rkx5bPWkQN/nmjc
c9D/AFVxwkvKcZHjAPak5bqIwL1bDiysoVionjhHtW4VYP/NtT2MkS/i6GX4OCdBMI1mRTT6fmWG
uCzzPOSZaAp14b9fcPq75ytQdRTFENYzu+aSJp4un33zrejLRpxqtdJbsIcmSQDChxQRGQPyk7MP
i6r6Ost4EjrG0uwnAsRwHfEszrgVPKuhhdI/kY3v8wT/wGJp+JvUA1g4mjeSu1NXVkiGuieUA6gR
aT80xQT7VeQ0JhMA00sgQUk70TcRtX3Q+Qf3jP8cvyXSgWGJjH38/EhnDGnzZkxgZfJMMNUbQESl
TO+6hrN7fe6+CYD/yXaYNPYCMkeYI056ns5syOL+JM27ouxyKHZrflqbTeoiEe0iYOQplGmqx7X7
vvUOlqPvu2e7F8PK3d0gGsUJw97VAYxye8t2dl/8/pb/oGad1PKOnTlu+DGPoacwHNXyhG6A2A4K
ZOs6C4fXLm9etC3q3BH6W5BoeGy2ouJv5bFxPtU9QlT9cKC/OwJf+IMR1PBdzY3NWN0AHV9Dj3bs
Rzkk7gyaLVmb90dAKn7Ltsa5CKbOeGuKGeXe+x6fXZ9nYJAiORXhmsViO06j24Z7d42fLgYLfmGW
//z6Ss8hkTZQHAtsItGRbsxLvxxiZdgN8ebE5vXj6uZFNPik2kUhuStQv1dP9fiGp6/GqQkur+k6
s+YSq05/KqIpE36rOd9yBZLBFdmDO9LRy3nQtHN4qlBFBfrPtUAuTXD2FND+8IaxJaIZ5IfasF/l
XRT2Ecghydpm3WtQ0jYMi7Ec6CCpXa1gN/Zotuhy6kHNrW69zsycjw5H/viWk/+sJ6aP9iTuBXwG
L1zfeS8ZNib2X/dnfD2Cdi2WS1dEPjD6vTSW+Is8yV+GOTjTm3VZ9Y6TkCcx/FkY4P3jtZHngxLq
CN1net/ypDPtjLDluNHaeTlky1JCHF0sPOAO10/MNzsxy2W5HjKD1HijM81/1K2rPVOuTfJuYXEt
tk97dVn9UQuNQUVnE5PDxGt4QMlvzCjTIgcCXDo4DVYaIXP6XRyfAGvF6HrycIF1u3P6VstaPofp
/owdSCsEQY+Dx5SinOAKoDj3uaePLGzd2PQtiB6OT2zdaCzB7hIc1yM30ODdUxEjsMiuMP04uz+T
iq4kcjFKMz7taA2zuxLYzk/6haZhjwLrg0/LspKI5h0rqO5OORfiZzS7f/AcRxoDKZfG2CAKt5NF
ZByNcSSO7J2o10Hr/FV5WcvKGwxwb4ygGIbFX99swVWH5nvgXDFYng/KNn4IaBo2MxsWAXmy6X3v
nzCH31rIXz71dWHR8jod6zHxpG0En8wEfXkpxtItY6Kaq7semqrnRwApVbNynE6OUkfjM/9Zvrvi
nR4R3j6bkvx+FvjNmWPjSIO+BFG+vagnHIZX0uIv7aH+TMtgpGgemBFFRyVOFxv2VgDwCVB7EpNO
wvu3i8Fw/g+u9HW5Wwe6/yPQnJaTRE7J5G53fqA11ljxkEZHuXVDWLVA5Du0d136zgOxIIei/1Rh
PpLUJ2jR6TtzXtcwXkgt5GTk3nGX+e0fI9Owp3zdqN0r7acmbWcU6UkAaLZg67Uz4BMTECRQWUVv
K/tB8GV//nJg3988ZQlqGLVG31mP0urQ1IMIcfxJxBH0QYh/KJ1w/b57LTR2N2ihKXzUq78lTAdv
qdqurVX8d1QyCylqaHtQmFLhcrHl6Y6B2CwXjeI9YVJcp6+ocX6maIqXjw1UOU9iH5LuzvpgxeW8
iOEGuFcDlCqPG784ibdin0PQph6l2JdxPQZOIbYV/J8uSdVqTTZXFo0KiaxQWhAA8pNqlMvKKGnf
4hfr6zsHMW5XyD1kzwJ/SdUXo3yjnoLUiZTfs2ofdGVS6yRgOPNMbs/Y7xP8wwrNVZh4LR1TdC32
M3uPlrmbCybsH58XEpllNHEtpcmrMYMX8n5US3GQj5QDLVaHgJdpN4v5GGxJPIhaR1mjlbHmWsOe
dN8tsiOcf8U+0M9ghzvTBT8y9OUrWL+unrsdiQO83uiJZdAK1mjMx4gispmyFZt968IvV/CrJhWo
8bzHzVPj0bkaqh8RXyvGNZgNUVQSOgbGPEr+7tShUvgnlVnaFQ/TM93oDCItCBIZ2b6O2MDwHxUH
nK7eVppk7UR1u5be7k9VeIx6f60svzvTt25oJesKtQZQUITsEBy7e99Z6rlculeQZs3vJcqLjzpp
4HfrPdWEGPkMz3ohXKTZBkObi9CZjlhoSmKoG25+i4U9e3f2nCcbFjIc2AgcKpN4ZwQt/MCrYv/N
DfgnkqDA5C/WD9f8nRQl11Fa7f+LBPlQG5f7HrlwAL1nLhn0Y/huuitQOe6OtkVpB5KE/da0sbTV
bT0ErEILh8tNuEEXQKjRhxrzM4Zdo/SpYrsP4byZmMa/KkvLMWapm1ltfQQ4Z/0NLpXf2PVpZ1/O
u4mvK8Mney0XrgU+TmD432e7fD78Wkl/ySAPgkI/oJEPZp85HpKkf4azxWDiODlLEXc6RMNBE4tt
TNnx64dEoncgFs6Lm+3XSj6tXtI+RFAWV2cpIndHkY0Ofa/i6JnVQtzG/AYr18iXagH4q+il9iQJ
34ulidlNUaX3ogTDgkvzP14oXjW31kgMyePfoV/cPc5V+QwdMzLUhR6d1KDJlP8UIk3R4zfb3694
nNhZTD06gVHjX/xwD0N5Y0cxqRMAJmY3AlfZjPe3T1amtNv6wevBLVFJecAVh5QhwM/RMhEbebp4
ioIkLE1+ckzxgq7fsDoj7pg9YcHPnR2MG17ntlNxL32BCE1ZJMUY/N9K8msE2gYcB0T1WnDaeIW4
UifDVIvuD4RszCpFrnHUOTMa4lFnDfPg0qRBNW8FE/GiEQU5dLkfMIQRN+q++jKoO6LzulhjvSQf
SnlgF5mRNIYWAcBGW1CSmfidOXyO2PkDV2JdyqY5yIKplPIB3qliQvSvK5JYg4Fu+SITstoXJuk4
hmJcm5KswI5iEQWjNckY40y+L0JW/0ivTBh8cSscmkthHUIkQW89nXYJ8DCbneD0cnCb/5hYPUR/
KZTY3UV31ghDbwRKwNMP7fEDYOgHaHCUd4Lnx7BQ8o398XPsYJco/Qdp2F0KJngfWX1JOGC26kY3
A19cY27kxY2BAtE346CCBQq6ni/I9uN5vPBtSTIVoFrCeK4cn++yv+oFKmMjbrzzYlBHrlLrF23w
gxIOcWbmR//60ld0V14j5E/c53bT7AtqLkoEg+COZf6JGimkHqyostiz1sxx2BOjJw2bDnTf37Wf
764vZQ/+3v2WCvUEpefjSDo6dG+vSJWc3oOoY3nPsICh4nMAEUBVf7XcqLK6YwMz5AYvPs+yVVQw
R9eA+OAWohO3CYkJKAgu0XVsXOpbOV54HRHEvRGLtFvrYcZQrF2xXkQyAk1PwOJlKfijWEQwt8OL
p+pO6KqbOl1L2TB+nYSLpJBueuT37uTSoadySYmmvcn/e/Tla7mKGbNTTS9fseFMtvuM+Pt9UKsi
/TKHzjlc4/t1SlwFSyfPHIRhAKAWyD8j8GvH7Q85564ncvVqPo62zbfJW5WGqOUBg9x45hvdHgX3
oOTOMIsIbuqhZEviN9Qc6V1hAo7hAAae82rtWpYaY8Y0TNqn9M5JG5wFP2P0nzlgKFd+WyfwZ1WG
vh5r/cvsmq8WcQO2tPGIpNvl+YSonkZQPAPSPJU3+41rHq0Z3ECMYfhaiZlzS2UVTB1qNNrZixHQ
tMYuHrTrZkHaARraYBneZ/A5T8FAhwDXaUsX+UoNXVg+xZtVqeSmVb1pPfu9ALp0iNdzz7sQ2zh8
5GiA1p0smXodW+f3ruFsIY2VvMDlCp5ntWUC8ITw0mUfn0XLx+JY5fdHNk6I2rg1LGkxZKOI3xME
fdT8c4AnBcW2eRkRFb/dSFIGNgt4pJQa+3EFnItiCyOjdq2uOd6L9jisGwhIH4W5Xyf8+FvjNCfy
MHKR6wXgkmPoeZhSiHAxDdPWHo/kwqLZ3Dyp0cpEZ8cS0DmBeVohlMG33h2o4f+RSO/19RorRlqW
4jpP6lOHcAtYJoq1fiCaNZEUKF3vVf19kPs6YgQNinSvDNifaGA8tttTEOVSRofwqnRkDmEsLcyF
KtaIHcnpjyZQqr/v37qpePu7zesN2f0OoRnZTL5FGA63i8R0yvOnC9a+50yOkX7ROrf39yFSgoOI
4OeEKcfCVADIqH4IG1BiGH47WLoUGfOQOdVh2zmnn7PDN2+Xp8kBfSfIBdXE50MwNr0mBP83pwCL
pZtTSq1nQXo9Mt7A1QzpAqcgRSl084bbq9W8+E5jUtklUYVci7pYJpk/M2hmtS6Cuuy+8f166SOo
I/jyJaP7WxRvCUPfO3WexIfOetoappZO5xO9THzrsEbyTjFCEwC26phcV5tGlXC8o/3p3Ln4S6Bd
eSgXHdQjqWUvMT6kzq37fZGZsjSUVuSXSxG/SU3gNukH1hzZFdQ9G/8KPSBOmA9of/UQCbPtMT3W
TijtHer5O1zy6YK8a9uIk04Bzruxg++0nvFDUhNxqqZqMNJDxsPMj1N3ZZve5x2NdKSsgJrpO1Wq
xnzf8/UJS5h8C32qUYJIVrV/nguuiViltUw4wvpFFU7u7zHLuBwz+aSMW4wEGTCSKqALNO1T5eyq
v8208Ck391CQuXYzIhiXfgNuOSRVXBoqB61hx2JAEezafZ8bMayRzXIj3lOPF277QzTY27l059wC
3KvCkjYyIuMlrQbNqZ3f3hcsEJ8hSZ2UpcItocI3cFcJ80oHzs3omNVBYyJK8Z+vOOxjmNVy9qIy
rnLTwx6ocwurAEUOoVkUINH83gCjoX5HN5oOGXJKQ/e9SfOQvJ9AGO85m37kawYIZ2Rw6mcttLl+
UJTzKLBQFgDsME9bXNQmHRt8tpPcNqkEWzR7gCxbuOIExRavBvpWiiDuptB21iM9XIr/z03UGpVK
3zA6mqBAHwPvHl6Q2pnBIuzrY8DwtxqbkDZcUID5GRtJCP8zT3n8iYg7KaE1HpHo26FMaDkF6Bxi
rzmjni2fCfEFFmr8PaO2ynzAqhddbwBGvIu1pB4r58o/Hi6f2zP6hLUAFb7ZwM/WC4+Q2hsLGOQC
pptt61FpMaMMJvXPuDmQtCpGxyoAacIlyUxgXVKJIYaXpCTBVXNZorTYzaDk29YeOoyf1IqCnPDt
vVmxEl24znNKpl/7MhTQ5IIHKBm5pPq9XAb0gnbdx9xKPHbFI7MX3wvza5dGKisP2U8Ly92fjsyY
hT1uvw4Ia7morrebBx8GV/kMsyiUiPoXtJM9e90kUwoMf2RYW4gcmbr6SjsuWwJDXtdrnA5xXN92
4LgO1/KuIaEB5KkE9hEnuGdesSRoHtdO4tLtPGWPC71bEnKhKGZP4pJ+V82UkjrdV1xIE3+FwP5+
lm0yMK5Cx1iMraxm4t3eNzDXqjIgitRvDih+G/zShME79vNDOweyHXy/k/YNi4QSpRN9xzTAkAkI
QwrzSQIEmGsEQZgCcw1MgbtLR6Gon9Zy88m5I6I2MLbTWCvbU0cGP+F/aH8BYVly2q3OFeyXnuE6
ysXZ+awF1AiTowJ0FYTJHduISgtsF4cm+noF4F8sKANz+9/rSroFnsmNt87Zw6Pj4TwVi1zvlb3y
jfrFfClRcG5MKgGrByS9kSb0Mir554A280Xf6jFgszxSUu3/hdRmbMvrjV0YByKCCLuY1pualUNR
WTiKEhFYd/2voNzQRRlXRbt3XiuT9YAplSPK7cR8839J7Ah+549iKmeDIj7OdRy++cfUXH4A/It9
OIqiqzi1oGLkTcb3/Iuj3iINHz4qcp7NBuLR4M6CQkqRvdFK08xz4gkYHz3v4ozbIgRZnT4QAsqi
OzYZtI8l7ZFj/SCQYJ6h8IC0ogsVt3W/senk8Qlglj1pqxvsrHctJtmBfYvCjSt2WJODL6loiI2j
5POABuxBZBek434xydwA5laPCALRgKPX3oJWfSaFm+XkruH6e6GrOoiNwb4L0FnGVyadYhFpslmn
dwKBkuh+WqE6UKjrltAuFIPuu8et2JEgCg1qSGM4yYQkAhyX9qeoOsIbpCxXIfxVM8k3My/DAjZI
2QMLLvI3VWctFLe/VNpLgu36eJgYcviCTSAZO3y9UtSyjuOycdQ6R9mcDUY8Sz0ocfkt7FPlO+6a
SNqBrThsJ1WGzPj7rzJuj231xYGlLlocsfK0dZuwScHxas+tEOQtw5LAjst/YLVHumPlknwkjcVx
dxonqCr+HXTdlChX1tJu+D1Y3hqvT2ype3TGaIQKRul90KKhTFHXBWaC9dfV8lLtrInQ50GA5shk
FPlFdzFNi0pfUaufy4IsvNavQHT65j7jkcgUCxopimMWL8XxiyoZtMmtUdYNdFRb+jdqLQD9XKVJ
8E5lMkwgZ3H8wRrUREYc94W4W0IQtr99fH1tKmSp6Ck9KaCpZdGHFAoUk6d59DV3qLKXKP+TEPSq
HTdz8L4edEmRbIsMq6cvIOEuEKJaRBrDaNDXN4tGDMxQz7FDXwRu2wqTL4FAbci1oWEQ+FNwoozD
UDEPSjbN0fq1r7MuWAUxFGoONWQCwM/eCwxX603ADGEYUMRonW1E/kQ882ufSy41HeUfGB6A89RI
c0OWk6i9t+RQDMOHOFASGHvMYvAa8bKdLx234j0RLRAhmBb4MyYqhQ04qJjuO/5H3NijAbhbbDA+
Y8aoB/gB7cLqCk4Jse5H6XvY+oDEUv/A+T9bmNZAOaS0TOnQecoGifRStevvpI2RNkQLubPCt8vi
xDca4u38zWK2EEXnXAFjFtWq2QjmZvBy209pB82lUhdTw6wtVCKqnZOTkvfdiFh+24zkfxgNf+SF
5t0DErkxI6sV5CH/1AjMixtMvsc5PQ9Fr95/qiMEgplgVHwPLjLgJBaI5tj19NreH/K8dicAG36+
mjhDdM4pPYTQ+miAzCNHj5TYD0WHHSOb3PcT9lX6tEbSuRF6tmtEuECYnp7+eDJ69iBw5JgkTyL2
3k+P4FdQlND02MX+0vJToFA8zGrR7gfcOa2hG68JpRuU1KhWQMbb9fECGG8MbrtExT6Qdrbq/seV
YBNTV1qTz9pfjq4UBLvp6DOA9VcX7/1Ckpcjo8MqNty/BAgsM7WJlhiqSej5xMxr4Qv9gXEtsw+g
fNMX4iPqWwNMwe7qBymsM7l6UB5Mdiw3gCQJ085FCDr9nmFMe72dCxzN0Buc6iCvkC9zk4/1YA+M
N0n+l1bvimRcB9CtMdjcPQeRz8xHIWnZaoadlEwE7JU6e/FEpbWnnNwh1hnLePiNjH7X2WQfMtZA
BWZs7gOC/Ms4sj4n4P7+FnKsPe77eS+GzRjQljOsvZMc8R6UMh+upE4BGq+gTbG+NaU9i/EnMRTh
R1ayZRdXYimtmCVt/DTRR2xQhgVU4ZL5SLyJKZaoRtcUXC7Vyjmtm1Bn8ui8upcDl62Y0PaJ8Xcs
PLOHQOt4cuP0VN/5ddur3yndCanPHdbMa2JnwmvbFmabkTQjDTEgGCYDCU6EAHCA0PXhFAox8OYn
CpWw53i1YY4BizIvmHwZSwntNLCnob4RcZsmgf86PLtjISBpV2zQk/UOBMBWXRlGje3Iz1ovTD3K
p4h/Aa8DUH0qMVUtu6cL7eQn1+SflLF6XE7rtjbI0RiQdeOjHSQnyx5XBjGplIrPYAcWO9+OuPZ6
QihbZIW0X5fKi8ZXujLJ6d/IRPko4sN0hpzCIyiSXO0yxSVrmtjAmpG5n6iROz7mBmfo4nVWX7cE
DVsbPs2y5boIKFa2b0ObElDa04o1wMPFCIzmOXSNI0D1KJhOnbGWx2O36fUpvcgUfrqxprz8Tkiu
SJ0jsUj9E1MfPdaRzBjcGAfOwZAlkjPEHWD3IKk9ZouljfHsXMwnHxCQqMGUx4BTIfpGO6LLVrGl
V5cq8lTxSjiYU7/PK9ZOQTD9UaiCBWqg5V8edTGSlZ1gtrk7D23fH3c0P3UtjeBGPmGPsgFP102y
MHG1slxayEeja/YXpzjRxnQ4Wu6++gghhUQmxVGtI24l2F8GLXQr0D5/rZcIL/+r2Oi2ms88AQ9J
+cm/f862tfaf2m0IyY+e9iqNVnVxQI0a1d86ydVGMtBpGU5yQi1YnDtrkokBLfbDOe0lFdX7brco
bInrVV3LCVHzTrknO2FJxlqq+gPjrylP8a//9XmJaHV9ZOMg7cIqxSqwOiAOn88iqme3xn2rht9O
v4QUavj9rK8gmoEru+gJr7ydHiuW//ghh7eLvZpAP4YDomqMp9ZIBTeSS/8oI0Ez5InNRmwkzqMA
UZl7yRzOwcUe1X99vniSEJ3zlWB4f9c7Zb3yhuMIMyuabk9KDmmTUlA3hk7p/AsBJRcFbKWti76o
p/sETVUKevcsQk+JH79gE/U6FzVXp8uQQ6TtClIV9+IYkBTCNA9Guk9kboIh+LqWZn+OCPfJtrre
Fnje6nLk7zBfjCXwvsgpx1gurNopr4To/rFUx34U4oWYRrutcTHCk+lNdvDIkyiGnrCJJx24d6mx
vO4l90p7MtwgRPN0g8fLBlrJ9aj5TytwdvNKPvKhfXKp5u1lf1lOmsT+2cawH1BBqww26MwV1KUW
uG12u90GHVFwktLKPc7W+crmvx6AA1dLWcvqaWjmR3JeMx2F7tYmjsjXSjkNzE3k6RYFB0D+5DYi
YxOvqPtsIH0ApLH5dW+J1BSJKxIIJ2n0Xl53k6eZHClLrPb9olmP3vta7R4I/wKl4C3Cec/A/czX
R5le3bZ9SgkKeqVuXRHKT2VviMIDSESogRWaMDqmacWo0fhhUYYTCximAFXexG1wKCorP685EKUO
jqVqM3jVYziZMxt3viKSqv52Bli6wdChJL5RY/RALu8XIu4FYqWqC6nMXS7VFy5xOh1aQhK//6eX
Qu79HL+SgnTxz34E97DLBhPY3JeqMJ48o82FY0Xzu5EcsS4OF2eXlf34vVKTnodxICix7vEjJppK
B2ZJ/LFGMGw+0PFQNEpsHwi2+nE+yTpGQqvjBCBo3UQByljIbiuMkOhZ09wFzb/xLPvRzf6QCf7w
fSFc3By5QUxMmsPP0VbybcSLb65AXr057UTv0tMffnzvBzvjbPbuer8pUD1XYBS4Wckm2uDZ3mDq
QVAku1kXfMi/2jETOoQEpHnTSz61o8HVGgVZBjAoSTXttkWgXcc+QE80RtceJ/qTjEne2p149nFY
Zok+MZDwtblucL4mMl8oLEtUPR0yWAW57UmDU0gXGrFQt8fahB771z0HgZDmydQ3YseFAZMNXN4d
KnzGOOQ8gh6roL5bVDsPIIH9IK0QWfoCZLs1Y6X5D7KCuz37hN8KeGuBJ3wjQEmujr1I5WXpuyXO
Xll5wGT9OPgUa8L777x047ZqqnE2or6gXJ0qr76c9htbyrelUWNsfasninb43zMfyi9F0RB1WbSC
5wJ0G4EKmjMO48wtYujWxzPcb1sm6w39RzUAeshj4CCULU3BXhq1iKRUF8sG5UHQdtfOIq3QT9fX
gVI3o1vZa2MjIGVhZGiU01WspXWgC7yI1WQ9DJxcaO7i9iKV2GqU6L13DfVIODDTeZtsFAvI+Th8
ILYJI2QZqQpR6CjVjC+ukNWAEWjPv12wOGRsW3/QgkNrx2Ud8EEFfSNacKiYinzObqdlFEefxpKz
mi2qcYETgKs8cbKb2DDF152wvukQjOWqUFG3ZkCqMscidTO53Pkn+MY5irSBNkAWHAJY8KLc5CHh
1tOGgOqDe08o0dfNscnIIrTx4EgP4UX3cODnhwdO+XCX7FNLyDFbo/lKkDMNUVdm4DtXG3VHaXve
XC5o8WO3KpgT/dVvVxw2pDSy5xE5cDxY01W5usLC91fl9KSdh3dba6FV1WpU4mRuVmVIbB7l15zL
6i8bHbLl6tYzbx9pDrf5mnvQlwkX98Afn56G90NcYqJXTBVAlObHoJ7/1eHYXsYceZ7KhVgOswFt
/L0+HMAEGDHbOI9uSASfTcHpz5x05+DQMDBb92XQr16IwKeB/4nrXj2dmZ3ohJ4SgiQWZMCFcFxm
y+CkAoBsM7lnYrgMchcZn0mh6HRnolUc6RKjI9iMqk4r604XYfcsB8L2Gd4QaCpBlEFICv6THBRj
JEaOOM/DU30ge6wjDRqc3Iel2oPM/aMdL6uN/84sF/E5a/QfM8N4be2d0TiIdeLui0Z8wxAmkGKg
VwTb5oYPONg7dT8DHEgm3n0vbTp1esoJT+Hl9OIPKNrTMEhn64efcr3IHf5htNm/nN0dKxQBUm75
t0Dsy9npB58/DtOA5GQnImeUIGNO0KTDbsdJe00mAelWtmYzJnu+3p9rs1ghZufjxDRo7bCwJKc9
sKMO2Bxu6I/Boz19TzBRmxt0rMdvZiSktC8BvvyqWlB9yOM0gKv4xboediQNzl8yJePxrjDPx+ol
IpF3z1z068IrFWJJK2G0lz6UEPQKqNtsnXg0hqQD5QAGjDHLqXn6L/8fjP15EYe9jYUG4AyQnPKS
YxDjRGZvSSSrwVIzj8+tVTQFXqDHlQTpQD2US7zCMqDiaw7lXXxOhX5GZDuvQ0s18aiLpRtFGZhe
I8E73EZ5rvqZ1DG+usp7hs+OHUpA35hafKFZUSu1uiaFPbPlkQ3Y8x17zIpiyhF0gZdXi+RlNqvG
+xwVqoXy9ZALvwMN7+SduOp97yrzsIqVkpHbEmBxU1vTy/heMVFClbAsqJBjLbbi4jwokSDy46Q7
7yUQGUK34ZeV5SCHVd3bYKrerFTkSI+THpcqAD21SJa+mNR2+y/nZqE0XOo0whK/WwU0XLX7tIhg
Cbv8g+NolbQ6LBmF64tguJHkA4CL4507juLwQdNrw76R0WC6c8i79YwU785fxUG4AkAAZt2HnsWV
csJZwuAB8P8/K/aw6i1oex3Nbx1fzP5I9xbnqyCkJb6I+ufIQiX8DNdTXbMx+XWWL00hM7br5v6C
2BAp2uo+Nwy2hC7bI2uM8K/zGxbnGkbNtGibbFlSyzV4x9EDhIaNezkepXF9zEQhhQhtVnATKfxu
3VNpxfv/PNAsayCaxJLDqY/MrKrOBHNanYxXMq4DLlNhPjfoXD8oQdozAl1ztlBm/0IjjIPHyKTm
KzNXgBcv0pPNle8QEErsWnC80IcSu4VpU2oXcOstducGTHPtzxfd2J2TAhKTEdAssg5rXV48nJu3
ty//xcgj+0o99AjGQ6rsCg325F7BB+Q6J3RYmQJ4eizflSOFbZZUI6DP5BZ1irniN4qsEG+Uj2iN
2tQeO9olC9BGzXsxIZNWIB7wiHN+iZqfzf4moRTp4hI1u6p442r+HqOMEnqmSvzdWZSSVezIWFRd
G+v/zC6sBPsERsylKhhVmxSXAHvp8yUDLMM8ywEJ5z5hHy9DgnOPnhlcxVCIVYKmwrIln58q5FoN
bmZg/9L3YdvzF+e6bhqtxK9w7AGdb9B6MUNDxdOwLmZ7HWUumF5Our4NfdEzorA8QPixfJwpSkIy
9jbvBqcLT2IaVuWr/E0Y3kqBk0t9wvBlc3li0+z77Cp3MkOMpX53g6CKAVwkkp1cWqVt+AQML+M5
08da5cW2SaYVlklzhbzW9GE+bqQsGqKaVrznyaUREgfGVkCIGH1sRqTAj3sZLNZD9bVbkcAeZMBk
kWOPaHvPDTUEX/8Qgq6Zt1b3smp0U1lhHkgJLx2O3s75oGDF2MyakFxNtrTkbd1ibh9sZX72gAKl
N7OcsfxtfLxe0Axsh9OsiwffHOdSj0zXN2M6Md/C79c786NrU4bA3MyoIS+lWPlYQQZLlFDkidv4
fy96YA/gL3zNelFbqBCOynwR8uD92ydshw/X68XBHVG10IvRalofamND1E27Hln8xiEENdqiZDtN
t9r7/Bhr9qnDZdqa+VO1FZxdAR9bul0yXVAF/JrZ8PllPP7NQT3E6e9aG88gZF0I5u6hpDBP5YfC
hUm0PFdpnLprdn+u6zAMbS6BdD8OydstefQNwpRWLwGEzKr5V6cmKXVVjSyoLQfenpJ8twUFXO77
xxP0FFT93kLOl4GiUTuViZTfFF1HW8tvFA1hRoAlXl39Vyvvt9481NUjvt3g4pDZ+2aJOgueSOpG
ttzvcaK5aJWNzyp/tMoWA69VH2w4sec0utHcOmT0FD+SrdrFPmWzeZlCiYmfSvlTJGQ3YzM5Vdi0
Fro9o3csd+HzO+ZiND31CkfAYdAfH3q2Veh3Il3bhqNSuZgkeisUnTiOOrwd70g4N3z+XLy0FniJ
6nfZokcKN4eCDFmTjM71o1S8zcRKKYfmKurSMNOVxp4sGZ4whO9ne4r1a0VQDouJXaPTN3XQRX0Y
RGIxG0uuYB+PMTT2vAcukFisiio0kAvGXBCc9la+iYkTLQBcWn2j40LDU1n1mD/X9lkWKqBknKJU
ARrY5ivb+qPNk6sIfSjTZsVhdIVePDctfKDzguMRik+QSCfNSF93B10XRA3DzwqzUU/oHAIHEVdL
NENZnk0QOwGeA6F4YPjNb0v12AzufkpsfEFJJ7iwIfgI9aHyz7XSprNrsfXWB6DAyIDp9Oy0f/yH
x582T1rVxAtNCah6J+w/AlNzEIDzgh3Cfm/tKYlwp+YD0sj3lhVh1s4ScXguw/l2qm5Qnrw4R1nB
/5jzJJsesSZvqwjxPKEPV9Qe65rgTvGfR4BsE9ws+ozo2uHW8o5HdJdjtd3OxJfO0wow5OoVDwtg
iUgyC2Dd8p3A1aFmXtgLpXVIF9TUGgmCEczWNHoPlZz4HU1vyR+o8yFZNkH1wv58mLTTrhuQFO6B
oBH/9AS84bdOvW49qZEd/uJ/N5UeJ9GWkSwM/xI39FfrCkOhSGTK48NLCCoaCXgJg5EcFPhGyKUp
QmQ2Oo11EPlEQS5ZHRxkrjq7mEmkFULYAngGzBdzrYmtEt4WG0d03oVJRFuVKER0o0xPNkV52NNG
HwkOZ2hGvg3zxuVOSltR280G1QIFQn69DTcSPNSoG6XmLr/TvHe494jYSiED6k4rtB/JQBeEItR5
wiJZDDg7gigrkjARiMnB1iXGf3NGnjBCTrHS+jsE1MG4rcJ+HWziAxZZynmCiqBsXLnqZNz0GepM
8h9MS2u7k2w2Ig35/I9JazwJtMnQVvzUYrrrmrA4eqhbJ7YbZV/OBIiKLn1FTcJBtxlztEL4my5A
M3ejVhZG8bsOBTfJf23a8jc8+8M58LcYhebsSkG+5yXje/gW3vO/OFlj72XiWe2pRrGk4UyzxZJY
mBvakrrHp9gRl7fWLLdAaW5jNwXIKBkHOI6MiUp5GtdG4DJ+lRv27Km8s0xT2++7oH5olsYtqdyi
1slOIAf7iOD0ezUaTbSgqi2AE4j6rTR6Mx2xkYxlmI4FL3zA5o+HCSL6iLhwKCv6ZgbF65oAcAoo
z/5N9qvPUbXmppv6cufMsw8VsYQrGrsin85JuwAbxKQLlfk4L/dbRkgcYwmIdBRqw6C6rH7LPrNv
hyVmAtAKniF4VdVb5wT1v/ZV0ehqeTBo8Kc83C5ZxQLt5yrUILPmDyH48sEcT460QX8K9PmBbLAu
u2AM1tSrMK3ywqaqyoE1mMMCq1OwUhtwOOXG4R/NjZNuG+4NhZDYRGtKlNR8usZnmyu8F6TI4ee1
+l5TGXt2/W9WYyH1NC2tTfzI7O319OoL83+DnkK6/IQz8AKJl6F73x7a4N6ouyuORr84CEI4e4gY
ad2znmgz9qFz3MndiLoO0E8OY1xx9RHr45y25U/SDB4z0Fu9qhLRZYS4tvZmCryAcJORPq+WfPWC
bwB7v6XrPEYr3eY/LtrduFs7yI+lJaD4hi4BFUlAY+LyIwiAvlj/LIn7D8hgvXMeswkz//ps/8XE
PYGfy4nn+8/qf9xw/vEaxldfh4xOLftj2jSKGCQpC0/7Z0zKF9D83Pl//PtT5LWDMB2Zr80iIR1p
Hy7FB6yb+3MPgZxDP5C6qS2sBKF10vf5Hg8XQcrN2ZP9MpLxvddN+FFPhBxzk5ybgE/2x6CgZMbX
paZltOVnlRhVhRj0jtRfAlJ483gfQrnOS250RH0GYLBRteWq3wcsKu/hIKod5Ww+eo1Tr2CQeShQ
LdfaDQO2/xXjU12ZGFox+XY09GVy5N+6UevaCm739MrGjgC4wyidX+u+Lx7xR0hL9KBTcdx1EpYN
ZC2n+b+rA1mwaYtnDZqCt6zjftIv9BhF58lDRhgm42UKjYyNpItJelA7hhztQPudkbH45yfBj95O
nZA5+s1qbAXi5JRFdBOxnvQh2OLgBaAjXpeqC8QO+XnulGwYlcKchAjCZ0ukEVFSZRqud3j4CXoy
VKO/Igm8iwIXE9b3LKSOwPNwKnzPnmCdbVVVtBvpf9140u7KJb+89swYYYIKAXVJ+8zHKnsjDJNC
3BTndwP744BAgLjpxSMYnX7o4ZvaCSn98Fp0kdKCJfZ7an6hdBcC1IoXdrRKvW3yA2kNXsM9+hFC
kV6BFkkza3uA9BFo4Y+KptW9jhcFqX2TrC/Tmz1YSWshi84ETG3mwTlDl3zejaGKk8q77Z71m5Hv
fgx2Gw1pbnqg4Cbm0ZakbAC5J3Cb9sc8Ug6Peu17wE4PFVuN32C40Hn648MHXdYr4hSGOguis0Ee
s4YN204WkyqWuYPopFyniAE2WnLGXOLpQb3iiRDSsoWjBascKjtqc4dLt5Qnsi8VegSJiuj/Y75r
Di3HxgJjYIzSDHQZe/gIblpEmVwLRWs+EredwO+730MpZ8q9pbBU1wvvUcllMvY/lJpJiIEMA1q2
5otkMS+JVFKC22gUoJ5eS26a6fdKlh1aJHyM0ZjUA15DJut9Y7+KobhHE0imqNQZKXNEDq5ZjSdq
+aOPGoyunU4UsoCZFBIEteVQCnrWaeMGONKTUlo/rffuDgohzYeLTJ7mwPwkr+/gYLhr3HaILCil
uBEpyf7Lc3Z6FJYQEc7a+Oy00/fvP0Yi5EW3wDiKHyrUXiSzexzpO0GD5MeTzYIUEBXAWEIT3cEP
Ic5VWxafZZys0TR4DXqb+sLG9LgBhFitx4CsjJ1VAuDS9Qj7zPKa9zzKHAf8HaK6W81Hi2Bacfqd
hAhew/7VOlm9arbJE3cudfgViriJaz+UzCVvFpQroICSbd6Fdll/yWJDgpKvhuFVJPPw5o3A2QY7
zw7iU3bh+4nl0DBsVrRm1dfdjcRKewCwRI/YoBrl1dtLG1br+K/QDTnKwp3zfCW4CuEIaENBOiIZ
evtPXw+wfcyWMga2RCBM5SEtnPVcnANz2Vj3ss85ruiR5Gy+C07dw8Mm/JMqKUM4MYNrJru0IHuU
U/vKDVRx8ZBHWVM7yNn9595w0eW9EtG0AHz5j+z7DZRI16e/6bI9tTBWhsclal8/8qj+JN4C5E4w
QGRR9HgFOb2V4b7OhCoR3EGl26UvxkIKxVf/Tjjd/plFNcF0woO5/CnkZQtIy4qN6pCL3NNIjxSz
Z7mLdreBSebNJC0c3BwTyzBNi6EIh3txlPyDto13nnS5owzVbsOTfhQhG4IY1i236qdRK3fAQa65
4nh75WmotB6uVwFEO8195xqiNX9m+LdUDsVhTmUF3kK1sQIo+vWqFYPeqDwwa5HuHSpGGQwxxBJS
rFjEqE2u24TPwC1vZI8jUBTOfXX6bJ/I1nsS6e6UKTmuDqvDv8B00sX2aDJZeAiK0rts/0acqyrh
0/KeLoF73zVIf9Vff2c722zll5821SRtt/ZaiWqyzCFovcU466TNz4XMlr8hvltNpf5se2W8y50h
dQiGY4xj34IeHcdK4wYN2ffaGAAsLZFG6LhzbJSKRykUOyRNtXbhcBqzzwlcbUi/BXF2c6v8lq/Z
1/ZCuzGb7Cfh6GKhc7U994lIcJXtvhS4l1wJ20zqP9E8FhuSz+hHR2wdXz0gT1HWDbmnCr/0NKGg
6iKQ9rLg2339Hns4E7rvjuAUSbfAOy3BmnXt6y/VZh1ddPTOXljTRNO6CMLJbo3AB9OIfzVa7Ypx
oC7lGlUvWCxBaNr5t95zkJlv7ImA9XVGqw6BUvHJq8xfawy/+wf2d9AFBzFrGM87fDy3oc72LXOi
nQW4b63zRA4za+qxh0eS+I/MzdsWVPs9QnGdWvmsMiVftgLpdKTgO/PADZ1KewGrvho+tXGeY2ah
F6ZBIW8g5Z+S05N4hO5H7wrmV4cYXSEzAgp10lusF9CzHkaMHW5vd03db9mkJDva0frEAu6x2ky9
yFkjBa5u71l3oPWt4pI7dqcIqFlG0aTjP7FB1OXrthmIF+bU6Uz7gSj2oeEOtfISzgdXJkdp6Yi+
ncpipckgncYNPe+z8KXbwGXzZp2VX5wte3VYqMSiCbpkkv/D6xW24HSCb7vBALlHWW71tJL+sfBO
vuQ2V48rfCv/+k19xDOsnqYgXVhSiqf5agThDFIgWBEqeb329kCRbEepMDiUeE4rjGk8OATfgnXk
SaFes0lPJI7qCgBH9BUir5+unNCkz0JG5mqCu0ISDJ8HcNiuZCZ7S/iW1Qg0u9H1xH9qbb2HZAHs
Y0xTO3uUnyHz4XjZx9dzwf5Zz9mxb4eCZl5k8mgyBXsPimyqkkKzmq7XBRYL+kXUFUsxsSX8NN/B
VmB7yY98vmBJd7dPPw2DDbv9TqvAwk2UsZkJZoveFSrXLkgyEuU0m36fJWcjyF4azzSkBlcmzpTK
/KDxKteE3qbn6X5ReUhGCLUVNMw9wlEMhT9yoaLlxGUcG6m43RH9CVrWW4pIyhsBUed91G8fSEuR
VM2AqOFrIg5+4EOxwz18jE6c3ajFwozspwLOJVIy3Qwn4tGDNIih4kppNtdlhmcMbwLOpaVRpQe/
u3Z6FYkWKnj05G/6q+B3Ba1V4pYeF/SSiQtoA0KYTsZZm2Ly/DQMGCWTTEjyn3SYm7OisXvqDavr
smdXsR+CPmdoicV8DajwU8Gcl7L1e/jzDmMSyIAZO8mR2kAIgJ3RLcoQs5pMqQpw4LUPaT8OsHsg
mKx2n4tccdS1f+O3kmTkJpej3pXNxgAgDbY68Nry/aOMG9JAQUpvEw4K59PFlW3WXHGUAIt/eju/
pzQMvWE3cHxsoWxdHeuvJP5yQQhufmQ5v5JlNDqmpdgHMLI9Y1ZA3vZJMSOSGVjGGj3DovuZ1gKb
wH5CbDlco92qEFmxtW7fOzbbSsV3p1m+vABfd5isl39obSrQy3yKfM1QD+uKrPaURuCgaG94AI33
Hb9t2AOzlF2lrdAiM4qyuUslRCsgbAyekoCvxZ/sJ+DJ9J4BqTgt8URBTuwtISctiNWlnNuSwWab
+5v/WRK6nEoi3L6HL1hB14CI/e5DuFGba43kmvLXfKOQHk1XQ6JU3NWrVrDr6+m5LkYZ5SkmyI3a
tt4oxAME0w3FDgk9Ym9cXO5fJzv2xEjSZupWUNBUWg9UHPveeQKRmfCISDcTwX4S5L6uQejxC2yo
qLiJItvvxuyUaS3l2pjNhXcJ0blwfIBLPVxOYf+FtMUXDjs7WRL0x9i0Oldzt4dW7+p9jS+VBq4u
MiG/5E7P6FH8TvbqcnIM4EX1cl7JhSoXC+iZ9WrValmbgJaCXT0bLE3jtVUpZrRA7wBKSFhRepvO
qVofwR1cQ0QofDJxcM91+9bLh1ZznEa5h8hhzPGT0Op0/z/NAr226h380wKGWylMx2Bo5hZHaEJn
4LJp1rzGoDbX6yd45EUDpx8IpMX31oa0MVxW2dRclBUcx/56Xlm/qLUmUBy0UkFJPEJ1poAqziNh
vY5orb4kZt4vSL9F2Gvyj/pVoSS+PIA0s6BlJ+3HHbp4hrRGOca93bnIVOejotRFgO+cCUB4G2Jq
Lh83v8IIZLYuT7UtAnI0YlEmABjazi1MYdEOlJoMN0iX3EH+bj6SjO+tLyouQ0l4u/SGB+aqyJHF
T076hsRNcEbFg50P7PGmVoqtqfk+xcvitSI8HpFJifQIJezBxnb3lWBrDgloDMCUzc9RZHlicifn
lTKfiNLQKvf7ykiUYDimeEMBE+7QNyPy1Snmt86KSYFSXKhe7pnz9qT58afefgFttqYUPyo6Esw9
7xtlYurFXg1T1hA6PFDs08iszzq9OTtu1mzPOsQPdOjiT+Kf5QeVP61iS+flL97bUg67srvq6+ay
db+fpgxGSfxzPcEejCmHrvy6mcaIf0zFa/JllMRVgE2L6oIE63Y8/Nds/VRE9ROvRpFJdfxor0p+
C9aUq/1JbvcRd//REMWJUjttbqlhe5qdYyCq8DjBWSsYOwfWCuh4nZcCJYyzVa0Ooc3UoQRQ/dz4
uId9v+0KzH+U0whot1nn/D7KwPKJ8cpu3Q3iga6FndTCTBsTfGiFu8J9SJiVRSsM8P/hZhKz8rwp
gfhnX8awYdSCOwkEV0nQgOEX6UHt44HaOznWz+kgX3OX9aP1Yqb6GD4uIfIQEqsT7bSDd/VwDWYM
bJIPKV58HDFhTHleKx1qCxNJHAGsARJwLZ4R3zH+12bCua1hZGqt8lt497co96RSpYJiBVTiF44+
MeeAiM3+XdN/0OoZnMOdrCMqi8Dc+2s1anNuWY+f0w/4Y841lX9iiqMCvoUChG/ta1flmS09P87L
jQ7zUpW1rQMN3SBnat1QCNzADPmB4vH7ucDFNPKtnGj4kO3i5biigqO9o30yy9vV7p0hnhOlTo0R
zCKyBPebmLAxjIklsPK4NiJPWrjOuMiU8bb/AwR37tX5B8dfDZSO6y8kcBRmY0FzVebP94hBjtvx
iVGu579GnQU4glBwui8TsVr2Ipfh/L4rmIvd8/bUXVNhXHl9QvLcCEHRvfrImTDMXr+ngIeMa0os
YN6vDdSwkCLlFZBepUahEJBE2+MjJ0zvGmayA/1Ao8RErX6tBai7YtJ3xrBRx2VR7avcw8K3d6+y
jCG46lhC5GnmnvAsUVIgnoCL9l3cLGDt2V1C3/3tnLocMILiKL+tyzc5PqtO1KGo39PVZTZUws/n
aLl29OQTe8F9RW9nnEwILA2urKF/RZpFtcWTI/NUUfrdyg8KzEMQdE2m0zNEPRGQXAfFaymEwhjU
Lh3ql6fFMSYP4xi5LymG28w/Ub36EuU1No8093X55kFoOuhgJgTbi3eW268p1w7e/kIvUGE2+l97
LoX1AaPCPLwFSCmSKxpYZCEGKdQvzQgekwD3KDv9nd2zGHucs6OFmE0eMRKyDgLC0k4QM+cr+SXw
HTf8hjVmKiKRo5WDfM00NJGkC4+6DB8M0aPP1YVUuMGZL/uInxUAJSNk2sUYDx1Tnly5MwNBgjl9
/CmVSE/lW1+eCnsVnlpsobZsvaoWs0qAnrotz4m9e9zIUkmMekGeuZuDTc/LH9Gkb3dcpI4R6cp1
2BOu00q+K3GHQpsUyisxLAniGzJsZcVatOGeGDTVe6OxIbXxox1iAznRbTwDhdfZayg2X97xoCBm
quy+Fd+WsMQLhVsQcQgqGl3XxARL0W6MVIs368N22YP7cZcgWmOjTmTwXLrauIn29fMPw/WcWV2W
/dRuEuZEgxOy3uk8wE4aERhsbnaGmalBmflh8qy+f9Fv6up1+DU0FJ5OkZ0YOfBaLw9+5MX0OKRo
0xgooPlKfVVf0Wd2iti0XxRE4xiZLRLrkDu1VlslZVMeCEtagAKJchMCN/mjRk04glfn4XMokZtv
YEa2jETtZ3nM3f/E0sdMX/ldBY4/SrwYb5dZdVBnw6kNZW0+3HlEUkCYj2ZJk8aZvR8BckVBfFnz
f1XkzSVazOB6WHbOeRM4dA/k26KqVnTUkBcFTAQ+Y9aLY4LUhxBOiAPxvC87OBtD5ZJsNB0vc5w+
siyIZ1T3XGek6z9fIOu+W8mLgJEXjLNEGIrd9U415GLeyb8IBxlsyxPCBWIhATkJp0ong2bP59d7
YA3Jqh/WfwRsZ1GkTdE1JYSjU70KruG3uPA8WzNpkPNfN9nqtbS2uqpZmn1H5subSevrpAX/397L
rsAhLtmhjQY3YiZ0TZtumflisdatJ28SRRahw8k9d6QeFHTnKOiOntkf2QElLTXatelnXn2MHYwR
HTseRgY0zr7ShanEbF4b9BlID6a/K7rDdxpwyfH3ZqhuF3uY9sS39N2bDZb2pE11i1QORmw0NwA3
NZfWxYOtE5yEnDMBwlTmble3N+5KKvBKiVQ3bPQGMmNWpBRTEbFxeRydqqF75FIOR4vb0yEQugLN
KPbbC1KCHsKHOLgwPJoS4JrRLc5AlPFCNZdcaZFbYA4bmNEGJVws33YHzeaO2DwFrLKzQDBap+a/
Zpe5zqKS9fK6ngUS+NwfSZ7NplV9umCoRHEln2OZieuXcZlbQIf+6m56MJkDW/3zm6obrvSAr1Uq
s/58TQRpA1T0C0VjD7RocL3TCDA+lqnXvsTmScRdEouELmbYpucgJmLECqOzCExmNd7AVBzz1wyN
a+LvoPVwQ/0z1567MKu4r16XcMyKg5sGxSBH6i5nlRiIwONpkdZ3o9257l9Hr3hkw756rFjvkBcr
rx93uU6KL7iC4wPLD4k3p+53xbj85FbG8gT07aRyN/agOudzBZ603H3Uw5BdGFfwyhw5oZclFIH8
qxcJerNfJLbb1vxhNG0cTY2eoPvLe/doR9HM/sG1txZQTer/b4Q+lrPReNKazcG5QAzLcgyBCy8j
7shaPXyGwjPzgMUvcbep1VAWZ4gymJ3Rt8+Lt8SPdxAU0PmjUCxYbIGG73CeP8fL00Q191fxgZ58
WHtXbRcDhUM+9mJLp8yg33q+k3jEcprMHC7g8PvKIOfxADMvnMU7SilcZs6iCfW129d8wEJa2Z8Q
7dLvD+aEYK7GyAAzpvdavrQ1cjXOpN9Bna/POEnHLIouiq7V0Bvtoy1PFKbRwMOpIAmK0/58+/2k
yxMwBRYNn8GZnTBxN/Y2jxewQeYh0nqODWm8ZGwczLHgGYS2iwZh09T0evfFsMnXuDEUmCb11/Nq
2soAx7B85lX+remtRhKSdQhM9DX9QpUO6HeqNqddMR4KN2E45ygsuu69Hdb44WEmuzd+uzUzYAh4
o0W8zJfK7pdovB2wdhzwq2E+vvPYxXRNRt8phWAqboxuLUaDryElr/IxNL+6Zvg2IDjsCsxQIJyu
CyUAqywO7dOPCTePyI2m7Z7QQxsEyPP2MX9rtxgSTVHcXBoKChY5KmgKWfW39QYplL4OTq5KnYKV
3l7gSbQYzY2gOSwHBYIyatty3RI5ujrNqKBJ0c/CHQ1gGXPTkhmTyMgr4Bwfk5irfxgxeJ+f3zKY
D0ewiz0XbCHpPv0e8rR/siTy0LX+f7J8W3PjmE+4yPe6BNEmmxP5lNCVgjAQDfkrPctT2jcYZjPm
v0FH9hVnSaAf2t4gh9ftRieDC9r/6VEY6bH15etuNjC36+Nf4sFxqXNL3FWa9Y0tmvlHnCDQMGfI
274xImjLSV+hRe2mfWkidNs7dLRUI2ineK1XY69RFIP8Hs3MfRBnHKSV8ikEQNeuErnQSOcwBsT5
bkKJHCXBZGTHC81jP4L+QIw1OqphitptQJijps8nyzTfdCx31fsClcZw5L3WVqZGxsSOHOxFNSPX
7ajH3EV3OBFapWdJVoQWrnoW2bULVKNx9gabKcYaaYUyH7/pc7znW5qhhM2SIX/ZxPzdK75a97Rd
VE9ZE57bbadCzkmOEvHfJIkSdZg2lXoAxoLFxDQWYUkc1ntooeif3htVMENO+3KcqQ6mfALIAWTe
M5HY3rsVcqd4sFP79fy4BPRZsDsVqyxTPNkVw6j5DrBDfaoaM1IEJQ31sTipBJeIwsQ8/kWmMqmZ
LwNGpH55l92v8b4I2cjXxuubrtI+EOxRaLVbJuwpSnBL9JR7h7BOMENpsZk5wGJNXIXxXk/dbgUb
zBZHDyrInvZlsSgFC29JGcDqichgDjARM0IHBukYILlnFfDk44AXysjU/mhiSRl51cBE5Hl5gE4G
iqFNeEYsTVyKoHwg2g0ZNhqgDpqI/CEJSkhNIkGla+MhGOOsHuiynU+zbUeox3Fm23Lws3ovRzgB
BNLTB5cNG/GihHpqW8GJJ+gSy0GAE8WpVNaMmfnWWER+nSEBwkWhOHKZHg9TV6+AmuQS9xQHlGgQ
G704E0Q6XYv88EbnYUKrHSXMwQjSswWV/uxAaVNY99GaNkF+08Miadl4C8Y5cuSWTVduNbCRbOIC
nObM/fMA3ElXvASQrEgbHrKp26ks1xFF+ZD/roKLtEIMkh8HlLosfjs6tGdoXob2Omdtpq6wJ6TJ
8ZBl+jOK2Ya3MLkJ1NBxOLgsXCjFqOaVRDH7ATmfEG4r3uHuPcuAFOWhaQ1wPWJ6nxvzjtXZUwE7
DX/enyQTIiGJH/V1gksdlLrRIg5SiUf+Kp+QIS5pf09XmHeMVgcI2R0ExRvAeXpnpOFDLlU9H9s0
MEWRfHX0/sTWVj8luyldzEfQUKPVM7+DUfhmMBwvatXNloxmYg9XtiIJ7Lmqk6AmGBlmDbFt0rI1
PyVGNqVGQFM9Dakjg1Z8sLn5Xlq0Dy427QMxLY4fxfuckpHUZzzetOUOiko7bXWZZXwJ7g28cbgW
w4ajduqB0xmSDmhZUygBTLaIzm8htyWhf74qXlat4jK2GrwisVl3JhU2jhwf5ONowLsBEZhBatEK
evQ7hXN49lFYho96awBGeFBI/N0aRPOnXMrWfJqf0WcyuXgTMhKI/uWzwG6N6i0bFqlQW6r1/ouT
tf23kKpUsZoeon4im5+yuL41cWgdRGHd4tblJfO5yCgfRrcwycKnawiKNLowx2tVcggVQtl7femW
uuouLgt1E0e837hDx9CL2PIIDd+4OAPpLdN08NC8kS4DuLZm2Ml3RYPv4kLgD2sxgvlLQIX3YDJ8
EGYxw+VnG7aponsIkzYb//ZoeikYy75ObQJx9lkIpgodcjhRRQz1BxUkLEfi+2Ajru/4dSy6rR0f
bOIYUvMqvzbPMdKVpT8YBOXzcAvGtqg6DRYVjBFYt0CT/fy+iVGxzsVo++zweXxlJua633s6CBGd
O61kHBc9s7rxbIkLa6OCFkOhopbZ8guTGTPjrA1Hs24kKRpAIrIVM6lsDxRDPfwF1CrctBfBe4Mr
gLJJU6IrUdLeFR0Sgku2yNnfRnH3NSihdejOUZD+R1NFBBuhOzga3KWXbZuP4eMaPOBzjKURSyte
exl5+HlgTUXvZMyHxA034Np6HPJTmAMF1e6xXgirWFqJMOFe8YgnDJjY1Ei/dkosu9N9WpC/0c39
QOgu+JVRFaKDLDBBNm+9XmfVo8I5Q5OTdc+j5mjTnK1cWzh6vFSetbZ9A871uV9ESMNcM9m6kp/I
E7CExx6jsHtHMY9vqF5VISDyc1NfoLfG90sbC2PW7zPR9qk5DucXVUVY945l1OEJRByHtKj0Put2
sz4LpV+ZOWiOXGD0hTTYHYnqq3oR5a+JEMta/utmPf25oohCdeaYeSTMf3/wmnDnnNi4cx3IGn4V
BGkVDnU3smxMq3GC0qaGJ43W5lU3WkpLpA9l9GjozAHaT3L9gtgJ0wI8TC7O25z8+0MGyjHsyFc8
tsqprUQzUB6P4Wc0ivGqgQAm9tVTqadAlC3o//zDTBSFtxkaq/1Fkep3qagjM0r7BooCj2I+tRmW
z7FD423MSmWL7Fsoh5f63QbUE+zsEaXpnimNNX6x0ojy1ZjIXq54bYN+Bg/U/Rw8f2X6rEdaUcYj
wezbtCtNoRuvE6MUCTZxA8v/xkrV9ws+JXE3J7cLUbNjue/Rk4mS4tR1Y8vS+n+WeqEhkIJbKscE
Gw7qvlYIjjpLYIzvEUdX4KsRi8Hi9Alax3yMxYyBAw/SqClfQNZRS/VoZD11cYjhYqXrGk3FsMgE
WSOahQYFXeV0Vu9RfqGnPbP8sEVxfkpRNM3KZv46g7RBlJWGyTjrt1gXFZz2FG193GSzqq379L8P
MdvClR5eMz1ABBiFcqjJ7ujHEKnNR+hnSMcD0UWGwU/h7rDAGcfr9S6o+/LrD5sud5e1HOXqKNl9
8bQTTi2TL7RtZd/CA3nhN86MEEpxiG06B+AnPIfkUct+5CIvZeOo6jsg89ERNgn5v2TFG04dKxLb
PmeynUMWYAi8K+ApQRxPBwB24F+DaH8GNsT6M60WwQbDfpImMDBZkvNgeR0REOem1EMd++xKvKz8
wKNOmNphVHHArdQOn0DCX+nJsFKeO4SDP1hmM5ZW4ZrppaAIHg0u3sGHb9lWpgvJdGlyMA7jJoHP
gLlucgbOYB06dRxieSmHayrv2TQ38wc73I5TFM8Pk0Jow12EoYiu6gPFsd2rLv7PzUQcbyZ5xB3d
OnCjxIeY/BOuV6TdgquQBVJnjQZBVgYz+DZn6a41I7DMZ4Bj2r1WrY6oAPCITNYbezSyia+egImy
QqrHnZ6zp8Nhg+QWikaDGaMhIIBbYBMfEfNrg1l1gca4V2NqByZg9eyBjzzvyBacLvaceQOHpUPE
0cczHOGXfp1WEcEoRioD5py4PXPMI5y4P1WcTzpNO5ul7YZrmYHFzSbU2uQjtJyNuMz02riUQhT3
ip3rQct8Uvg52CVNY1z2Gf/UEbvwBX2uRXSJNty6WK7p/HzDENW2ZsStmX4VpnubKgFc3FJiS7pi
fP2MRNzXc8vyIQuT6VXhktBTMBa1fUsRc8TxJxp4ZMuICoR2jzEwOn91Ay6xQEm5Iruv1TQ3t2cJ
JiVVBsBO9cKmgXXHdo1F5LGw2ST6seN+DBJWjyGtkQYza1PP9SSxfHfXRMorVNTLZb7TFcyCIcYJ
IhhHhGaqXAkEVN8no2d0QGVPLmy+4sx+KB6uLQVWLhSq/uJkB5kAN9GuKFGo/xt8FAMyRWom7UXt
Wf7/OKBK/wfWTorJttSuAydOvelsuKCTzZcXI1/cF83IJG5e8XeYS4NGFNjJO+TKy0A2XpX43o7m
VM0dp6NPZWkCuULDi1vSq0rh0BARm1yxCCyhJSsg1emZHw232+rkmNVL97SnrjrxJaqpJcE6B+4O
7Chq50yBvBmD7tlzi1lBq576NNZX7VG/jwKWp/XSpd5smOXiPZONHKuoH9zYnqLrcA8L6aLSiyCi
emtPEymOz5YZRrL0yycQjkUzxZUdYYn+2YTFMLllFKA9c85xa43ruqCpXBATgE/OmoaPAXabiBCA
2+pe6kEcgNz9r3sBBNM0wUASVjzA0e7m9r9RJFp5CvLcPN3kHELvEPnrHe2Iq0BX4wB0woVJcQyw
Cnp4yp6+G6bRUyk9dsVsxUrEQFRP/bEvgeWAwc1oqLPimQcb6JxWhJFLKZjGc7AL55fPmA0ZYMnn
UW1O/RWuAIg3Zn1piB5qEeHdGde7DdUe0E4AsEYTxJZpfyBpXSD9SalgoLbzVZAuKDCPwyxFdBdO
vMLjyNsPPqp1PQtCHxbxu7aW0wzSN5SERjF2rsBw5R2aS9MAjJKjqsju/yoLOaWHfZZhk7RUdGPc
Ce962WT5U6uAGRR8XA9AjgvWQu9jn3uhmeCnCM6k0OYV0e38hzvRe6xTE5BsYzFyzoXbuDIfbH/g
xKObuOJ9cD3H2XDwEnQ63/6qjCF7ZCuqLSuHnRyvn1RDr6djeG8apk7HMZRt9GgMpCWVqIzlE+gl
FYonaifHZa9VVPwmNaeZwEC/FkGBbNM58iR6fMFJc3/IfrIxXVHRlQq+RyWCgPj5kPuQk/yw7sNm
CiYLUvOodD4hQiBGEjQ26RdlkVsRYZw4GE508nJ/PULeUYaelHY0C//UR8qRDy5tU7iXf8ao/1bT
DFGgC31Zg/2W8uF9wD9FEw8guwsInvNq66iT8USbk7mRVNhM17j7WEY9rPCI+wZkJFVI2SLPXOsJ
eO+33DBaUpNlNXNRcI4wJ5Qxh+yIaA8bSER+n2Vz1CvrlfThBnneud9unzGKL4mBqM9b1bG6Xrs0
E90vGAgvoksRGKn6nDykRQ2VrBVb8yVyni6Jh5GefgL9c+S2vdEoxL2HHfSwp0cZe3I2e3Qzjx9i
PMYvxWD2Lo7KECvmenDqqunFAq4QcPGRRFUM417cpLZvWMimqWLQH+/gCheDn3cvmeeyijjV/XNT
cQx4l8cX7G24QWyhDSAr4UlP3KnB7I1o0v5psPpDZ0XmvWQ/Wg+JyC0W1VpGINV+o+A8/Iab2G7H
z+YzI9LeYfsCTX4zqj8P01I5HHWaJ4DEpwxfq01RS2Ki+fFEONi3LzG9Cg5bLPfMUrF67MiO1XR/
N+45ak0UWV5M1p2HeWzMPyNI9nRAbV9FLR2BO2kOmbpMU7WNl92FV8nP5R0yfwRco0lh15jNVvUX
StUcbecfd6eJ97ELZjJWDXiukmo1KwVv7GU8UjsRrvi2mPEcaQtgRENPeqRZOg2t85XB1P00/6Tn
fMzyy7Wg4E1EbWtR+6MGYpL6gVyIe249KxBIywyQmUiWIxmPEYJGmrXdVl7lLra70FPIwcpczhAu
lBLZRhgmFyWuIAjjIfhvXZbQcEO9zxFqOnpcpvEwvA+eaPZ0GfVro7Ztr+SgI/vA65EqgcBLCQiA
SEYUySpLDE+uELhOgzvxRCJn/Ufykk53ji01s4DGGm8yo3Z1I+Mheral3PPhyUKmyN5QTUp9JEK0
IWu8Xr60ja4tPr582tmHiw1fbeuXx1vSKxsZopm1ULDJ4sEeYT4vrbowJ34lQjQnRjgaIYr8fTRA
oF46DeZc4Fa/HYBCf/Lw5qMws0uvxz6wt5o8uqjgmOP57sJmt7zk50IzJVhYbtnyyv98LU1i9ziO
aq/STm7hmnYAKRYX0Q3vJgb2Ax+ySM7mMgksYkt6b/la95eTs1qSZVsZ2h/oSbmvFVDMShAVDdIe
B/c1Clrec38uSAf7PFx739FqasEprEbb3at2tc25gKpP+PIkaTlc95/bUUPEb2I6wdOx8iG/hKQM
xMb5MbLznspde8B/SfmBqlaYswyjDKEICvkqYexMDEAEolQVKa3cjZedLhUCwULhJkYTGRjrqv4H
1NyG+iCzQdgnKykLom7X8VnvLA4Z3TVmr5/2lOFrPc151JJURzGymV4rG8hbLV+iX62uHPmjJloL
NwP8730eIU06rb+0Dch2QC8MW6TFkexZ8VmiKnSLKMIgMwEVCIP+Xl+Gx85qKxa2Gr8quoTFep8x
0WXFq2HRE9HbrTFnpr9LKEiJmdoHWGlN67w+fkjrVIWWy7rl2OeIk59m/pPhX7VkditZ67I5BN9n
M6p+xnYze6gLR6xXDrf3vBqebmHXErJrIgX5MHKVRCKc6MDJlGYjae1Pp0nrGtXWe2m6Sdjyz/um
xKVL4b+Kyc81M2GbVmMRE22Ca2+D4PqYiOE0cpB8hTqZB6JdXOgsKWSjyHuFnPLNRKEzxxOqgfDP
k72Z089tbUa6EAujXHoMRtb5acT/EInKLeoBrgPBJNiRmvsV3s0o4JTQAmElnLTl8aUfDZIWHcXs
lWRWOyGvqJDXFBPiLLK3RRqUEWif6W4UpxCaOygVq9rM+VFWjd3U+eOmCTLAIHMbgf4jzMH3sS9U
mX8fBbnofGhmGDJcjHNq7+BIfGAyPvZNhFpaNge2EjhtFfCq6Lh7UD1thgnuTOuzUPYXwkb52kPG
v0N0SNAh+hcDI5aueu+yJOHUQtdhbY2S+Qso7n6pYYhb4ejYBZbQPt1IbJW9o4JoDtoJ8g/WPoeI
4c6JRe3oqBy7Ay+23t5LoZ8BPT2TaavKT8/VTh1m+dA9RAYgO4TmlnNBnlyrm+f/zYxl//K3XdyL
khAWx2aSUphvAN2qF7Ukmv4kJoe/S68XqFRm3pE/ZT+F2wV9ZqIgjws1FMXcsa6BoT9Mt/LcDgIP
fv7jYqXexsGlCqk3yXTYT3xlqLeJM1y2RjAPvb8e2JUL1qLWOtGAFsOUFGfCZQqbRRBuixA98zPH
PaMqK3aBAM48IE67Y1Pv2xYgc3eKLG0aVX1CXilLlLVaV0L0erCAIkoYwJRyNeAV8IEXhRysqjZy
a+ydmWGYmiWJtycOlEwHd3TgSCaJNcmGAgmKjazA6aII5YXKdLkayuGKehtiEh5YH50Ew7rGMfXb
JdwN2c2bPqHgfHVhnXCvS51eqeTttGJY0sSww9ziWakyw/uhZUCWm9u5KrM7krYqtn/urtUpNmoA
jl+mT3DECz2REgay1/BRhfwgiiBGmBhfioVsTk14AQtENYdcBKA+fx6bV6RGGtggVXjFMJY4Xx7L
EDSJEMcxZ8qCnlYC2qFn3vJG9gvlFKAeWshaMVJeIImuwqJJmo5TqMR5tGz6XgfI9Dvz51iQc5wf
JPWLr0zCWqIjK2JZ1SgxG3j0PgcLw9XYMVilbrMWqg6odZxrI33DCIpjWRPp8FuMfPcrARfZkfb6
ia6j5SUrffBcj6/BOoMKn8hVjJ+xVgIbpulYD1iHI7OvWLWnGfZ3tS5I4nmpAeVB3iEBfNm9AOpc
kc59QPHUpmh9rcH0UUbx7oLvVGyLhgb876bHY+QDbPz8WoOqDlF3rMGE4lwl23Cczy7b3Ez7Zhx9
G4lv9Amgw6osxuXMr+s8+UA6IKSLecNvyodzDP2A3a4+utTc23xwBXLCJJu0E6kkzPKFEg4aJU1w
X4Nvb13gfryTP2ZMnib/nbA56b4xR4eHj9zJe93fqgDC+FDdOF5yNs00Hq8krCjAsWq69ej8bFMv
EurIrtHiH9BqzAwRMpTRL7jGsWs384jZmuTNRT2S/670RW0yZIQWbySZhaqUTwTae5xa/3MPPZQ1
jIZVrcLYwxXxhIt5w0PyGhTeQLeVKWzTEf2Ta2d5lcWTCdRV2EUoxOG/Oo87wxGM0xQ5sngMjuPu
Qx8zPUNKHsUlyH8bD30YMqwljb0/gPpcQDDhBcO0XJqXM4TYU0vF/KeNbcPfL0QGweNEM3r8gwz9
lLKqY6gcBrJ8ER/pl4mxFLj3rb+Ac/f1/5B+xoJQptNq1CqjC1Ik8110j0DlDtTJpRSWKIZe5gzY
a0ZqZyO8jswxUeEEz4ZafWyc1w617UHZR32Wef5YRYvrvYqzEdIp0pQWjmLMbDlL0IuFaUwX2fhs
cNT7qpn1KD4UL6zZvzxALOzJE9nccWV2z7Zdn7HXwa8FRuFT2WYNemgoddQ5Z9h6Kd9yHk6Y+5bw
2Rnf+yjf3T1xp//jRlKn5il6rFC7hVfDrrMDoGbfAFpR3UhshpHMZ56AOnCeN8FbrLoBAdW6dm+N
qvg26pJ5loEZvpUPg32TP2iVDQdL8LA9oB699thObBT10Qn7w7JluewXoLaiIb4KD9jcm7we9JZD
p9+NP4lkPDxiN5MHeqKi1ucHcyKDAi3qvI2a0wEzUa3zU8T2V4gbJGUKFT/z2ZKRguJGKmCfGpG6
G2H1aD8KT73GIHO1hBYqAVcTqxG8lty3r8zaQTrWoJg2BPAH7GpfMo5AYiwNd0fVycGBJJeIiwF3
U9iiZT9WBPR7DNT9qsJyDungbBDHRfvqAIyb4c81JjCnca8YehtYxxmsS0+Jx58QweX6G5gFq/2A
yX9eaUYBZ8Oxwuq+Pj211xKhROdBHPSlYqaKOkscSYJHOFUxQ4p6aie9WV51chRbGn0msYc4ORwk
NPPz5Ako5eKiMqe8XxVD/WGwU0pb5NGYEFLsHz78AAJZ2I+UqifY2BZTb2LRgpy2SPovS76hwvbG
ToDaV/VuvuNfwkTuBVbA8XukZrYyTpBPFgeTlNMdSUK/rY8013KrYOQcv/yxICcoHqNMGIdvP4yT
zuQ03M4HcvC2wacj6RtDsoZLnrB08y9nPHEuc4zZ/4aiko2iWyJu29G4Fma403Rafkl9ko31Eo51
OgyiAZkxpsYKQs2rAl6EWa3kEzaCA8UOf+Z4Sbeqdyc/3PIhHz8ahon7U3sDMW+LuJo5H06vqL8k
oTJ2GZA0q2i5Xg4IxGpHt+/NdWNHx9gibVli8j82ayWgVRBQMfSiSXWFoOOw3wZ37h36tOoh98BJ
5YdxpKnZojtBe+l0NFESNSdc18CzBxoyA/kEsLZGmDke66SpbCxpyXgzNPp+aGL5Z9lbk1vkKzDn
XkdOv2z1PElknbXa/ItC3HAOVYHhZptffjzHKCi337pXN9776FQGtCcCjR20l1BwfpbP3UN8f4p0
1R1tj3GlphdteFc5yVoPm4cpYMYWR87immMEwTcvFRlHA/NO000kwIj9aXtLgnJjPUjsUnBx98ys
3v2stoHfkxAqvDFVtipeTgF3COaI/lC91SajkJGEhBPbsBh0A8JEC63JxxRy/9O6LtwcVmMci1EX
huQ3+8UryVad1uSXnFy2qrQ0soZRVI8WPieidnDT6pPn4ofCrLF9SSqhySG1rYNjRujxu/ZlcXZ4
00SbiFn0qvhouj8Ka8FOxgIEa44K9qHZssRSxpPxjf+MEtJF9l8dev4E63xpx3d+JjrTz9UnZM49
GUdwrSFwfyh/nitYRpNnv/KFZlcaligurSoCOrOFxd2HRh0y0/LTf6d98JS0wbMBR798iovFjrpo
1TVP6XtuM937HrCpD1XIsPhcChWkLYO39dh0x2rfiZ6nsPzq7bC26tWpMFYCy7HlX/7RPqVh4BHE
rfHxJCT3/nLRP2vEWEj6Su/hxzCD6RJLt6JgM3GFZNlluMhwmCZH90j5POV4tckfxmpzB3syhgVr
PQKGZsrkZe33DIkn/42OFeqGvgnW2WItWAVkoqUbxSaCsNHX9/Hw7AEH8pMshLhf+hdBBMe7adwU
WAofhha90Dm0rqD5v70XAFzpB7ICMYKR5mcx5NECCllQDC9JiGNWHYwGhkEMLEP7Yx2BstukXscE
1ikwp8DfFnBxRk1ITOA7IHKJRYCvRReRIKCoaFnd4dbiLEMUZoRToTk14DB5JZZY9NjG0wouWreF
UB0soqqRHa7tznSvxcs3Pb6OF1Rd4WZMO6DMC8PC0lyc599O/dyuqVIgpgL9D0Vw4EDAA+KX2e06
YPcxSwrzWHdmHWSETwNpqb69XU9oM8ffbvOk+Jb2IJmRE4VZqFq8LU7znzEpnF6jFANQweLo4zlx
2y4yVmFynadxC2LYLdvi0pyhYYwsiHPH9+KQHFydHXPCrXmxuBtgcenkpLj9pprdGVVGeiZDzoBs
JQac5fxZd8ay/5PkXkkwzzvUkrxLQ9daM5iZGRtfxlboNKEvk7PoJBH+zad6Ou882gCjEnk+/DuF
69VGx76EbRNWy7ggMxAIUXlxqnv3Wbkx9Y9dz5grUIuaGYGHJoxn63MeJSXV9968ZNRzkamSAX/2
ihVyP4sWbs9SOFQQHLPlyGE8kSv2Tm0FQG7kxEY0bvEhoHECdPcb2lJFUd0y+HSJh7Qky4MG8W/h
BiRsKPUdiOEpt+HVL+je5GAiPAGj0e+0DkHrifrJhhYVJcKp4brV7ZiJMcmR4km9swmJ4EiR8gHx
h6zCRMqDksMeFpLRC+EFQmtagYk0y1fXUt5rEQQLp0CUo89LP6ElhZg1ZosVEWFmJUdBMVE9XTkg
FLbPTPvfeE38Y61OyI8IdvpLd9MgPfVlv65+8v3RY+Nniza/rr/1RVHjxylZX9skd3QP21LHg3oG
MOH+EQjCOP/mPZ7l06v8RgVmqVRO44kTaK6bgZ2u4ecTq6TKLU60VD3+q4XUIPtFK+D3SlxXJt/O
MRakZ1hMC0Rk3Hzvi4VGHcCnrCCGG6lf3UZM5Awpf1xM76RoFQ+sTzP/E+2TKPrG8p+8i7QugClk
++8Z4QrBY5yYHaxDVyW7JEUXa7uTn2XV0/nDmVyTX9JRbYJUkQ1fCWgiWVC7VGL6aOimRkIQoeZj
LDqP5v2nlV0+8raS8v/5reRTsnaYLn77xDBsa8JsUuUMy4Arq6X1vZTKh9+pNVSPTPRDCuymZd0H
0edFQP1WfrwEo/I0oWpgyAcApf6R3br3PGIyUVLcNPTJ5CCk9cIvWvrGtCT8opIioGiGexngDad7
/5EvUtBaVWH1XNODcydk3IedRZ14+U6Z87enx1qST6MkRf9uwSlknCmPdHeRAmSmsVq4qS1UaiKi
kIJNatGEqkT3tOvA1f6y9fIODkkUWNXkAK8nSoAsnHUt00g/HhvQO5vxvnvdKnFTGGHs0VdxByBu
/8Rfa87qk/QEaZr4Kkra9V6owKrSGBgf1bJI+dpjZsfZuD9eB6/cxaYq6UvnhvpkHPx/IMqCRtMp
zlnj8a1kXFV6s95ijvjvcMvZSt73jcocqm3tFYixjJEzLwZ4LUMqN5va0xCBw5eNy+5dwcrKjLdm
1/79FqPqWuDJZc6s0AuxLBcbN3oPaDYCS3qdXi6ME1FCUyemoIZ6oEaW+q8yDov5cZvRAMY83fdh
DzfVRC7DvH5BsxwLGzv8ID9KHQeqUXo2Dc09yVcDZCFrH+t5C9PNYfyh71lZAvRl6Th5fmxXWyfk
yGlKW6BBIOVdkl3tXHik4M3HcbrLy/xKHX5/sxVzNEIekVjChqXKfZZfcgJeMwpQ47EF5jdoZDEm
8lb1JXWrIZeZ2/C52F2vE4heFPAesBCLmsVl5w12M0BKGkrXqsfIZQBtH2yjc/UkIyJwT55GlncR
e13aq9HV6jWFY4C4rk1iC2BeGYewZ2FDySelNmLyqt4m6+FNrldPajgwp2xWlKFZHzn7Po9oCex9
Xc6SRE6JogiI8Gkqjj3/g35xBmAEFAZmo/DBezS9W7XQVioO7oe6CoiStCObSwlVDBwdJBbF9DP8
I7DTP7k3+5jPVjCeS131Ttsw2IbL4St31N/znDMGZY3Jzkg8F35SAFJcQoo6NSG3JHIIiGjznf0v
Dxkqd4IJ+9aBsL66S9Wjez9gmDitnv6NFQ9uzVCpD7ropAbTSUeenTKq09C9xNXkbQ2n1TG2nGTq
+4AB5DJWiqLdzwXuP4DBuP9l2nxEDlxzXTMF8svIriczgEkmN2WB0fNjI3f/sJm958bQHzfI0Dpf
87DR6jAbzO/UPgFDh+ic+4VCbTaIbh9DTihFVGZrc+PTzWWam6jENAQBx3ZDjU+Pykuk/WRjsVUV
JluaGCqyjSv7VAZAinQpK3zowfwisc+RJo0p6+zN6rTC32LKvzdN8U6QH4v9H53o5uvpLJgWhjBe
Lb5SrVSGMBBadU85tn55VzCdXTH/6Ha4IlWTOHncZbwKp1pT7pPBlfCKRdALsorHoA90rWAni8uT
MMUd0tcVv55ktT1/h0D4qatYTtstd7x1/UAD33PddCEpptxivON/puKI7MCQ0EnP6aY9lC0q/Z16
bE05xxigOtK1Pi/gqU+oxvtROcaUtWav0YgKqxSLGq6IV7wM16yk152PoWm6aKR8H180Elb2a6T8
BR8wecr9byViZcKM78GXQSYAIwrTtEaBWOrNzr/Mev8EAbOHeFCVs6ELMBomaKaW3Pj9suWDrAoJ
g6uFwXYVpt2uOfi5pmKefkrKGqyilFNBGb27rnwt/iKD1t4T24VqxkD7xAswif1Cf7B1j8VtHcEV
CNRpY7wJMZOgpm/561jrc2+j0mI4FTXfSRmwXKeVJYV9gOWMEVKbDnr/P5xHZDZ4aykxRTEF7xUl
yemJCcbkT1jPUz8EZPP9UI5D3eYRvwZ/WnSrQxRXFSNSnxNcnD/VchxFJZXX/FOJ25n+sOB/1Voh
7jgq25dNZFYZW5t8V4W7ZC+OLSe6P8Di/Ruh149pcsN8wuKWxgLL5Ach6NWFUaBrRilfJkIkSPoQ
S0j3e4GMvmCaLg69eUWYx78yP7RCsmqZq30is8AHd7DYUmMBqnO1vCG8bKVvcNVSTM+ufwqBVMjL
c2g2wweiIagEwtH2esEWU55dPLQfrn/e2G1X0jUHfvBnn3G4z3f/TRHsn2UrzS/IIs9ibPR9z+q0
LpHcTQbvC9/shRNDZJKfKNJsEzv4xcZmI4nJWSF5cQLqYs7mvo33TLpxlDaEQQcHxWipI+oppVM2
Z0Y7uHlinkVfI6I5T9H9q2icMFzhW2PUsvx0ui1OKLiAZUuR1+Gc2IEY3xLhaan4OBmGTG7B9Avd
YrT7bJGemVBaAwK8goC6B4qAFcoX66Vvp0sCzsQ8hz/HNLEJOeVi/cVmk+Almpvqjyo83Vr1Q6Ye
UF/jzXwGQF88ZTQmTLrqRU++REojiB7bYLNp7WkpfbiSjCOM0nmVLH6RZ9oG5OL3hRMMLw7lNTMM
0ULnncrdh9R97QcOtI/qu7aE2CHdEI2fGnv6cPDzmbDKFL5PIbel/4hqMVCULv5NrGSWhv/f2E9a
B/HzP3MswdTsY0Fzq0hlYEIF6y1J5Vv5HhT2OdbANCR+lVowfJ53i4LdoeVgMf5OncSU98c3Jnng
mxr5vTLwkHIotRmzZn46nXiAF6UAfYcv3G1c7hxuxt7IvyOD18ZeoKWyenrtgmqiZZEzQR62FVOo
aC1Q6eLqNldy6XPqo6M/aTKvTy7bYZ++LLSYtO22SElE9Ugv0TQXdLMhllDclX5BQfQJJY3/JpzG
saQVwon++SBx4ddXAVtZeaCFarbJNL6QlrzWgPg5StRMd92UNUTzD0i64l2prFPRnpV3oBC4YonS
/+VIolzK+SbnuwdTkJkbHFV3py2f4NSl6OfOJtzqs1u3jF6KjwwHpJhpokvxv+wWV0vnbz/xjsOr
eGB4gMCKH6hSrrqtY+9uV9uZlGFNK7dI2KSP85ImWEkzP6cCctLzS0Show6SlAVvX7lIxo+5/7Y0
EIXqY8yUHR3fUueGTi3GemnasyQsyXJxPh4KHaAQWRfLyADnNRwfAgHeBbnli95xgBiiPudvR3QL
QUM7lrj7ywSznXf7X3PBre1St6bsQuMPdyMoStaPSLOty0RJ/PYNQ1py6ZRXi6xxc10YZCtbVqfx
r67d6mEiV9iP7xMzIFkdt6SSGczjmUsq8toNxMcLof9Mc0Q0L4zJv8XVPgGlh+buYN+S1OyRFzjI
oleyN9MXbEkl6sHHRIVY+jJKIsutflLORfuMz3m1ObTOJKsN40VkQmkQkMlBhyDvQR+7lKEdo0Lb
h+2t6syiYsL1R3kUEbxTYHGhs0EtMAlNiQvac2pE/FbHHu+0j3sfeCOkmaud+XP8r2N+5DZ+SV9Q
CfVxN2XdvLmIFwkf6172vHF5SlJCYal/4g9J5Gr7pO45mchxBAGOORdcqmpWnYGQiUi6f/W6B+nP
Rip9Y3D0T5864jJhCzoNafyvsPaW5pE087xGS0Ta0AyDUBq3rXCWw891cVL0AwCikQnKrOT6h3Vh
/+4jQ2M9V44nEgjOAiRfRRX6ETj2N/L1KcjW0hVh277VQudS8iZYKkm+vaRDR7+1I+0GxPhQOg5I
dj/5SZa630+vkBvr6kwOSxJYBeOWTazaf1zKHe4GokgfvseQBPnI/rN2YZC5MtUa0DMYosQpzJqZ
2JQ23+JpXS+RhgUoHA2PgCM1XgZTCFmxZ8pWKFp7fsf5uBPOwwhT7NVxA6ugUo/vOfDE9uDC7LqT
QzkaBLMOmXSr9z58bvbZHA3vGGHRV1rRSL/Qb0YREfjSj40tRyYipClCHGWOjlbrlcpa0fFIBMOF
eYXkaN0SiCX5yxXntPO6fwacqFE1g0RMuoYctvFqYoYUCN4z0Yxn/wv1u9Zobr+AWm9f2dXg5Kr6
kSE6ui9XXwNMHqxOmyBwBeOkyxzrKm7peI7G473EGKjTw+wyFqyIwI7C5PsLEieyFAQVq14SyK1R
NZBYKjqRnOYbkQb0i6GrSmbcQoJgzytGT5E4rwkdU9B0dkSb5R+hLAB21hR1jiZoVWD6dxMw6TRL
Fz5GEr3zBV+KJ+15NGFdOAfHAhEE7gmAbKPphyl2YBDObOgbXXx3GygDKrjciYY7mQxPt8Mt6jLZ
6oor1mMrvOFRxb2PSHslnCGw5RuhUrkzanx9vh8vF6A5iFogBV3czNlp9bqW9i3YH3p+pbOekjb8
Z77hhTFmhBnyyzqb8kr4PMEddsACIbsS7OjmwJHxzJXMkE/lXvOfQL2fQ/iggqNZL8dwhHFEtjMS
Q0m1PmzaAsX50PyUaqhTPIdCiWVZabFUEsrQUkKxamGKjAolcX+QNx11RRcHQbAWybh5YIOzS8oW
B5rANoeH8Azr3fL9vuT1e/l3+CukEMlQif+3egixf+X63J2GKkG9rRsx8hfPr4zU4ObnaE8JSmey
Fv43L9vd+1FwjLiklh7bCerrTAB+mIctUe3sVjHBcSpkRx7ZQmTnhYrmZjvjq8iaen4AZosSSLjq
VjQ4fFdt2dT+8siirOytAugLAZ8Az87cbVV7o8VrDQK99U/6OPRtUJ+WuUebisVw9Ptocl1qRGrj
UL3UR8SjCNBJ5cdiBykiukknGABwIOQZp9RstntulB1Kf7fYcZSJszAV9AMdgIAPKa+MWiwa/bJR
IHPlADeKkmpDqnsvONZLEvobL7D3G85huZ445Cfpil8tnFAxQJy5UNkooHOtRHdazJikm/99mM4w
7hxk2avBU/IXzCbfLILx5nARLr7MXPRnxgqTRqiLoqXoGFLd79z2R0EcARMhy0Bwx/kBsHqrDPWe
y0pD02JbxYJbDJPmceCopnkhOCwwnDgFtzEN8dMqUe2N3tcMaSsz/eBHb2DmqS4FTdAdXZccVjnN
t3FhLDlL2h+tnJJK2JDxkAQxQKSUZa7tyJDAW6Dcx4S1P/A3Ix06em5pBCvKrYUqM9djrHPxbI/R
lQzBzc5joBwmVvUsuXtZwe70rR7aD0sDL84n7fpJphez+O5LVU1n0sMdakM8ck0YaPkkUhd3+/Xi
CK0muurJwFZPX7YKlEiNnfqlzIXb/OG25JNTZc2XqYuqQG1kW7L0XJgovJraLIibePk5hTXrBv5C
nC3+Nrlq+eqwLmxfblLjy3JqS3JhDjoyzrYFfyrvMOBqEe1OOLnhWlve+g+/y0f9DEqea+VvFsvJ
i/bzrMjZ3umH4guep+q6k8ho8nOP/yh1RB91mpztNk3On4yx5cnqP1UwTHSbR52vLPowXE7E9cri
WrNKe6/j7X7rsBFJRrZT8Qz+07Ry/1aiuuHy8Vgh0APddm1GorXOB7E4f7iQ0XsSlQUnx3wc2nnR
5us0r3CquOCXyyv9BwCBe4kf9P03M/oktjENmAiH0kRmYxO7s0TwDrrlp8DXJJACf9U63lENiHP5
bv9BGUCCIusGEoH1wONZQstu6dMTSnQSaFUDJVO41JGWW649HMeACtzfVVPFHACAQR1fVoZGj++E
YT3CuQZwwCEpeVx5kNfS0qkmn9Xo8bvieov3iO9ehJzBiSbyZs0rGoe55QNCPtLcMYS0vBtba2eS
AMS1L5w8rWkRIkEUQMm9SXmakkqGf9G92tDVFto1kWWvy+0/7GOFr1icuav00zZyqepWOnKf6SqW
pyQfhPlMOEtlyXN701whzMpnpJrf/yfc5P+AqD2GQEfLO70WRbmJZVUMPyErK9/NMB0vcbE8IAzp
d+wxmkOh7oQJtajNey62nKGmHTOvrIAdu7v6XceQUbOMvtNfIqTaPpecF5DU01KueRyFrt7KCfmv
G/cU1OyS9w01qZQfezFAvkp7iBIUhyjA/47rlHft3CLIybZ+CvnPsNphBxGsy94xnbem6j25WOHV
/vfZtnVrnQn+2hOPQplAMMc0t/MgoN383jjawhYNmvc+nvOXLpn/SfQZjd/PxpG9ZwWM/q4tHIRD
JZVjoHDAV/hCuDqiOUe3pMRfxqHbA5KegqzoIMsTsttEJGaQYjFBA8sOV6RS73gDSvXu3lARbouh
xXHHqkvRdpjNAI2KZxOtKQKOZj3DKiO83YQisQFtF6f/mVqAjqeBhKSrkOcCUFWqmH51aI2/2eNS
dO6TF05DTZS5MWmyvVdu+qMnBIT0r4W8HH0mecoroZEmSgJxu4fxPN2+PA6kas5QhtiU4xjz8j1X
wkFTPSpHx0pw0EL+xujeywQC2qlc2+QfbXv7AzP6+5GEt3dl+vsvpDSwo4qEGfMvNvo7ufui2zVl
J5cFbMRQO2VntmFJzlSnf6Z2LnVUdVhtYnTf64eQJax6CI6B5GAYW80LzwO2t+eEKJCeZ2Ci9TaL
hXOugCpyAXDWZPycAY0uOievTo4CvUAiyfzc7gF84bI0pmrMKghb8IHql49/j1++MnB2pjlr6+sU
C0AzTAt3wEJarH9pflFW1HIDc/A0UMi7f9ukVlykSVxm8QGstFw8O7y5rL59qgTAp4nmcU24w/jJ
K3JSiDrqKOsrpw5XsXPHSFKIsYxekVlEX9CpHt9/aSbZ6BgbxfbgenHvj/juEwzNQTsbS5HIuBs1
gcPZ0qbNGoFmga1VDdgy/3c8GlYEAZjMeP/Ze72GmMzvMXt1DvyFLelZv58G2xryu6p4h1ih04C3
i2wIaGksViUPpTAlu32AokjKmRcrly7PbZVDFI9NtX6Rmka0mrVB6MkRFkuPQUITeWux4PQiNKUo
JyFOKBYaROnHRgR0Uh3dd/5SCZ1kF8qBcA7PS0jaUr1nlOyJIGhS1F6XGWLfDCJVtFMPtH+6F1g5
lUxzDnN3JlrBCdGv+GAvAjwEhEMBcIi2Ihn9fFBTWAZ52vPipMliVaWf3ePBQErK6keN5bJzrNUe
W0UyRiLrxgdp7YpXQPKPMWmeN89SFvXDSxQOQmoreflWYplwTtEmpXq7kN2+PD7XpM47Mf3AIOKc
loOZyN9pomXlgBmeTNzV3tK3KB+AS2Ix9IMtcTzUwFZu9yWSCcio+5A3fY5gTanaPKy6xFmcyMS1
kEH7Ecz65pUGiLaWtgy64sZwKfDoWkr9xQjHM6TNz3D/h+1Y1lGyq4UxfPgEsUHlc2Bd/tqPoj59
Y1xESDVV32g/lNMbA8UwZS6ZhczQZuLBy6KFjAWwIdvTMKEuDF6EfdNCnbHgZ4NM/NyAh3RfpkPe
NRk4OIliHf9ZVQE55jxMKpm9IflpqCggHQzsx+pdDxdt9B6KUO1h2tXBaH69Jbli3RWC3z9zNtIt
THpLhGxEfhZ+yvcsKrWreoQv8DOR8zDdJD5NlIXpGVKu+jcKkwkI5dBMAPjeal81pzde/ajYrLfg
wDZ4eueTVnYenXCL9PPVKOROlUe8dokqPNeMCn5xBR/1bwvuXJJIwDalT/3RcGin3uh11qbCz08g
5hpD6gsRZdmHUCETyjMELugbT972WgShjCIeKo54g8cwMHicQNPsKncj577haFN7V8UeZHTWzwGW
+iGwy84kkXQ9n8SdSPnPwaLjOut6OLA00JWZpjMSAv0P6TPFYGjqYKdIOkL5X8eviRfaX57bYu6d
fG58iN/xd6iymSznPalip+vgbKZObYtYmZVbIvnyfpeU1K0rIRELhg8cvj3XKn/i/kGDKBkssavo
3PIR/MODDd2dMWkB4/5upvvd/3EzpzlQn7Wvfv8oDQ7GlwdsZNPLG/l6vdyuEUuj4ThBl8qCA4g/
/DdXusISo7R6RK9J9RsTNQ/XWc/ex9mt9hy+3WT1Tz3FMBQBYy3AFreuqXsD0XyNDeXeblFr6V3h
Lz/bFV/ePVdDrbsIQ8//u+uw+AjGRLMjo47n9juXABst8bFQqnJpbwCiahPVSwaN4/XoL7p6nu1/
/1FYXXUnf39Mcb5RuPP2p/x1wYbs+uX7YfWmQohKSXDZiAi0xuNOIjLuVHoCoFLggPz0z8wLg6te
wHHGImKzBZWnnjjxPkZV+Sz62NEXZPrkw0mZ0oBJte9SBfCXE02f/oIVqN4k+NptH4MG4ilBqLXq
tOxQ93S9tV390Nro0fVyO+eBqsRef+dZxnhe6ldvF6Poatnu0gqSDaSTXpsp3x1P2BapOo58UTji
/CD+SVUHGaFtJNOsR3yzYmQxwAOhs4Tit5k6oaAZ3Qjkyadurq1rDZkfWIKMkM/5jZEK3RE7//my
EwcKHCLhz87nk9Hg37i3VMcG1eISTEPDDIImQlcoFRw5CDyzU7h73AadyiUVTQ/fy6QA1M/P/sJ8
7Evgj6Nng5CHS0htlPVDHPMxQ15jYVKYlPiECvHWieT7tGoc2rRWDtd/GPjrQ5iVZ4IlGC/QnTd5
BSHdOQKEK4l9+rCcQhw3JfOkmAXuhBZBETx/8ShhAfjgV+Qc8WttmYwnQP0fhezefpG6Ef6dOGFO
QCEmAxF8AGoxk+wpbsmV69DvTKhtxRep0vGdPuMHLigFE8uqzAqVGpaCuVwWbbubhWCARRvUjsy7
MWTtsCYNCEgss5ItpaeIujHhwB/dw2CzIR1P1gmObuopLf1yuRUb+rQ88WF1KrUgztiTobUMOEWw
MdlWhBjw2yloLBXRcPsDk7aA5xtKK8TGKJVcXxxZfb8t5EyomFOcj+KoJzV2IxlFd10FR3OQRCc8
+UhbZ/U10VB1gU2AWGObb8xX0oD+PFyWP7VEg3JfxMABzO7oTVtfVllM6c/2CBEaKGwK7JWItIZu
dYZ2U5WH02Sffz5I/tO6ubz6wVqW+lSe3U961Jck+vHi679qpU/CKIsrtinJIWmMdw6bny2KX7LI
CbhRCcEoUK+AWt5v+AIQM5LP0uXBp4gtJ6U/XIpyWhmLojXlNKKc0wREdchzk7JQPdYUYMvCbwKr
GLuepQG4S3Cne7oN+Ub45NBOXGn2CtLHAc0KYrw3RnDzcBDx6zB4lvFQMerMxeHVwYPjl5D4w/7T
FlXNfBcJhm/u39iPEkfGEOafSPAp7ov/UmQY3GLMzq2Vef1FIkYQauDePRrodoA5kjNU/kn4sM2b
obMxKdnO/NNvVysLd0vzJkYBOcvC7cX3PekLhLEMKRxCeFELrjSK9lcTidPxfUbhZlAmhdHypMz1
FdLWEgl1axChuPtU4jfyNBZOVh4x5PDZ/d0211jE0OzJTE5PWfmuoZMLqPwi5YG/Xi8oNN55vjPx
vXrtMowmYEex5aRC26cbM7rLWncLlMa3SfBuEHyT9A9ToyTNJm+7bwKXq/bnGXQynrwsCM8xJVZA
ucG50JjTxR9J0JcrO9H4HYEeUqPe30Gm6w5aFBBZ5WN7IosvSyMKPZoDIvhIwfprpkKTXqukWlPH
Mu67iGx6bEH2rRYUbPyNLm9bk1C3wy9k3m5hXRhJ9YSviw4A1uk2ePObqwHdiIkZVqiFeoL05H3a
j51SrJtPoll/0dC2IRH4aILw6MmPbpvtjpXgoH+g0xckNUJIbNqmKTBgbrDYm9vFh6znFYoIGXeY
r7ET7QZegMgV/SX5zUl7mdFCawRtf4Vv1UNldQHdcbOdFNoEp4+o/gH2OuDVn423DYXt6ljWVa5B
x0wrTOgHrn/G25HZN1GyUnDLQSZ4MSY5R8fS8kiMUgg4RfmKbzNZ3aUwPyZdaAdjstTzQdfGdAz3
Ah7jwOzY0gTy4QjUxo0oH7w3sgvrDOT/2OF4yDDJ4z9ne7udBbisEXDFOlFYCmtlpHuwOqEr65Ek
d3YA9gwC70gEtV+ypckb2xMUYR5caekDG0YTkbbbhbIOSfM2S52V3vHyAkx3c6C2zioMamAuULHd
z6mOrwJSBIXTOfGKHnmh/ch+P33zn7xC8ROYX6HMnM4UZTVNoYVujkD8JKDoyTZTLZ57+T38xJBC
Hx4EihA2FEpFZLgcHOuVn+l08xLHE2s9RhiLR6crp8k4nh2RcpbxUTLWzmj1Z1hgta9l3e98ElfO
LWk8kuBI7N5tm3/1b8oKaOdsEkFVAhEHN1mF4kcvfX/3o2h/Smtaam2GCaeC0WVnPki54N4Y9rIQ
/J1TEjU4wYIEDAsxBm4aZ8xREWFT0gMRuNsY1gjy6thZUVDCW/j9Bq8yhNRecVvTmT1acVRicIDZ
pYMT1zHeEb7Oz20IQCu/hP0QqoDv3KpmNovEOfyxDF7ZjqL4rWAagXIhnpAF2fA/pSurKWP/nZO4
jluDBxmEy3qKDsO8DVDUjtcc6Q4jeASblQLMusdsO2jb8VKkEyBAAUJifX+JGbdV4tver2GMroX8
iggEpkaU04oDhlcG9er0O2F7mIzIaYzraewrBZeREyZ6OpVOoqyfPMTwi+9Lqz89n3uUVxfBp5Qd
PcDjmVQX18HeEGwIWX0ki80qrFSHys0GbJtyEJXn+RzHhuRfuAHuZecSBwYxbjJuBCyyJde0+Z24
gtEKRs1WY4Sf/sONcBeh/lak5IGS/U3CKm0v7XpsV+dTcljgOi90mAQ6Ez+SSMQxL6o8OiMOdkNw
4UWCv0c3e8lkL9TNhsQhjG8e1CuFj32+AbWFjo7QTgpiZDpQ/7+aDxRdTSMH6CAP2k8JqSgvwpyx
DDKBzgEvY8atU5tmyiwYULYsjSgq+El+8ZjpEd2dtJUW6NvS/Gk3LAjRGYch5H+VlRDwwWX1FbRd
n4TImrRLxwdQFAD60pRvvzqHaeUZ8YWkz9POaPPyIobi9AAxTs0K9K2oIPqZ0y6VDO2syB5ZSwwh
pRiql6vBO4y8rhuQbvgceOVQ6cKrZ89+kfbGxZejhLOdz53/swTSzCo17LNbnWGnzoxpK3L112Xn
wMnuc6m336dXl2ZTGazZz1zafdyK8oQxxT8uwFKYFMBo3xO7HSIjynYwEe8p1wQpBLJIaySs9CIA
GSppNdBpFjaqqD8Zo4Ms8PyURIXTVCWucVNqkwDjnEK3ViUtZ7Cw6IjVaeATe9k3IHD3VfzK6ncw
OmhCxpsq20chIgl6L85wTDZNRh4NMpDXz1/xGODR4uUt2wtxyTmN8hByR32kXbyeUhenadXyi3zx
wYu/lFBdiwFQnUP73cgrKvO/Wrhs/l7SlKf1lI7QkrRo9x2gLP/o7RJwwg4lPObMVdUmsPx6NHws
Yc8/YLoWvttLS55rM+ZTmq0n4NwMDRr+LwqydEBKhTuYgW0xF0zk9bwc2S8hAeEUXfe+8GKcxNzl
yELTfkJdDPG5wO1T5mAx7R2ecE0FjKr5vOEscxjIIuVJO8sJi+kN+mtWkJsOBDZbZZXZgjeEXnj4
hgnpyfIZ9H8dgCTVJ+JAnD9lezN0JQ15tUISogKxYKH8mBszgsVLrxgJINF27XuKuz1ISRQ3yerS
MjEZ6XDEc9BSqCkV+Zk/ZkiRryd0Op/+3TJwzPvoXv12Yc47UtG5rpFa2ZkxKBFnrEg/Equ1d8pv
lUlAMDRwkXKySuCypScZX4sxUM49GdPHNSUcBSoHFBqGAMQgcz1itEngb5JZhhp2MFNtXM/vDL3k
y93HBJywBYrb1wlZzXkvR0blI+UKuycF2A9SiivQtPzGZnybLsS//JmHXPrfPMQrogsxgfmZXhOR
sqa4aaGsQ5B6lGAYLPXDZwqt/bNblFGNxluMkB8Ib13mf0Joujf17pZAlCaqspV6jqJv/NO8UB9r
PQ7aRGHjR8qKbsbu1mgkKtKR7A7zGvkuiSSh1tyrV96SVbmSZmEbXukuWCmFeegmIjPJuwm8kuN8
GeKEHozgyUOYRaVRYbKebO0sS3VhBRkRhwxtuLftuHcd62a6/d2lkqRJmE7P/4S/bDqA4ycFQdql
X4AyWCFx2RI0p4MdiPeZ3OsHqpGUSC8lbbm+iWV0Hti8JUqRZbYzybDS8CLdiReapzl/qXvHMI11
vMBNp7663li0WlLidwT5LV29EgUJIX0s06OeP1HC3QloOPlH9eLqMpgyuftVhxQ2ixNRIjU4EM/D
rWt/7o4obscOsYFWJlVKIBqSTx/uLr+3aRChPS2Bdhn5DwYVDADrbbKjuMGTcZ+VQmFcA9BKOuGJ
1/BTYHJnFpelNRXomAd8m0VXBR9E2Hwzo0HbujSAXdM1UCbhDZ8o1KidD2jz10PHP05OY0taWvK0
TV1/dLVWP2XL6mmj3nAMHvlyMBBuwV48mbL++RRqVtXbtxkntpwTu/0jV10dFa30pjSlqXqmcE/f
m2NNtoNb3nxOlxlr1wp0HlWdIl7U4Rlws4pY2ETVeejq0KtmS5I6r1SE/2NGscppm2ktiH8axWjl
VYfmHuhY9izovCd3MOg2bD80Sd0BE1hZnIVaB6QvjELs7bI4khs4alOkiLQARXO1r5mxURflBs7S
if0NcxOoZ/K7dvDywEYnJ7cYAd1OjKu2B2HVPOPv0KDg/YKRkLIT5kCRmCYPLWYwediSf+GUZA9D
t9BxDFc0+kV+uSm8Gs4MSIriIbGpBHM22LjjTQPXc65B+3DBotAVn9VSPY60y5KX9PnxlKeLqufk
m78lkn+bEQFAHVPjV58o+CiAnehV1YKYquMOsiqkwEvFpJ7NjNoDHjjrSE5XbKvnrKNh/QIZc4l/
Q7Pd0d85xCe6HqGOcWzh3lAijWKahuUbzQwdfKsuAEknG9/V7y/Sj06oaZ/YNPCkCfaKZIT1wLoN
yEo2owDfPbHwyvdnbp2BVi1lr6eOJ9kC7KijYc9iF64UwsTPL4qxJ3P8t9YWnRh69HN+n0blCOEc
9aQVVQbUI4LXZ0ETShgd5CBCpx5zvrP5o/zAE+EGSDXSWA53iSeFA46QT53zJPIE/0Ppl0kaEOrO
CVm1SYDLKhOjm2AhbdQuqVMiPwl/iQ4dU7oGJcBBDG2vHu2+f4hD5VDYuiECc7RBlaPYcTQsCtsd
8MNB0m7bLCjpCJrsGAYOstZAWu7DAOYHORDrTg6nUCuOSloM9imIH+BgE4RjZK1lg8JDQpzZIHHX
KTwwCvToYPfi9WJxFPruSIkK8qCq1GCjEXOo/Zs5Mx/aXcKYlPTVZfcbb7bKTpmstYEo1gz64bPB
XJEL4+2FQfq/ovAcywDDY+wkC4TKz+8Knmq4PBMoSTWKj3XN0zDTCv0uGIIUGJvImafzLdkxPTwD
sj4m9U2Izx9qQ5CxMSVOziuIGqOelGFzPpf0OZjHKD3VApimWo9QUhnsmmT7i+Tr5KwFA5mybNXl
w+zPqf8kZGG1AssKM8xbaP1/F8FIbqWpWredqy1QEeTqYsSrZ+QEqX0OyEpMqKwB3ROetLdjoW2T
gdycWRB3XCCZ9sr6gz3AnkeIZDHHo7WkJRBCfQw8o6C/RoSrZqgn5utHYWv8E4XemOWKKOG1fPjr
vb4h3ER9L154IG/X7HPGcMHw9C9urps/aEk1So555+b7MF8gonARBeW714bdNZLalMfOLXDF3dwQ
DeYxM1qAv7crqYD6qu7/tmUrbtjEZWHucGO3DucFy9d6Sz+fMK4SJ8VmUFV+qhoFDmN267MM7Y97
/iB2FRMLmiXDxyjZDXLm8kxzF2vquCpZMBJj9CwKKTLQQ8IjLRdL1VdnCoNrnWYlXsX3zqJxKgrn
kq94qQQ056gGKVBFxlmpTv4TQkgZ31brcZZkdPH1Q5Xx6C3VL7B5k5/aqPvJAqK7ijSKmcBGIfp3
OS6ERVM9ItGjQ5O5FhnYpKYOg8wG0mz6AB3fC1YFgKnHw+5De7leLIwBsdfUs6W5yqd8MiqafsXM
aHc6Q3BnTIcAVYduRlZAm3MRZ98GzpSQwWHvCnJ8lK/S8dCDsEtJxReYbyx+zxvI8bVjuC2Ed1d9
hulW8B+ER1dw6rR27Sq+soRdstVtsxLEftZ7xbaVJ2DDEKNkoeA0aiSrZ1hKfn+Wy5y/RsiHD19n
bpTpo8Neq/O3DfB/oAl1GG+S6CcSrE186yNcqQMNfYdIjn1dHf+2jmjM/s/kdQMgVtjzWAlyO0ti
2EvrdWvXt8xpMRow5m8MlJIlHYIvJEym6K0wicO00ZcYhm3MH6p8eRMrSyK3FDMt0TxCPacwC9u8
mPKUN1U9pU3GdL8HzKxXo4CmVZBSAs4JyLCUvJXiPIGdAn5KUCChwF3/oiQSaPQN23rY/QxpmTDE
vq0jh3G25LdXog9ZWfAGGIBlZlg6x7jaoFX1/7B8C/Wc0EcfiENxFgHBELrNmF4JEbt5Wr6E2iMX
pHVRuHJc9zcZzOZwT/bzTvl92M0yo0Mr5fuBV+LJi/6590BCbytkib4Ken6PaEImmDeE1JP863xb
/4lgSiLdDYYuZp23wcomVBx/6KpA5wbe2me/M662uqExuhc/HeSuusHpkEqSfRFwdEOwrrmhxefa
EMFujklmU6HsomSOnJcPGShNrdCZMzuLy61z68Hzho8HpgdEJTlnVat2yw0HdHN3fPHABanL+7bT
HAhd4d0u0/3yNZoleD/vKjxKQ+QBZo7/kdpIOXbBvFIt2dWNDj5dQp5w2jMps8hG5qXPPS0IWfvY
ltzIkEI+8T4eYdXBcdR8QwMEC0tlK5xk7rPFrdhTqQcZGndmaI4QIbj28t5hU/a8Z/htI0lVMdnJ
IOs03rscXo5oLeW6Qx4UHbNcTfTspj7g+6cJSKeE2U/2LeFy1va7V112t09Ea6hYZE8vI6vMsw50
e0kHnQ1k3ye2NIhpdZzg7Pe4/GkYZnaSEkqGLgeVmz4sXDYPgEXf7B71QLTo6Rm/5YvOQp8c7Inn
5bhuV/snq5IwMUqEPaCdi7GRga9kZWpg9Ig+hIyKdj8pfTDpV1RmbVwpFmH3PN2K3luovvPKnWuk
DNbCPggRDL8CKCD18pkBAjmiHa+Q/0FY7gdljmkKufUvv1gtXZ2cRZeyshtUv2ndCD1MwW/4Cx5c
kvy0m909w8CNv8cogZHPkRZJ8zD9+eQg61DiHBr96yEFppS0Qt8eunXOOV2NU/XZJzd+XwlktvB5
x7F9UoNiAwyEaL7OX0e3MGeZQSyJ4GmtKdkAVIjMNiTEXi1uiUgvB56xRNJ2kvvLesvLMDOcPfsS
uGuTFwUlHsZ1OszpfiXmblog6CGEtzCV4/N+VzjXM2Sly5DalvHt6yo1/PWwddsuZeOmRXtzaeE3
WTsfZxxofPnLV5C8fQ2xafhkc1W/L1s8zJZZedZHhq0/7D8rbqLLVCOxo6bw0m/uHP00W7vGrnx9
SslaLL0MtFGqS5BPgKNDKQrouvnoz++xGu/c5FprV07LAsEJcIXCLFhHLRveqhbdbW0z1nAdPIpJ
FiGmWaV2Wef/NJQuCEt3HxD/MVPnSYVfjMtTRicQvxg8k4YLLl3m1yMz2omUKIC4b2wjlB8Ku6F1
hHcpzltNG5uLP7rRxScAYxDfFLkyN3TYnx/Jf95XA69Xhzmv+1ewYeF05jPjmYB2mSMAIOAD2IQn
e51IPDdsnI+pkv9oouudP0sfkkgBjtUkrcogARQq/sNI8ZFmqD5UqnUXlR/Fa8XwCqL7YDlEmIBd
dYzz1tQOTTntdaR+eIzUaQqyY9hH1o1GD3OUrps/pZfgqECU/0ufVF5RmVAIXBXH6f2kijqWFsgA
2NcXF9GvVDmNdRyASmUHgswranA1zRPOu+2yKpH8wt3+5sqQcxLSigsh/OvnlCVsrLvX0sKN2YEr
GDZFAD8GE8XdWuBpoqOAJOS8ocTWf1B/MjCWt3I6Nnn27nc8/e1oURcP+256AcrT0uL3qGKKn719
dwwVg/O2pB2yT0AoRQJ8ATD49Eg/AQJvEbSyquoZZQAlWLr9GOzliqXI4sRVUgaYC7EvD135qKos
kWSilf/EtBg5+9KIQ1AnK+AZOD/j3urw0g1Gh1/4H9Q0mXmMbgf4WucI5ZkUv40dxyVObNoJmhy1
Qitme0H7fZb8DSgk3zcFO9X0ZQhfwSg5G+jwQL0lh1oSOTSeq7+8JHvAaJPn4p1adx9MkArcJLOj
0EHr1rkTukbKlDlH4zseVftQuadglLrc165oIjXe6l80FxvcA1GSw3AsRcO2FLvFPfjHndDHrZMT
HZFSrXmHEj4qzq0nl90JwQwdxpZUGUNQnZGR7f0ZVCvREjueN1ONf0wO9hu9ANzuXdWTBG/LnIzs
6IHp5Dum5LaH3ujsT7THFsi1oBX84iKWU3F5fjvZl5u/2YhEhylMUQJWAG5bdwZmsMTmUBM1jTxw
o/SzLNHIBUGe9Ji3sH47FrGILrALu8TihShfgHT7AIwHxO8HYc5Gdy7vVrw2J+iP3RQGqCiMI+Lr
I32zuPPipgwotJnTdwlqdI85feYC8aztauCW3wH1mKMXURsWOX5mONQRzfkDI3/k0+Wc/m+JaRgF
cGiZyLD8pj7NJL9eDMIXp0tYjBcDL/Hds/kto00hkRo6Co23LIllXGqmkbGu6NKPocRUZ+zpevGy
UxS0+Fk+5lyG0NnoMFc4/eEn+xhcpGbM7ViqQ8Ux0VoEqiyC7hkhcda8BAxU50bGEKqEJgnzmcDE
O8qTZqauPlDCIWVC6tz6Z0m0+4y7yB0AzUTbWMAQCRNsRLi7ChxP9s/DjOAjJV7TAKVUkDNEaw6X
mNEe1tpuBZPxhtlySD4oDxlCgEN/eJwiBhG3i2JZD9gpawVneQLBM4lv2cI5gJrZmbdHhinsgEy6
wBx0cy3IboY/weL3mDSd2OpiK/USNoaQbnM1om8whAvToGi6hF+jIXpsTJr/c3ZAc7LwtizYtE2i
K1jDQJFY+GFpwfAOA7bMD17aeMLGOP1WyWcassRsWyT78VQ+d7svpCeoYgYvy7/ajD+lKRgNtpba
1DS3yqpK2evZmBfkfWURtRTX86cQJiVUl5An0ScQncV797HMkZrjAtz+2pap4THVIu3Ld9Dtg4jr
5Jq1L4KmApYwa4UHJh+CXhL62TbyFwt4A6vRSJ6K2rOWaa7cfV1btIzY22HyvN1rkgoAYJdBhY2q
nATpSKE7KuaNEkuIX+ccdqyIMOs+whfuq4QRwcQ51qHIOHNwWI5kF8getytYPf3GsAD02BnBv/ri
zlG0WA9GVp+/uD7ezD9Ze/DltVa7k/Ea5xreFKOQP7F8mAnkuaqjZqIbpD97A08jGw0vyg6eCYGQ
pwtjf7C2IkPsZXTU5sD7+WXzmL0B4KPm9urm+vxmixW3zuHr0wWCguQYjDn0eMUQ1NWLMFjoyvvf
it94dywjoHiG/cISadJczCfYPFpRicQj1WzBVIMQlTAGrGRZ1CAmsMYckdzQBzWtoh9UN+jAEL9c
2/ZOYhFPziFxfArPB9dBo5q5p+zIlDuD7gCS0xAH8k+rt0NwzEoA0i2yeecq15Y0Scpgy8e1koSV
6vgRfoLlBR8YAygZEcK0zuvAhY2TBAC5ttPrFFrqubUpPddqMhD5z4C9BBYiUO7cluG6ZniWHd0a
qxWI+otRXfr7KDHsAeLTK3kuQ/wKzkbBJef0TNwrBu3pTD4VznOQPLOjUudK4nbwZ5Qn/CZmxvuP
0JmnGcGlBK8DFJr7ghgmbG/gUQmfjwrZFaWitmSmECoPLPd3hsSYXiTHjRphwyc3b19vkOJgDjOi
XIzOlA6VXj/GgY5kbt4lfgIkT1Bh8UDQ9H7iwrtkLYWhsKPS/58k+QsIkIDzk0FFWe+FR+ZIkDWa
bPV4Nb9Sj2/cfALTY/OktKCLijwlpifI/iSjvWsXcl9eMzye+cholVzJh3h9hjkmkhhvKhOA/3Fs
tU8TxCb7qU6FDSpOhvcbt6pnbC1rCOKVWykXvt0QPuAGzx0d8l0xxNILvTAPcjvgX/zMnAKSZdXs
2oOvvjfoQHgEc7sVXfYD3BYipInfXXw2JZr9Cb2BSImzThN9IFAi2Hm8ux2mCJHKhi8mwsLngMTN
cO/tRTQty1iqz7WGoorvQVlPH9QiDxFdF7oGygZBqG2sXHxKZz5OM5wXsg5jgOFz/E0heBd26C+G
FXgBzsV4zZuMp9hXFqSTHc2jYXSFuvqGrKO2itQu7ZdA1c+0o5n4vn8y6PV24xQqBI4wqgd4BzLO
EjtuKTUjeRJ80/B9A38qeEw96d9aLhrnYRCkl2iYugmzL7Fc0rkM7rT6AKq8+WY0EWKO6cjdR85y
RPW+pZwaSsvM0LsDAM02grSSNKK0vdVl1husRLbac25GaWonUmts2Bt0akcSvu/Ej29YxP2NITTS
1WTtn6EMSqT760Jjz+ehyKE2YG1NpfFW2cCTVduLQeUguTrLY0t5VZaFPlOfmUq5QNEzkSl5pa4Q
S6ZZrRYHRtrbc9vJVJXNhoIrJSA/t3/PIeUiZRSo2l1howFre+Zb5FlELufzGxZVfrljlARXd3wR
CVxJe8mn59y7HoqlN/0xtwuWrl0pl9XWX7GIG4Qk0FLd+06vYeFXVlWYB1rt9QwXVVH9XUHAg49L
QcV1LXFraVlrxyLKjcJZ387dpWSKvpchMasir0lbeZ3hw/NmnchlzSSpZK8zDKNzq1ITKYVTnbId
AffWqKOMqgiASR4N7KgXMvuzSCpw6Cf81Y5HdG6BkztL92+FI9/wn5ZlKh5+nPVrNUNQFiDjioKE
YygS2W7imiqbM69qmid+hmHFtLrf36MG5lF5USLeSs1w7roXqWPw4xPdoSHLyeJKH1Tqx0bS6mIw
w9+VDLU3IFsub2HjdRwpHq2SFBMrLPUXWxNZtROMheFQX/b4BUkoymOkkEjSaoQH61Syk5glaZCK
b5atmKkaO0o/YAggqDW8/lBGrCeevlJ4biwVSqapMEt9rsnIp2iRM+4z2Nvac/4sDQavQcgIKNQO
EC5k3ioB0V6CM51f4pyQ9Ag/Sgq+EJ+0Wqm9Ng4xZWMKr1AxZGXqVG3+7+Sz+jOM0M3vm6qj3ZOo
/IBDd4ry3PNvUyUhKWOSFJPVd8JabMk3XjQKFrs4S9bAtBQBgmv9SqaP92A8Iy0i0GDwJ2kcrOvd
xw2QuMAE0EsdCtiq1Uae1Ntjg3FXdQFr+di7+Ietbl7CeIE4I1y8l0F/PipaHkW5t3kxqWRpDWw8
olgWgAW07UGgse0Wbk5fPDKrkufviYKBX5nNHDm7RFuUjjIl1V1D1utsFtXPcNSh40ibCol9rAw9
MwbKCj08ry2s5FWt2o3fAQ1yFMRqOmgP1rTDikS7KJwXcRNMN8t8NIellEIEGWcw4h8Y5kMzod66
2htd+iBMLt9P6qSX6JaU7QcizmBljCn1+QmDrFy6ErL+i8cLhibd3HnFM3MtgdXhNr5PhyaenEpS
MEq88zFeZkRbxH+qQ43SAon/kUzKaTtsHgZs4dhIhYzo8rfWZuJLtLlRzNFohHnciz/PPw7sX3ic
k1OtcDt6QvZJ9v+x7CLwhNg39rK53uys4vdK+uVBnPO3u0Dy5jWc0ZHu1ZLChv7Vbys5QdxkWlXJ
XUTtb7NHOJ6wB5xg3LbDJ69wkw14pEnTikPRn9tlAxyBsWANnDxiezmoyeOqk55Ud2P4LpSx7vB3
jivrMYeZZ9Qc3RdSH9LkB0HQ0d43xBNAyJg/QZortz61m3kAkD60z05Co3BfcAkREZBnVz/j0/XO
mT8AMY8PpVAWFQbI2UbWHT2amYqxQwcAjDv8hfu9q6tLF70+j2Wds+Xb6WiWfMSHHt5Q064tcgFb
aHxladVk/0D1w9DmecXG+1R2RSWfrzd9AwssQE2siQG0jLMgpmjJZMMEVS7XhsffX43WdTq+bwtR
1761xD1CvWfakFIwuRhBKkgM0Sklh0VZeT+t9tSq9Nel7B7YWNjxK0x5p3rapokLEeLZ9wlBmpKf
OV+1tTyqgK0Ba6qP1zjH3Ry/iPbCCsblje8+czJQPkwqxUw9PvVsQQpxgONMUXNsA06AH+DvKOqh
2CIo4NCV3YNx12Xe7CERllyxN7lYzfqE9g31gX/zSXz/rp3e1/laC2R35nd+zIVCPQ2vuvsn2ePi
sSagozEDiwPE9QCrx7bYIzJmt03RXnAUYEtXhy/QAIT224L5DlpokMG3dUIzpTplmSqyWH6B5HXA
ejMMv/xyp+qFf/vuQ6rAtfvwcGSVD13CW9FRXpWCnFapJSUIvdvNujqSzwmC2/DnxDvx/UhVEhgp
r58T+J3R3hLja4URnta5ypgDxXoxGxfOv4FOpJr08b96OdFINEfQm+t5QafxutaqkFtBXNTWlXXU
kWIGMcrU5KV+DHzQTS57qpjnCQoF6Y2wWv4J9kpAz34LxjHpZwbukwAvvxFtcwzn7LaKrY+14stA
icx/hlYI1mr4aWDM1XCDlmffUIzLAg5wF6vik5JtPK2gVqRPvdudV6Qyt3SrzhBfos9CfzkX6PqM
gPFzKL4QlX9tTKtcHUVeIx05Ebl9KN/92AHkIOwXvqX9HA2CCMomr+Me0vsIm+W+RxN783BzM4I5
SsyIbeviC2WHWZ3zxD2GiPEEy9uCiWovddO3HBXf29PDpV+mPcPu9GWwmwtSeK55Bp7IjQyo2nss
z8QTWokI/Qd3+CU4SudHS5oJZR8gv3O3//VoVYPivlCBSn1jDeIGwphf9hlUjb64vhEKa64tX7ej
30ArWZJ7yBWAzlbwy39F48Ri3vy16opeFoEaMSVlCPUkCyIdVnpXOvd0FBzzxS+vteAMhfAw/3LY
7LcWi/nMh5RbZMnYdbIFuD6N8ByVibJFHKTyEbF8eiN115dV1Z3B3YibKjH0K6DenHif7/ly7oXR
iuG7mSfmoHc7pk8d6djGoPhlNs3xKziTc5Xb1ajLMEOQKja4A1ugHJitwGAxpR7EwXkuD0zGGkfV
bqVWzZf9ecihPYJR17uH7rhyHCfdKyjr7gCHvb1aXG11Z/YFhagU/e4fvVfLNW4jX8Em12fpsp7r
Dho3y+I+XJdLmRHyhmKciMJN4d8q5Pd3h8rK8olQgl7t1EW8/6rsNGYAbv0/p0Yp4DMbrXC462fl
kOzPRgZ4B0y0ugETu1DCShFZaOJezToJPsnBSzH8akWEPpsuuX90RDVFrdr0GcZRvjKS2TEiDEf1
LPHkQmwNK2+nPeeuwyfa4mz1onYBS/zhEYRB9owM8MGTt/F2+xGO8f3m2eKyD+7CRj2z9Uf/m79C
Yd4BSLth0ONvxXEYkIAM8tFIddXWDPGKQcHGpk+ey4KaHleH4+FkTG4HOqdYzFf2EijNaz548+TO
eTnMLs6LN8Gr/gvGKsZKnWSNxb2yYDgz/8Lwu0YtGEBEZfUsxF3XmDb54pd0nQn3MXWwz3PKljPu
iAUlDfbGdqwXSrWNtCF20S4Ak+oALDhnJnZFVeLsG9/tNutzq5y1cqyHL46dh9txLIuKN5FLFVQX
DOp217qL5Z6FJ5PNGE8qqdEMtT1buAwn+7ADpoxbvn0j0cp/a6I9LXSRIZY9PdmaBwg5boi2VFw/
P3s7drjeIt3s8o4GocfiUINCRlco3YXXwueArVdRqMUpHShi/DZTKStBYtIcPTWppYyPHtbFXzgR
F7/tATFCMfj1MWQ4uLyMRDRimtinDRz0JaZ+d8QlQueNw2YjiNdIw/fhT/fUfflKjLyXWrJuR1a2
uC+TGZZh3zKpjJH24PJjJpRbtrqyiabthlVHY5TQazDhuUdu/vykl8VVby9czLeJfrUPeGs7HeIB
bCR803m4Tj5Kbg71ZckNwFTWUGvn63uYfLoCKESVXWbFZGoa34de+2k0TLumBpSUU9lNW45h+hMA
jlCNgClk12q8Bz9vAkX4j96hPnTynh0z5eJCh37pzuC3loIjliVkPZH89ijy719pNwXoi9mfpfr4
l7GWMaLoRtQhJxwxHGXMkSd7rY+mnNmsJ1rkP08uQcsH2qPyqKz+5/whgqP/reYgQIGP9hIlpbKh
hMGRF8qutV6mmBu1Jv/HH0lcE39QlMOppN3DR3xvqpMyhrb4lf8/N15uWa/CiRACpIOUgd+NJ0hr
Xheo3k//TH1pE4c6mbNx222sIRdmxBEK1YS8bLcvv0Sb3sZ56tbjC0E9oKBcAEsQXSC536PGwYYF
gJwETuWr530DdKYnuGj3TXrzbTdPnRv1z+X9Iw7gVJ+Z0nozOf+3/niLxxlzCvkVCawHWge/swFX
hNGiBiMPnReAxFESZ7EpbFxUP0AsZVgVZFbQb4pLkt/tt+mMORoOxSHW3cvSTZaAeuZxjFXaxIqU
1I1dVVFGDE/CP4iVLuq8Lwbolk0EIJwGjSphgbAjgpsmqiUyuypbPXj/86OXqlvv2bfvE77ZdTGr
kSeleAPhiBtxuKTMZJKz/oYnOvW8xeZAszAyrElguHZ7QUbE1DxU+sTNIHvPQQEcu2s9/iyNXDHF
le3lmMlM0z2Y5cPHNlsvE4h1nb7sI3sN0Hxe+JRElTBgqwRD9h0zMbp/r0+BxnzBtptZahprjioe
hWHnHxd/66xnLZx+YOTy17Wx5GhOy1gksWoc27ulbTssfEjq9ANfMoicdeG7hxd4ABRnd2aCfpvW
4+FoFXKkUUGeTX3YNePTPjsMBp+ipnK6fltecZK9RgtsYyxFNM7EIQmKJgW1qrcnQXv5NMFG1jm1
FmwymnBiJutB98zfquO7Mal2KkxbSC0iSmXv3HbS+P/HFxSUG81AzTtSf1QKV92oZ9ETds6VwC7z
Eh1GnHAAAqGOl5AmN2VNIy1T8gFrD+yjBAGQa2bW/SfeD2mipqNn/nAGAqLKX6l1pWxA0LKIPYpR
RF0CHvCHqfTZKONeGg4ZIo3z/n2aByQxpmCtY1IOiajcmhB4WFnqLJ2lQ8Uy44VJK3UzfO7welYq
vfI2Kwyq/LcpdXPRIKWqxjdeSrkJra6/CXGZLErpZC/KtXhKj2OduQ8UBok1i/UMHnGsS57T++ZV
4EWBYRqwGxPZpI3xkexSJrkJiWukoPOxdsjSoASgby/9bTk4xJdvwospABI8h+31E93dLBihYb5r
WjUtH+cNephNv6AfTBtGC8XOTYARK86Rg3DHAkV4Md3Gp6UH2qzNVJn1IZFBRJMAJZ5tUAfqE4xb
5lFQkqN+bwctIX+P6QUupYFhezue1yisKbd+kjoi70cBF1afeFDzQK+caW8rMR0rOGqizaQNH3kJ
jmBdZ+vnAaX2rMw6GP06RelfmNU46RHmz4rGvAu4lq5wmh3zwz7/XYhrRwzlbctGH+cSaD4C85vu
Qx4RR+H4MOZQJPAcAeOfBBcttbyrJWQfw70t4MJt8UfotgxLNxfspc5LpLTWeYheozhTX4T8eriI
QFq2UQGHpJg7mQO1aaXDy+UdeckFpUU/iL1ecLH0yVQMWZm8pwQUZXXInXOIsG2dADfCt+YP8kd7
5SxaWXvq7BQv3USgTFbu+LClagFoCf5wQ35NASfkNYI0WKvC8h9d5zR57FE7Bz+X3BKLNPSoql1s
p3Z/CdF/9Tq46GbXdUanNTQZcNM3UdkKOqBAZGJyoBMnqltP4RFptZKKCztIRg5mTwdfFq/6XRAG
bLiSu8jfz+sho5pp+dwmlhTml+/gIiiuvVlOAaq1SqYUfIaJD75rEL1XaFWEop5LPgUEguQBHjUN
ft1U0jngUgT44KBYpV/gAaYd4hy0oFYE/50Axw0JyQbZAoTE2rZRcHgEbXrtrP6fr6aApJMP0GCT
esnnSNrnEVBggdCt4BbwonZf+yW3Hnl56xrmxewkNKic63U/oN4EfDaIVGoZzIrLIswjy/8f4FUa
wVgUCvp7zQ7pv1Re9mOTYZR04XH/fb5TtQ7KbwR1c2XuyuFoOagD5bcuAwuvgwdTNgpfo1pEuVVr
t7yqsB03Fi5ybpn0bZYPMyZVpmc1j2Om3InNKVFYpS45XXfLqM6rFboott2IfgQHUxDlGNERZn8e
YAwmcwEWIm/KV/m6E+5Dnehx6ym7fEYWjBo9Zo5QhqFnoofVCMMNnYCEjPirXeRWsHGgTNEgtGqo
HwkTV3NuY973qJpMeh0A0IPDnlOi3OnT/byhuwWKEXtfaaix8lecmCyY7MTTugyc7JgXoaL+iJKQ
p7Wyokf8ixt5h0vZ8nZiYotV3fisQGuDjFmE0edIYO1pVyv7BEvIjnA68r8RNtEPf+KmCyhSM0mA
+9XpnC/ITUQwfmAwLSXjUhKOVN+6efQ6zbgJKsBtC1dFwMlI/DUd4ZAMEJ7189fzgb6Ti7dP6Hsa
N85DuwuxneSUKXAypNckLE8vEHWBleeeHqHNlqmbKMaSZLgXFf+pZOXtn9FhihCatBzomGMfIp0B
2JNiep/uxcNb/tW9cKu6p6sNMh3hMdL6rxgGhIoTPSm6+i7TrhTDFgnZ4NmsYw0pWY8HHqap3/uP
Bflie0aN3yscUDPj4eMmoZGjYWv5g3St74VEbfG8a3kY2s7l9DOxnHf9LUe4eofmx3B+TgsSXNFy
3XTIyUzerVRCWsc5B2f8+GDFbrJ1lrlq8o6UKn4v38PTVFoMDK/q9y6Yd7S2FPvqSv3B6Nh8+FLT
YWqIeNd8IdX9f4KSaVgip3Zya4bS+0FLqlfTZhvolPTLHrftJtp3MOoaHvOT7XLFwT8Lkwd+qKFB
mgdRkSdExtVMrO5ARwT0hgkvd7MdOETyjdDVt4gw0TuBCboFgt1wsTZOm9SLLuW68+e8cfgIwsgh
RUCBMExw8ow0vTVKvWkK14rjpGG+k//T5jORKJzhZav7Lia6qNFomAFSXmzhTB8Cq2CRT+ssxMgr
5ts3+J2O6j36jIanTMp7xJ8qH8sYUUpazcjsBjgZUVpNop6E1womI/vYa4iuu9cWoDwXslYzg40G
07js5umxEVEsXSdbRKBPx3cngV0mfCTld/EWwipQHgABC+AO4WMgclZR69NV2nFqjK5ZskA1Twe5
Myt4yxypGPOLf0I1thf60lrxaqKu/qt8+NzMeMgbj9KztAVB4hIX/vpvNfOyNPLyo8vHSYJ0W297
eIfo4QhczoVhsMwFm0Grx5ZDGd91gLoB6blAXPUr3S1VF2J9lewsl35lxcJYbPaDIq3oyq/tnldI
+NziIqXypqlMw7+5FM3mCuj661GoLm/HQga+uYblvu+2RwgBlFCqn7pqKkOSzg86IpmRg+iu62Nj
otdiMXP/VkuJKu7eNsaaRx1VGjvbWTkfXj8a6XgpM+0Twy/0q5eMkwi7mxch599QqBVloDYEIW9b
+sD36FRbL0WFCg+uO99T59tBuEACUCR+zs9w22hShL+3rY02fFjdE0+1xI31qhBMDAWkHHSVmlK8
v6dByNd+HFOSh3sgl9Ch589V1z/IolG4vHv28NFSXQGniUC/ZCi0kNlBBUlc2cH4a6+T7VCc5e3n
jKPzWQSgZcsP8eCCxDWDHrx2NzEWkXT3kznpsvmaSsK36K5lSXqNMdMp6jR3EQdimSDJDtC+qpy4
FTMRHIfK2u5FpfBb5ZaefQmAxGwHgcIun2Y9FDWcR+ep92dSI8Lx9bFEjxSSU4DvoHu6qLFz+brM
VeaZzvJf9ItvtW4VAoTzfAWIxRQmLJ1WCpJsgl2Guzpc2fmV+sNHb5QPNkHTaF4o3R5b6EsoJ727
arh2tdG5+k0bky4K4kH9PygB0vOjZT2XUcWP832S8ftgsqvg5nsDDHK6J1o7Cgls7GZ1M3nKFoRO
IbXz4hY3G8l9eV8XYcu65CkGV2wHDwhbgGpaXIXpjZ5vEBop2s1nWeHpHYKDmFE/kF8E5jUxgOdb
WLJDU9UqL2pyWkb4SNuSs7YA8UoawwhDxSg9bwOz+d/0uEY09JezPnFCtyC7aVt2149PtVoodpq7
1BCVjE4oR5FsThi9HL9lQKyFrIPJDf0L72zsVUss8Yc5kgr0DkdmPm+M6Z77rSBqPsbT5JkyGZu2
sj/61WiIqCBg2G9k/SC9ey1gn+QXweja0CDFjV4GFmY71Und05zF3LGZW0RApwX6Rn4D+6Vp8Av7
kNouEDWQas2d6zrrNbcWTDtkBB1RgMINH+l2ocYp9atBaUtNKntt6AJgf5TWBWZa/Qr/D+hGSAg0
oU6SsWF6XFCziDrJQbo+rmdiSpP3dXhIj85VYRnRwbuG0h38nluY7gSxFmMBnO2BPqiLIAdDC/B/
b/Nf0ijXB8Odtv7QopAyKXuk11q9NzoN4K2n3eeW7rx5Sh7w4wgA5WI0g28BvTRpK7cSg4GUbZEv
v9Nb55abq1oZ3/YhD+Dcf3JV70gtSnn+OQD7cuUKkHDX4K6f+ocyjL66z632Go6kXIVQuv/62r5d
dcuPqAgmIzoyVtOm24Hrw1opjhu5764EdYexqC4rolodvpfw+RTdDU5/7VTYkvxr1ZEa/fU1Q8Fc
Ii6UsQfHHo46UheGhJuQAhnghTLOEaIE3tT3ufcqeDd/Xwsgy1LyxIzfuaGVp3fmgeo7LTkHCsMi
b80M8yDlUuP7NNShUzGYqoEI9XfShoQ+2ohDXAVNngmww7sUD70/JTXkDlrcazKp/UZqDwRryCdE
XYvnDf3hB+raXAtXlGu3BQTLQzjUm2PaobRUAwO1lokn0vqGjNKfperW+yh7GUU0ybHHb+jxcprB
nzUBz61UkmKlhLi+dGaYTaNbxlB6ef+svlAq889i7l5v2MKJ29HAL+B3bOcwKJDPK7jFwCUPR8qZ
upTbahj5xH+6io/VkxVO0H0L9TAiG0Y/yl3uuLD49aY6l/2xzOgX9Ohmtt3LxjxOpBK6kgVVhwMt
dUzYFfzwPI0Wn9FC79kt92cHTNmayKXdM9rCXzXxDylQKfiT1+WzpPxQNKV3uqmfu8nc2dzFu92c
weig1qvWqWXQ6mIJ8ayYQ9T0lIzBRibSgLHEXRyz7d8Dy2wgbzWdGJWZhHf9Nl2ibAI1WR0rAmlb
e5iLYV2mqbU9MRhye7fKrIuNliG5hePD4KC/dMD9vwdQGmngNo+qpfqv3dFX1a1nJxvGmyUhOlBE
+iSHarkk7buZMz/EFVduErCZKfGd8X01hW3Jalu/pSxD3Lbrn8N5A4EigVh11LJAFHZ9/69gb7oj
9ENhNu486eytMghkGHG9yOS1x4nq28pkHEjECRQqLEpIPgKYJ46TOUPbh0WdwgInAh39rSNDf9ZL
YQN2c0Uv+j/Tqk8dObFSIUKwgT0DdiHw+adDrvAZ7bcx3SbrVS+8LKkEWLsJVaSkSQrJqAw3hZEe
dRHSZ+Abtq/3ErOjV6MxAyf/5rqOCBICCTj8cqeca5rfsXmVgfwocEnuLmcB6vyxbqOANRaLJ0yg
GmP2hcWMKd4c5Vy8JS1A7TVMiPUPttiC14HVGvprEi+TpfFIuT5JrBiXfusq+YrpzEYdA/odassE
BysTzg86k0d41bMB6QeOmUG7JOsCl7yJYWJxok15zZMloHe+7ruw+5pv0+EITD+ONkYvYAnTRc9a
MYosetCi6HwlHWS39mUYT0CsDzLHSk9s3hz9vYWFmIWqVe3+BCSisNRkWlHt3xctGpkyIl93bEHm
JHa2iErQF7KT5KNX3EweaGO5t+CN9UzYG+gEZ0OQ739y6xmRsTw99uzlqMdlIkq/brcWzVds6VIv
bQUo5QauSxoQSzutv/FzD5iL0Bvt4Gx8hGo2oEfLrylggrVheEX/F2WQYOrAKpCoCHWqOEO7zMrS
3K4KGNTTjHeowidGGngz4y8uipRVTqAGVOh6Mbvi497SgDbxIHq41IdeicFPI09mqgatmAyyi7H6
AukHgJPNYD3iAE7VD30LUoH0NrJp064sDB/StSY8qR5GMDRcczl88oLX4YLtYMEVuh6UUjaslXjB
Hx9rbfYv9X6LKkKisx9OxJrTMezqS3iUmcIxtuta8cXpsLIQgUEVgrVxIY6yWbMF6PM77iet9kqB
mGwjmhEBOOg7RJ1z3l6/0iabRmHkzoAPrNk44z8n3s5webnqM+6stTVbWDKXXMma7+hhJStxNZ+0
WJ3drSO+Qibg07smkgBdBOt5cR+IwNDNVwmOsDnW7MLAzwnFupxeGErKh3zV+8vR9IJ1uMxHFops
W6je0Dp27OxlJ4WFPz/gqd+w1Y6kSuzC1wSc1aKqJAwPNOidpEblxFXtGtljnPS8FLBc0JRs/rCb
RUQsRFOcxvDruwxV6sHWSz56iBLWVUC5oF2zx7b1lHyDXcbIBd68c1Ll7OMn4yvs3m27tsWOkAF/
wF2hub3sTJwmA63J+maB6PS18l21QjwJR/0xp2pH4k8USX02eoZg296uu49Pv3jXqcSmgTy3t6yW
PMAY2JEv2glsyr+Vhdtpk7lf6o7HlTRSnP1iTvYfWuiGZtCoBCcQLPs0LtUY0UsMd1iFuPCmgNR2
WXARsbJWcVf6UdQdeglgCRXx+YzclCoj13jXiEuTjTf+UCvPjePA3YDAk5wYnUYxjGgmWCag9Ulb
+8GG1hRNtL5N2w2LOU7E/nwdvLRtnRvVQRyGGtDtOc9R7p+0IUmXamTzuMUMY9ZUqH/9HNZ7pM/t
FAdqpA1psIvI1BYuyCLQ2HtIJ66lkD8WU9eCqbDkhVnOgaxBEp6jbhigfu7G2RQZm3GlQRV0pW/D
QycDQZt2FcOGKt1BAYHcenRJ33da7t4v4t5Q7JUsEtyumLHGuY4BblI6iAGHSDzivJVvU7/SgQLv
oCB2DhB2pPhiF11YNhNygM/cpMexG35RLa194iy8Bxm+ENiILO2lQFggRtoXuM5LT5dh1FKRcsM0
ggamNDViP97hXom5baTEvN3mioxDvrXgKtNXrFVwT3hIgRUHhMf3wBHjWdoKNozo43byN6x5Wxj3
lVGr2QjeulJpZnQMssJZegOGfxdHiF4KR+SN2RjJU/GLNveF7rE3lMPFkKBXsgup6+ZVSRla5UO5
J/IpwTgdes3YJT3KJsFSczoXLk1aA0EdlC5SdveV5903PfyhdBMuPzw3Fu6TlEyHb2S4YBxspoeU
VCW20uv6aSAYFDEpaTYZAirEWXVg/gw5Jh6jqxP0UwJ8YStEPsWVajv50DZocT6Q0aLHwRmRewGA
bHz1efUuEdlOkgt5uhkK5ulfkxBensjf9pQ/jgvVG4mNRs5eILYQZ0gL8ScI8uSkJlCHJFHc0d3O
VcAfFTlTR1yHsklRR1egmfUr8NVGIuVgoCoi1jHFj47bx+yyHHFZw/uIARIaKYSJ8eT/4nYU9HWu
sQFH+MzRrjSA6ralSozL9wcCZk9Na+ByGj16sAYrWvmFvQ/pggPI3OpRWGY7+DgK2IqM2fb/hCYl
mU/ir+SJOpQunBHCLRcTbv6ZSGDkD74imKzO4q3BS3uHC//+7q3bXmamkv5H7znVrIVM0AcmjFkH
2gsrY0zkVmBZK3RfOdVJ5qa5cpDrAwFAvw/62NB5e5cl1P3v3yTfNekH6PhZvd05YGBTgiMfEeM8
Z3wMHwY+i4sOiGHqvBIkL3eDuS7ktWic4Y/4wIxbwhx05EghVci1stw1lqcFrga5lnNbMbQ7Tyb4
4GoMmJ+AzAKxoCC7ha50uhdELw76r6aicXijKdoBvnmMAGfG+nW2N8dAnnkHvggO32E1VjykUEvf
heQlAI5dtNNGitOPT2LYlrKWUcJme8c67zZywSizUq6DctxJKh1xaCm/gvXAoZtt6ARdjgSCc4U9
8DDNuw4+Cmcz5etuhgwFOgwp2PbzREOPS5JPN0OF4+8/UrsSW7a3I3akt/ALZ3PJRLaegr2DrWFk
FLRKwxm5yKQmIR/4khyrgHvBwT+Qpq/QCC+/tmrPQQuudpu1orcNJ4c4mrRuqny+4u+m6eBQ2WjN
eJ81TWCdq15RfFxTrn2bP2/pi/silFSWHuvoR8rbukVKlC/1YETwgQx9zCo4t/Ul43Eq0ANP8+rx
i3PgUYvHjF/6fUF6xyICM3HOhWoF/IDnjfWYPBOmGKaLw/qh1ydx3b/XnBz9hlui6k/TtC0PGQYd
tcftaxeQBGgU4PoaYt4pyMcHaMDt8hV3DEB95xyuHibTUePbnFRKcRlTQHEWa81FHVwtJYtetdXW
I7AHlbjEWjszToxarEf4uUh0jquGNiucCIdPzStJZyGy8LCOnEAIAw9Rn76CG2jey5ovzr10HIF9
9XonZtSLybxgo/3y8lSCmeTjDLqtTd5uP5Fbc1BpALkxVcm3XaG5ZvZjkox1MdmDtwmU5H4FjAYG
izbguMu51+MCU+taroVxM5wIldHTW4PQRXsSLgp2LCBqSE+b4/Ewc/EHGgrNEzrAMltYOx+IYTDf
5Lo3UwsugrwN/Beb0/HfPKAzZYxZnvohbivLUIVSJueE77NYMwZhQRc41qGFDb4VnLk7Abcte11r
boHrun5KX6kzYqf0YjlnAUsuxtBTmotEaypfcXi7d5WjNfAV8IEXqrnnindtCQYfHhNca7CTfgfJ
73b8IpJFB0U1Pieo1/8bVErglSvwKTDsYTQCDGkRJ9Be9BYSkj+LbR6fZyxWTWMqPuT0f9CkHrIX
02WmJQEOIO9B2vIInyWOr/hMBMG8HyAurob6LleKbNG6noAQEQ5HXtpzAgnGjmt0+XfPOEILNI0/
K+qADq1S8G8FKkLM47V4ij6Ir1k8nkKZXbd35dwUoVfbR4T1HjajgU7CM77f3gjPMQm0aEEobBXQ
9QXvDN2slah+XuuzckzCOwb++n76D4j6wV5aHiDo/fWs1RTfDaY90JEJNkHNLN3dNitYVTpblQQW
0iD70F7Ed9CMGHCBgt4tpirOjVi3+VAUcjFezu355SLZg/kZ/eGemq42SzIhNCT9fgpPGvnbrWoi
ghiNsidSMpBLzqLzOVwkl2Hr/0oO1Nr4EyNdQn0jL6Gxs/5Z+pJuhUryYqjzPUan5lc2Cf1Cp+m1
Fuxylcc8q0wEMoBVax/TT1ol3w4ImZtPhw2QzjP9nQ5vj81FaC+Qnb6unoXxnnZYHlIfCWpQueVh
UF0OgwXIY99oxvPud4c1xsBDiE22hKBr3y7sUbJ0SDJ+anbBNz6Xx/rmlX/32bCj6CoJLBS9H7o7
cHx9pQB+RAmYFUQYHsEkRgRO7KA6Dgc5iinUq40boyTbAfKI8XbebA+1N445WIU6oihhl8dQvrC6
1TAMbRofo9YMxctEHltrBYz9BaVGq01/4G98SlXBMpveMamC7g3miK9IeIBOyuBwDUqwnSA6unba
7EemSgJlTVd2sgajbvvqa4AYVkXbcVkrSzPC7tbNC1Q3MHUdgu3og6D2YAEBmtgpmq9jkutMh2vI
ES+8L8uuUghxqakTg2hCv85Fpi+wZDm1FvrANBO5Jaj9o7uJ1Tg0Po15QeSH9gXNoqPXNYdVFp8Y
sVfM/SiJgKJUCNLCFzDCKB1A9CyfsXw/ygJQEI65DAfZ2s02D7cX4Q+frwjS25Yo6LqW/dU+ZKbO
WQfSo4x0If5WhN7QZlbBk42nFuWLiUCMG+K63H4FT70cbW99l2N48HT+2Wbcg9YrNW2Rw7g9fs3S
f1/+RiHQjI5Fvlt0KgVD4zZyYB/YZo6SlTq15gJJIYhJvUMoMqrLjtFnjihZsDOW3vQpnwWLnLDd
lekCjvCXoNB21vHc7moBDh4WUPH3uvBCdpzsOJqhkVa6wJhwhKL5FdMzxCak+SitvwP/oHEK8nsF
3KcdTl1R/uJs1wWcwLxoIr4r4uFIVONOZEi1lPG1YP8NGXj3B5tPQTgufSV5vJ9FGkJqNiVoWfU8
4ZMg6TWlHHEP+5EizeOwniBdlTKvjEb11oZhmWR5+gCK1nvMxUFbXFUHibBtHzZ9KKQF4XpIIMa8
Rw4C+C8bbV0Kku/kNYFNz7g/2kdrJXh9RRX8ip6dHOKAhioS2upD9rV1joxU48whgXpWtZOWYzCc
rXble7LmeBmNpz3aAMEBs0OaAZyQgImDRae1ILDVl1IR2VkVY36rTRhlduvvItGyMPhY48sNYgt0
1szW8JQfDhGZzZz1Uw12WB1p0WlzLFGJY51bL8/vsmfpVfK8HS0UIXa7JKPPkdjNmXqWWnC3w4bF
fn2keK8Lbw8hMDal1sFUzy2ZRlOPMou8dp4/BGJnPKsLWcBTAs3f4uTmaXb1lZ0i733Z+uAsGQJD
cryV9XeGYhbPBu7/BQTdFC/0UtJKObefFm7muChHTayn6LCCurtvS4C8dCDMBhwFBJo8uF98+TWZ
LV4k3YmXKJGHtPKJsqSwRehcK/BeR2UDGdaye8V7baXSwoV/0XCghr1P4JfqLRS/Dn5HROFL/tju
XUoV7vjK3i/aeGL7xtaphPUzKGeuKjopOQE7pp0LJ5BFxFGQlyiRKaJZiQhvj7DqCclfqx2Wj3CK
bvgf3gBL93tV4N4rjUlZ7Q8s2Bqp/TiKyf6b4bXuXoXgX+rpz7m3qO2EFVJcsOEs6XKY7LuYvGpN
dr2NLvajGt5GdMkYGld3/1IHqq0sfBdIj9gfB7LQORCpVbrVShGnrdVFxhT97BsZCoc5C75CfHxu
gvUO2rkAOMCBqF7rHttlui7+mDwvT/MxNrYKKy8nTW/0Zh9svB2zEQD7h3DN9ubiL+KCBYuvhBpF
mNdu/YmJsQZT56cuPG8ma+PonvKQ86CUeuTkfatmf4D8kMYlAVpDjyU6qEQHn9PWjLHP8WHV3MXC
jZg09B7WWhmJFSxwJKF+cjsgMucYZzDMBGuGnVGaNOshho7dqHmIfQ0t359tRFNOLQ+zl4ol9OY2
Nybv02FnZfpboahqYbr+eBpWFuzxfrG+lyqVoAIAUnsJgorGBzFAR1XapOYL+YPFPF2RbsTGLCeI
A0xCzM22Vrz9G+aVmsjRG35isRvWAbi5DA+Y8slPn2/p+dDVVlvFzbtlcxx2f7QqZc/yclWhIzXl
3juhu0KZWSmgBBQY5ZuAc67WiqXNz0OQM9i/QUoC8YfKis6fg8clFaRYkaPbmtPfQvE6/yjuaPv0
ehzeoT4DQedzu5fUXFrzaS0eSvZd3vTqvz/L6haRpAdiBtzJqFFxWmueVi8bC93tC1JZAIbri7aj
0njh7TOXmkyPsi5JRHkUZuut9f6r285NKlwZXq7oGkoh2aax3oweC9f1iW2AaH7vq9tkixudAdpf
VpGQrItga0tESnfAFxKEFN0uR0vSGnxoOhRoD8eDIfjro1cPmNWxd9w4k5KEtnORAWAO7O4sfdkk
zsEPHVyCfzOSX4tacTVjFmia8I+ylDuBxzICce3mOpgVF3UMudoqwagWoyTQjseWLIZfHzCd5Pmy
Qe/J1ctnDk++qkrL05tKr2ysY7Ggoa5rTePj4xj/FKO9BmKveJt2pPyHs96uGItTu5pRjsYKZ677
vELmnpb6JgWcNiskk2mrIAbFJgeZV9wa9KFEiaHXUjLnbJsHx9zv5gJ+g0PX1dC9XR3bhXj2qTpS
qwDGt5Jzh+CkwQjbKvFEkI9YNzGjTK0P4wJtsydgXHnmAAXAKWH+4OyzkIpBf1OY/wT0xJqB1YgZ
8hnwChAfmfe4C7x47sFfq7TAGH7Z9pt8Q+Eaa8EofhLcx4w+JiadSYdWg+THNHd/9HluxHZ7MfbC
0VlJh7HGmKajqiWx9DrGUrUP59gKaO6ZmhP8W+Db7cM7gz3qC91rzcRfx7YFTqizA4jnHIQXXszC
N5yCzNF+VB7mtQCs3Z3CNhJ/5yYu7cgd6DN/ZzB1wOupvXGSLKXQNxPTztTca//CJk87FbGj3an8
teMfDgp07HCpOcUGfpXZHX0oJRbEbpYnw7QjbbB6UrsT8dFKvfZxaKEqQcnA5rvNTUuyc5AfWZaz
jX4Zz55zTVHGUt0usl41AeD6s+TYKoVvwLJeMOMVevvVp9HmRfkD8Rx9keqZ4FWG7hj52cBXN/ly
e2LAO4yMhcN4XjWOTEepVaS19GHxyQGlmcvJ4ppKY4T5qifm54cw3gzkNT/DGALOEmhFGyu4dMP4
269V51kfpowksgOz15r/tT6Cy5UFSdxFjON+hVPLzbxQAFtXkruINRaPOjwkojiDvWn3no3gkLub
3lO/w8rSF9l7Bg5AUpDk6Nn5nPQDen7Xz0s0YsKTD7milakaQKbojMiY0s0vXGM+PZ9uE943Bt5P
lcAjEaQSXZ//ECKMC9+5wjfqGDurE/ytA82HWsv3/GNhm+BYOXjp7/zHr8rmbLgQV0rK3Fth7Hi9
MadnnCJf2RlBwDu1mtqGFedGKwXITVWUzULLP9YNWPH5Pm882mpy9U+d0jUsZLNhRCBTQseNwcCS
ZcQwYtqE28LDwIPKFiYj5toZ50E1AizuWEsyUqCd25zTEVNmvpyF4zMznt9w9//l7LtyHD4TFJKl
E9HWW7RGcvsyjNRh0XLJg7YM8r7UEpj4rL6nXQS3Pkree2+wwag1ggOk5ubjcmC1bxyrezWmDAUn
CPZkuiw9Z/8ehv6k+smbvhHN4Wv2/nqz0wXGLDHU5nUmafz3LLZJJAokxFnOIlVZp6q7DX3jJsmd
tIit08k/DW2LYSjLXNWi+ZwGf6Ob+06mh2CObQpFFM8oqSKOirJ2j2Y3C4dIDSiG5HkjVppNxQzC
LkEL8gUj6y9lZM8bAUHD3cyxsbsP7AnDcbE1eyPkdW9yaAK4AZxHaG4sgfJ33EwjmxJGh8XsENBX
Q+dMOHr0ukboLKrfkzsl8AL5boyXMuONmsBCPFchFlRbCEbk3t1a5fXXMsc+5OjCQzOU42SOG2Jg
GWv9meFuUdJf9mzCTY6ZCBBQUVxYnMg6xtcvzdgjILaEo+Q/77JnjM8/00PgSh2ACrp+MyJ50md+
StXCWfZ0MK+c7by13+Vo6ajMdr0DhQ+vVp47VKa5Eq9FxfJbS4GtsWr9G92/PFXsPXv2eWseaLiq
fs37yGJIxr0NiXPIWMMbldka6dCHQplXszqalDYGyLlxIc2KdHGPF6c+qFyIAD+m5y6U3KUXkX4d
GmzeoWCzIC61nWyjTzIZcsGHUuWlO3GS1jAL9280mRvSz/En1LcqNiOi0KeRpDUW+WiituRlh2zE
9kS4PlDKG94wrljubI/nRTEt/f3pXcVEP+q5xS2FO/oFfFkFYY8jbsMvGWoJzCL3NXN5t28ha075
tyYQzMLWaxgKsU+q4GuLVLaNv4dZ4w6CNnjGNQK1zfdWw6KoNZd6wIsWHp2GPW8fHZUBe6s/mNFa
7b5vLt7QZgtlzFnFsVtRYeocCXY81n0J4AixT9H/PXnQtS/d1cKtgPnrnPEtLBIDWKe4GvgN1d2r
9dIs9B55VI2SdFv4b+/++qX7atqfEh/U7Ul0U6HgEIPksNWbZdsH59PiWu2vKydIe8IKyaTqv5CK
1a28f1xVtZyqaIkCScesnnXXwJT2Ek9t4fLe6ZUDnWZpiYaXS+4m+mS9vUOyNRgpDeeFQBZGFaFs
fx8RNetu5djT4luyb6ZxH+2If4XtbD7Sd3RsMUdQSp+Dm6ldG/7cS6//IOo13EuYrQWS9hUjOThB
WCgahO908Mufp0mX4CCDTBambCjoYPxjjcKuLsbc+mq29Yk51DaRqglSwsDVknFDT+pJ9nX09zYE
uxgZgNGAqrwyF7kFPt8baR0ssAN0I2gjt7WHs4C6zct28OqsY4XAcLEebZYQccyBeDrkk5sL2oq0
mSuh0v1h4YrkOycXyAAQ1Ebp/wG+uN84cZtcTphQ64omd4PXwSkLbtIslOxpwCx7ctU4b5N8VOw/
pPG8XyOrtyhZxce+XPIXMmkCZ9uqdXDWh+EdoqYtC8EJJjc/r37ZhTWhmXZuJqmbP9SASHuyO6al
Wm5UgND9I9zyPcPHp7c8sDfShdKP8vJfMnYZqlBqXZyyrbqVQYxeiLUXOLZXGR4s4Vuae3sX1eFx
Tx3oe5VN/PuBqF8nwbsu88xIzoM0v8fOw5A8Q4EgFebE2zAPBgKVGsECf3C/mCzZQmuEnINvgGKA
QTKnkcXDE5H445n40ljYg5kxHZ3vN+y2jtte6KheCGpcFWLU+Bsxln5tFhRZZ2NbOOubMnEyNWT7
hVaBcaPOYz/bq+Jj2xSWbgQnieyFDWHrK85IccNvndf5/25VisNYLEL5ySTFlUFeIHCcZVt5Rzu5
+HJrw/4mtKmTHFDazDS2t3Gt90bXexWa1y8GYV7Cl8gqaWtVVq3HcVkkBHo6DHnJbXt1/UaqjTQc
jdvVeZwFunm245Xer/+UIMhvg1GT/y/b7I8Kg7vSwwFCxeWE6JQJ9i2kxzh39YFU438uRdSR8u/1
yjh3Lmxn/Uqm17EePmL7bq1BIO1+uH+/ssqik6JOCU4Khk1/D6gAfIF3W87D0M/jPfCggTM5Fo3a
cW5LRqypOOxkD+Nq/qZi5aTFm40UTku7h9/6N6GRbkDfaAmXf1L/nQcNwsCji0gIALHomOXL7umt
8GtfUgK4yskDuyBzJPk4ViBi/TpzsljyL4RM2jVF7uVTb6XSWwGhrDW75Unq2IZ0o4VInYANc69v
kEFlcfQHeV5D9fuP9M/CIPYJqrRFFOOg5J7QB439uFKf23o1TnjRqIUU/WY9Zsp3BHFYpXG4s27x
ZHkIgfGauryoOgwXjnQH5/vtbD2+KqgdW76qLBtz6RlrJ+tmFRDHM/iIY5Qp11+bFnxIPx1UlWoW
medHs1pOEegoFlyO4DTEv7PQM5cQ9e15thF2oyFVkgsSywfPzOO64ba8FZGm6L9XEqP2u4Al+vDa
eCYOB58crgi5gMLiyMqwK267SqxXMOAivy1HzNApwNUcDybc+hvud1iYJdkqUpv6bcMow0aWaPIB
dY+cJWlfQbLAvXyqkMP3xZ8V0r/rp/5X11NYP7EF5RaeurAVWD0E8ARq/bWsDwQBQMmcff0RgvX1
XQAxUcuDqGPc0Q7AU47uVwq2SvaIp/7VPRqKFioRjBnsJ6D5BGgyWxIRREL1VhMJrsGSISeBqWbM
WINc0RvPfDGl8LCuDu80E7EX508h2BXrhEv8ABmKsaTy/7Yb1jiXD9mWBPxvt+fOCdra5vRHhaCv
Gkj6ixtgHtffv2ujv2169ivMLt+JC8jW0ixPdcH6MmjMJnA+8qYbDqTOgJ0/tiobFkvb7Yc0t1Vw
ZCEebq9nXIo1Icq92twuryQWE9IdcRBr6csrHx/pVtMXSp/oPKzlqRZj6gK7UGZFbdKsUByPt5WN
CAkli7Wvr0XvAxvUlXzDDgQI0rgTAdN98lQ/7tbI5vmCMp+5EeGo8lyiqs+JT2iSSL/kx+gQU5Qz
PqPd5KGBQSjitNAkOIfLygni6nWDRuZQlE1hTC0k293GuWbjpXXz8tL+/gyehUZsqFxWWcRkeo71
9Css/9ebQ+w/EpylKm3gxnA3I2dFWLSV6qANmyZo0bGhLsljrRgov99Twplw8lTfKfdRhiL5vq/f
QTePWtGrpZsQVHRMrjduRNJjUjgIKWvZjq23MWgDrwUybNpV2snQzs1z4jUhBq6VBXqGj+k6rKUT
x5Awhe/zFjLZzOw+HTs3Fq9QsTAgDxZYRn08Nrl/mC4BWlQly64jxOh7HgCkQ/wkdSh6tn/0C1Lv
MPwUh1B466+8s3ZCeGHetOkuEgR0WWZlY3i51N5twZ7F+kShbu0LBnGze5qmxE/DkMUV+TT5hngf
BKtS5vDTrbdWr59Goi73Xr0xkcCde74QOmRCjlBwb1M64dheaH8+jmhRqdezBZd+depyl36S9IGL
Uu7YX1Ct7+lVXRkfPMQaCPyOjdLFDeZQHSBOTa60unjB+UqnSv7cuN53/NIJIfMkSHW5jekHlVGe
UcoBZ37JTFBbh4cG6UvyH7T+dA0bz/bPIVl4Njut23cbHjr0Seyz8dE6/YvKsntAVj6KM3QVFEVu
k5EXmBSz4ioik1rAkRkrMoH5CenU7KDcFvMZtlzJfqHes7QPdMG3qIAn05Y3V86aeZ+oWDJPogO4
5Sd7VTWiz31aDyD+xrThSMdqk7+YdaRrdkDuoAmvhr0oRU6Xfhrm4cEZIlyzjozPM7qbvpMcS4Ko
XOCfEXwsN3lalYffQ/G809eYbucDBTsnswmtlaJe6c68CQlGjnEsJljPpb7u8zY8UWKsa+s4rrO4
EzprpI+BJnWcqQrAThXVm4vh40lKw9mvmCLtascQ0/Yw7K+A6YcnB8XEh125S+OLjwa/j1VbkgAt
aEBzrmA0+3TbomibN51ZMU1FVzCD/uyqNRV3j505Mj0A81957gAJrPDiFN3C1Joo/BPq4Sqh0d/m
Y1KbiLB3n5wmJJlFDZIwjy/fGd9z/TS8ag18Bbdqb02bgNFA/MuRuR82RiIX0rr3Z6Pxwr6g01Bh
tudOBDBi5rYZsKYkcRdadypoQEcFRS81q38FApne0a8jFDflhhJRrnbe8aZjSvCTORIKiPhAataW
RW4iYX13ccK/hX14881rhRKYuCQTk6Fo/kHFDp+azoBFpYKz7JfCmikoFp3k+DwVDXZ1cBPkbExO
FZDK61GVCcXWVtYug7LCU3HP5SvZlbULKQbEhLZKWK9TQDmlE674aTMhflgo77o59ZbYaafk6NfC
IMnbjDpOYnmlB/CCWBVqPgUG/nIDDO+JCWK47Nvm13yLoXr5DqkIqA2dTasqA8dg0FJH7lKH9eaI
PpWJafxe1z5qjBGuX+ATW1bJZUmJm0MfKLV+ML6Bkvv0/Trmsn3bbWNegPjWxh354gZcE/MvmyVu
vCSD1vqhK+m4JGGs3ll8/OxIdxQICO5OoeFmtceC532onc312O7kxHjdU3+CjerVdublLYCmIeLj
fq2/EmxS1NinxuwUrt8JsI/AYUeS3ZV4straspy7PVblryeqy7rOgoiAoIcfKFcuSP8KzIM9+xNP
cXnloVJt9liPxyFqjnvRu4yb6KJrCyMPhL6zikyNr2iSbuj2fkBvxG78K6yy6O84ePo5al2oKhrV
p3D5Ps6gsG8EMCDiQWUpI2mA54ptM7+/vfkeRqnpbzc8n3Yh9vO2iQI1cTsebilg9+PFegPAIWrz
M+ezWxubC/hXmy4lpdOMQWkIiqp6JBN1DH3UqSKwq7LAMRFCahrJ+vPKpr6jtuoP2Fs/67rSpLPL
Iv12Or3FfM3lWEJI5SRTMr7FKav7k3oq5H1GiSidsJHlaIZJMASvEdgSe0BuFpGwEIJdXM73+Lfx
DVEeLC47MoFzk4OqhEJkvWs4LGR7O/bx5ShYejPezMq/NYz4m5XwDFD1uphYGlMJOE15zXFQPHRe
CdCleYORcaLGK+OR4dndOAEmSfd/Y/m6B23KULBDtdOg5vUV80IPfrenoDziLgJ85p1pIwFl3L5Z
EvyHU1NY5/9pTYs8QBFbxwEtySarIhe26dt/8oxmNc9zULWGbZLP+wk/A8ihbTzukGo1RPG+UYf9
duDVURHi5WVTfbwpPR8r9zwhfvNEpz2DfFFT2AWeVV8jEa/AIZaGHadpht1rqPu9Y67Nh6Gqfla5
Cl6O0Eh6FkEC0H0eGyoje6g9KpCx0k6mFVydmKPNwao+41jzFGw6bkWfiBGevR3zIJyWAX4zgobS
nOwAMzI+kJMWhGZOfbagENRHKxrq9cn25WK8GZ62tEi6/5MTQXcswHJFgopnbA4cBUAM236M383i
siSfNMs48LZXBXjsmV3V3bi4CLLZGFw3vQrBSx2XuVzLo4FbKFdzCghkteaNGZKQ8rvPxxZQenAW
Nuj6DT1kwWDqjbFHBVwKUEQqB765NSB2w+8w9VsI1qQbe6gXsv+GZ7sM5nf6I6yC/MgUiEjYRE5G
Tj2imZKFG4Td21d4YPgmJBIbC6Y4Lwja+gFSqUnZnUlkeu0PQZX0m5AZ3qEnAqQvy1c71nFcCpZN
ssGULsxSI3pjle/fHtsXx8QKKFuqwsGB8oxK0rEDoRmw5+4RNr24weREz/+gntT+gFfkjuL/dqS4
7Wh4XVuXq3BRfL/LQFkucRG/XGeXacsMtcGoMQC5Y9uSKGSsD8sdxT0KdV0Bojt+j/4qmzkGq6sR
voQFewbpsJ3s1HdxUgYyvLml6Ge8k9raZwz4xeDum5tCio1mXIrEwwVd49kk0NRI1rvjpceSTz66
Htj5rkp+C4cbPlWrI/Is+rW2/dEpRHQItGttcOhr+oPOVBgofmycRmmKfe3PHpMK71iMwk3x0ZbY
Z1Ed6LPaHZpXXOuklYvwFCp0ZbYJqbSfo3cJvkfS6/Uxx4IAywr4SoLhcB+LE1eobIP4NC2YKhmn
BKSJagJmIrZV9OHEW3Z/WIBTdPan3fcHd/NRzgy8ZKnUOSQ91zjekswgnJ2N6MHB8qZLjaAhArtm
vKH8Pgj9xeHmOiJvjbFDaqC+V3Gsp2bsuzNFsgOGPxGQZvLCGV0LQD/yMSVq/yFoyQsLFqD27/BX
KtTZQghqx6YWdkYTNmEFV8vCVoYAXqbhqYaCH9AqBjY/JdAwLN7t5X3GNeIV5NUADT4TETXxh7IY
VHmZy2rya5Cg0YF0/OvS9o/+69WAyqejEF6rMxDVRdN4hIbnBdmlAM/s+Pi2iLUOITC55/DU+bNX
HyiOYvytNP/hNjpv9u3hz/dHzQzhuTB7s4M1/6FF7aVR97ELh//n/SLuP8rhz6xtGWR2YbU2rlVu
JfAvW7JgSdK77vH4/Zi17ldPix2HUKeOnNt7Qeo0LDfESHjKnwJclXiXBnOq2kDiL7fqoEfOoHrn
nhZbR1Lji1fdhYKl4EfF1rO9YGZ46tYpZWa9FV3sA2F86o0zRG3vJZCdpgwBmES28Cm/5Y8NocNW
bERwhaSlVgjyRTVBnFGNFz6ttaLWR0nfITrExa3G5skwq75O9mJbwn8rBTb2LKOB9vAWrFrv/Roc
dTkhTrBQ6VUewXqqow4f3qZQr7GNOLRSqFYmCC+yODKC8O00mnHhHJQTsJJXA2TS6BeuJhO0RXEN
HCgi0AZXPdAqblKnIxcWlD/Afr1hdSf9shsN9h9IdQyVoLrE2exgt7mXNEegvCGkKgGSodJOnLHZ
qNAazYET/LClndOiU/qMiCf/T9NZsd5uXD/Haip20Q/cEDpmKmI4YyrNR/S9u/+A6jiBr34i2QLL
JSEsVp9aq2PcYDuN/rYBKNqZF/IZD13klvNF+05TyIiZFRMNklHLGElguEjKPuuxwlKTXcMglLvI
A1lQ+2AchNvAcg6a9xYZfqivwgAhLe+ZqINTC/T8BV+1bjKWZdR8gdv8pnvdpPsyF17zDwopeg+y
YHq1+z0/UwyJn8J90ThSMTInC0N49v6fXoBfTn1hTyTsk21GuknqwfsjMRxVUo0CQ9TuT9VDEuQ/
Nh7BtfgAopokj7ifVnVmrr+ar50RRPEDcI9VyAJFrkpmjYGz1Lk5cmfNDZu9E2CTpf9PEAQE2VmN
nWnSt1Qufd67rKhoH6ujqCwB23eBDzalgkyWEF1uEKlSMRXn4VwtJgOVw+WQNTa6fzNIGiH1/eUV
7W9FenSjWxeuEnGRzNRLi2lmYnDJJansCBw5hELY4lbCEOv1acEvL+xNTGFX177smDP6DxtaavTV
XVCEEdrYGmKd86XVvBk1ddIP6Djp4bN1stTWSOhWIvbRgx7JvLScupSYymFd3uuIbstYP6+s2Vvj
3gtJ0JMKF4ePta6XXS/FFEBzApj+en1DNtIHi73WFBfIPk15NJM0wik1mCd5gxigoMi1Y12y/LZF
f1ajUTOOLNQ0cJ7QWDSQiXuSPsGAcz+3YgPmt3mJNb4RUDqNnWphYFJkWRsXHXc0zUxlLD2RiqKH
YKyOqnkmkvQlIhbKWUGpo2+vVFiKNGp0WK19bMTcpav1IyQ/vpvGQIQlAQw3v43a/pTbl2ymSnwk
FdxOFdt9CjTzayqPAURMbeC52y3mkGya7Ax5boj3YMbYDzinsgOa67nnD5maedNni1zF56n/qa9T
87B4TIbbGZbI9rQEGu2WfomE42ZdiS6peC8c8D1alagT1DaFr+REt1+aW4wNF0fl0+E8xsro6tkE
Egr3C805zBahz3OccvYXiYZl3YfQa+EXpKvYF6PFGA80XW1JPmdw9F+q30Gz6vCTKVXkRMWgj3wZ
2o3ysSoGD5QLWCdV3KzoFGFMBT5v1+QfZG+LM3ClgLssxfK2W0hDmAtbFCfiLQtc2wd7DtbbkUVf
I6bwqlqd+3u0CACUYtXDlVK++y6V2//vR/nJ0Pm8Tb9+wiAINV7If+/VgnFv54kSl7E/I5T4uNxW
QTtr+rZKqmwKo7pxCRrJkRZezV9k61JK+pEUfPdy11LrmBSeDAnfWfM8XGXcN60DAo/eLn3dPm5J
ZnCV7RNo+PwDQNJchXduFi6c7eooK2CRhYda86ezTygoRrZVaap1LdrsTplSpmB1F+rKVqxAPWpH
R4sqJjApX+QYrGHcNiXQvjh2AupcMqHQZ3pphhGoRxej7xOFRdxIJPTgsu+CjmFQXK16/Srv3EyJ
mRwtgEayKQHJXHU6yv6Gk9irW/KlsHzg3RU3pKLz/BVDmCxT/nOMBGlhgw3b1bZiWH0LFnWV0ZNK
5YnY7gIPsVZugn55O/NjRQnUL54IxU914FD9+OoiFGrf4Ndm9WpupUdvW56uD1yLvFHgA3hqqfEC
mZCJHCsIIccPvOYpy8xyOJA2apzD20An61UydZSOMh611AemrY2PKVmn+gxG1FlRr9aSWKWhu3+E
ci2GJwXKkXzaGlkgUO/PC7XKZGvpq/7Mcel1zjJ4ki3sfLcwH3iUeXJ2och3KsMUTB1+O7242Sbn
+EJo0hwRRwraqY5XusB7zBIRIbMjddGrgzMKUYyJrM1iMQqLKGfMW2gYnTpNFxcNfMJu62AB/s8s
Af1Z87WW80wmcPI/RelOyM5EyHX9dTQEf8ZCBacGawCzdxSfkb1xA7VMb7fmFwUXLBHvfhAY71c/
dV5tEw3h072GHi7iiw6lWpzAi580H9vJjw7IKtQlrP0wAHyzZewN1JVihAL63BKtYoz6ITuiQ6aI
gu6yvfrG7A/nguwpafXeu9m6nK5PUc2Clgi7fP2Z3WorRqLotkevOFarvgR5PJ6kQjxaa0Y/5GPW
fD5llq3u4NI+U2Z26BMqMNk5i8A/OQ0k2ITk75Ub8j5OUEf/2zvsc9p8O54NJGZSqZUimH3TBpBF
lsvRHxgWqJ6+wS3Glzyl49HsOgxL3JmDVvDuTdivYPTr9cL/OdOV1K8CR9/Ys2VP95pQa9NRwUhR
2nfc8aKjPz4AhqEJVGJlowKC2H2/C/8yAM7vA7sHMcvOvs8WswJ3fZwuwSECtnImv9Dr6gsWHoGo
E9CDhhP3xlVXCnxSilgpbB/vQfEcwOq5uqCLJIZgtHhyppX9eVqWt3Ql4m4M/RaMA3TWQJSK6jf3
uscvw9v4HQMnXfnB/S8nm7WaG8z7PJMYcXktBEyJRIto9fpd/NpmrtHIR4MOPP6RNdGtdsNxgqsG
1K0ljdMg7p4jnruGsMhdAK0TyystKIVR43+WmTn+4E4Log9i9gclj43BVaCNCBd8zYoHqVpdQfVl
VjHLLo4nqT/BCha9/wypMhI9Mg6FQXdNEbe8O/JsbQ6CX1KdwvutLpLMRWQrn51a/VpLYKFx5X8J
dP18iMi3GzvB09btXBEZpxAvp0JMAJoT7bGa9H7++1iQiuTNfWT2XTT9MSd5Umu9PY/wyyvspUw/
gLjLL4Vi3nEoAnjM7IVvNsril4CO/NJBKXRmiBWp4w+nrwJ8SvLbt8Jjd3pyOnINDVUlkj9Zw2go
WH3YQ8NbRUH0iQiZR2rl9FAO+IHH+kzntEQCcvQ6Vi7i2zKjO4YjntPYL7UK356gUSctQgSeFQiW
9+F9FXolTW8Ni8WRtZT+qcZOaKk6J3rniukm/Z5L6E34PTOphdCwS1HckfpL6/u07pwbjHERkSpi
kJqF9x0zsS7w7W8BHQLnpIH9ppsBHqHE7dbMKY7go6ZAa0dOKL0itEGx5OO3HMqoFcNke8AqU0BP
6Yt8IbPB2Xtns+C0HdoVxKiAeBFgN2EySNrxlwArjzbHjR1oAecHUUD6ORzJHBL6tiPIO5F0uyLa
3Rj4kvXSCASqkIi/vccYy0jl2q0T83Dy5lrABomYGlTEZDiYSCQ1nXzghAz0RW8B0fZNerwJNP6A
LJK0URhyH88SBO2Cu2KztuJKenAKyTO0023URRdVIIhxPYxo44WZaTmWh8eTRDZqleVWedi9rJdb
+56B/92x2Lt9q099eHHwrsKgc8BnMgm2T7idhw6BbAClMye+yrf9LyGkQMQl+O8p/1h2obuTXHV6
zwNFuBoh6KjovM+2Y8iCjtlo+b/CtWftvg9bsEBeyea+AvhVa/IIULGjnU5grvuUQxsuXqmxSIei
KoNr6/Hujgqq3IfqKTlsVILsgsvHBB43V+7dk3geBSKN6SYliHgcNlX6fpZ7qJEJPjv/lMqsfaPX
VzSkm+d0q8k9nixeWwHHz6wVZNl4UI5Vle9NTPz3uzZTo4UIMh7qeUOR5sO3i4ZbOdqBIjAjC9aK
Q5L0Fx+UpPTn7UlyyMUtNiQ8XLa7dunpREYtruQcTmQgXh08uZDhKcvyPK4XxVKiIcIGdJdXLQro
+MkDEjiCnR89gCrDp+Ls0FV9fSsUooKDgS/V/vYx21K7TIAX37YpumBr4XHwwuK0+/lmhO7TfdHh
3uOOisE6sOuLnZ9Ealh+nk2hn9E0UlFkcEYJqQrP22qn3wJ54BdpoIkV2RSl+tZw8GHnqGm+yn5Z
7WtT84cPoQY3MjBwicPcnB/FVK6wm7+y4uYtSE9bc02x/t+dUVHKVycXkL8At0hIvauiUUDAvYBc
T60dloxiDRErO1kOxZLwPPpUMsZ6tVcwu6VWmbgM1o0RQE7iLlpm9crbQK+m8K2jnH9RzhrBlP7/
hvLWWlj1d4+cViIm6gzNdBmUyRSdulVb+5B1Ys5+qSR1ByOwG3SHvDxyReKYo2NJ3RTySIrMh0vv
xHSeo41xS0sbgPaT3c3Wf0kQSdOY/sxHmtnIJTY/XhxOZ51f4FPaJtxNE/ZR7wRLNvh6CyTjkCRn
Ixx18j0pzzHJ+P28Gwz+sQD6EWQGIOhbmk3L54DkLRXM2fhvblozNCSabUghT84pv9B6XapE8RF7
U8fQQYXH5bAgx4qMJZpGqLvD+n5kZzXkcaGFtT6yHN0n+clx6p7OG3nq1Xt/Jp6/H8hnxdirDHTT
0JYjM/rV9JmGNaqkzNyOWn/WeS5iV8ilwYXDgHuypTewKsvl2vUJW7Yp4RlJNWtF3UaBEK4/TRym
y4pOSy+qoPTQifZlVC0oLUt/8GsR9zOfIDUkPSP92MFDHPi5GWWQ4XVTu0rXDeMNHt5E0eRekMwX
RflqyjX7EQ0oOI6d3OoD4uU29CWLv9EkELYgJIA59rA1FCLxRsBpwsf1fTsHXGj1BSdGDYK99iTZ
KX8GeaKMev++G++AyAxcVhmWHHK7YLgP11LYBlWbR9Yv4fSzRS4yZJDpN4GNe9la5S2fYUytELOL
CyY8KHSB5Egb4AEHdN4Sg6eTdqt05PFGEf7xyOpN2X9NzAAT60/GtrBRGo45fiWV3RSc+iBCqQFj
iDCHFaN/m8qtyWzJTeyaheUjJaETn3A23U35c+bRYuJoRar4j2i0bZBtUxFHIXpkztD6BZAiBDPx
X2l/7DDX3SU+v8SHwpA83wFgVd9QfgAk6w2NOscvamc6g8rJ5Udr+krUBj9hGj9P8qdoureXA7yT
EZPMhCsQryfKs2fUT0bUjMWoAXuL5qAuluOVpBHIEx4Od9FbbdejKZkNvewYVB97YUsShZ3By0CF
+AH7uxzjGwKFTD0kjga0TBy09ZqG7UHk1/xnfT1MjVzBUu7vxGGcXh+JlX6N2yBPCQS+9IUiYEen
xGaez1D/lYPOk+rnmp/uybzMHNea3MOsd+RWj0ztj/K69qAZ/8XUMBoOOKnUfONErKV9Nv7BoxQ6
TByHE9G8wDi2tjJIOwW1IlGOzgjPCoAUSD07nmJI2d4IAgS5HJLdhS5KcXHHbvm92Q45MUcm4vXa
K+15ch0ZSRE0TcglItZddj4QYlUowVCulD8KAqVQgDB1t1F+FBDOe2BhzhWTrBFs0DyziHoEwGUT
hNJzCeyvCz9OcWAj+Yu6tRJp6PuBvUfaIE3lpEGYpajsHvU9RcgH6b392Y7VW/YM8T5M1IhvhfrG
OtbFNyAB+PUWWIQuftD9DMobPFWMUtEJVnniXli82lKX1ElmAf7W9kF0xQeNp/uCUvDmpuwVmiSN
14GthEBF/Feuj2dDGEUKxODGRNavAoW4R9XAnu4dfYCrufRMAXW7d386b2mqsTi7QLy+PoMg74JU
Cpd4cCuiW/vvz1f2ftykJbQTgiuQcXxr5W1V0yTsg5sWQvrBzmMdNPlJViUTrjwb0g/PloT0UMEm
EoqrabxLU52CkTkDGKpxHxRvkTUms/W/9rIKNyoRGCVibRTxXR7SWN1d5KwrmwI+QSLDZBuZ/Jo6
4cVwsO0t352z7hu+mdnyiZItqxwcIQaeCpSeqagonFfdmE6g2T9sX5TeIeNLedl9qd7W831M9LjF
HKhD4JyNcv1AJMwPZNQ/di2ml3FK2xP7wag96I2h+Qu7/D0hSLXTbDt3MnDFDmRJiYZHl3DuABgP
oWSb8nW49qOiZ58M4uYzeorm8+nPmVHpMcC/l0jKqBAStTR92bCRlLD4XxAyYCe4v6Xp1WN39fWx
J4gEN2hD0pfMaP6LjB08BxSI8iRoUUCQQf3BXWSgKL6fS8cWwzINRxBFhf/83XEZUPe37pWG34u1
JUFsWPG5XJbUOuv83QbEc5pZI6Odzeez/wRRY03r2LzfF6O1mehytwzgP2qmcscTLuuH9RPKZnfq
oyiSXHOiUxi8NYIGrIRF54O8VVIras1VJZlqgfAOroDdArpvoGai9eVcNahBShPVI87UbM/YcDd+
12UwPgyimPsloO/FdIT0lXWcncldc5zel1S+8uIK6/6rTNjHObtTcGuCdR1tgnAlJrceI+DV1T8m
tfWtWlp6zJt7D7O3w+CCDGcNNpb5V6orU5if4XlOZYavxBJPPyotXq1ebL0j0UXoa9csSOcRD0eF
Z8F8OkkORqnMimO6jHJkU4Lgr+D/+MsBboCpunLse/kKW6zeaHSzPE7+HdLqFiFjUyRBW8OhMUxR
XaIXUEnxrd85Tatob5qePOi6Qw7y0fPc+uxTDWaGQaNmzBVbvZWuv6m8sK9/YFuBYEervGyD6AVO
2nLNUjX5TOJJFfdQbEintVhK8RBJapvgIYmApP6SGNP3cJRE+Yda7XdHlp05fvEUa3qdqnkJJGFx
VzX1uQGfsfAP3Tf1EV3CzT9pQrFm7iwegfYgaNm21PK6QU24k4bl4sZRifyeg8iaR2pPMC4/+khM
DHW3ZGQ+yIbvfuud5CW6hWqWQ0/tZGBXlhdNZQZdcf3BLVyTNDZvPjgpeMnVEfjgqz2t7xJyuiT7
bBhOqM2k95zpHMflJOFHfKL5OTod5LJohS8MFoUJCZ8J2Y92y2gavYLaJJ8YPkhly6OAITcre4uN
Snssekx950NZWmLhB7f1Jf1mfcb0X26wv7/ueQz+gQrRxsxuehkEghsUJIFcZ1uPZvB8BRk6kgRZ
q9pMmkBZpTr/SWcf8kANffm61VrRkVwTOen+mQpKvM8YvUBSmeqt1LaUKj0ajD1UQRMb7H6ArfRV
rjShIk0b123ctwYvRWsEDmI+ILlNkIKBR2pCa644JMt6hbjIXEFJbbjrRF6H6XN6YEiUotT027dW
z9uIe4iycP3dSK30OdIn/SWy4g5AlQjjcX/xnAyJWEdIsV613OuzEPzIYe80dfNXarN4UVpEvN2I
FIRBgRhmaF3UWz+q2G8HbOXvFMXygO0lXQIODnIXNdvqauIb96wNvT+bIrW5wPHws5jXLCYlUid9
DLqsjnb9z+JA5N8RR0Q9XvaNaCvI1Gz6p0zqHyKnyiRSTtnT1rqsiL9B+EQtHL+dUqkKrTM/shKp
7DRC94/qABD37Q9z1I8EMPHSnF6TyyF7AxNMJFXF6NXpmmFKxgM7o+V2yAtEGqEXgnSQUedcnaC3
yBdwOM6IxwoNfAy3NFFNkriytrqpsWCAZRScS2ZSu+8MRUt/wBbYNHda+iqgJLfvQ4B80lQN21l/
2aKptk9xsoEEhkw9HtgaPMeAzu+pC8WsB+ct3WvcXN4aWmSraYX806C/f791D6ijZiMhH42/ewX8
mR6vwS4kR1KmIGDwTNvRdyt5YalIwzvfp8QGZg2+v70uENJf//+J6QaF48fMT8tAfOqS3srgNLRG
0PZSUAdcyMueujdnk701dSpk5QSn9ycOpzaN60f3Dz8XtJMrRuxiK/seurX+M8z5FQK2TS7olChE
ErUgQGEGLr6oYJuFsSoNaE4IGiA7DMaC3lnc3XM8WJ1j/rj/5goN4qCwBUs6u5b7qfED0x5w1oBp
0oZacbS78sNd7zLquOWwSI5CdCOU9bsA597byIq5Zp0uS8LSa3nk59K51xWygthyDUEData1Fckq
v2HS6UYUw9SQDNwALt0wO2/UtBpLvmllqZe6H4w9vRu9VzVNr5Y85g5Oo07dNuyW/6g6xo2YsBF8
6nvrNRbdL10EarRvCegURHnAXEZnl08qagsWDBmccrnFKj2eyBK7J0uRu7jayQA+hQvGR0GRSiRv
rBWF1kptZi9uFgP14e4B7abR2EQBXDPnuWD+D3++9vpSGbmet28QSDo/Fdnxq2x8CvvyNqiz2tnA
dawGomPD/dpl8KdDRrbLYi8wVQJLqUqSrjMQ++NdtFFwwcoCEAhUJ2r0vY51RCo4SY36bFsKHU3o
KdRNwF4rdHNoPSVYr706518ciuNiUJVcfLcS7PUZc/8IkBpzQ2iqj4BpHQhpT65Ah8yGqSio/aYF
jTB7/blbGGNnlZnJ1aaUF9OHxkOqHdIayHvMgvaEoAMyjf+y/gr7/8u7Oszu3kXf3p/eLfBUn2Pb
YpgNpj8qpd7fX8gDCBz7TwpBxq/FkbMFENfwaA7Ulg6FnMSGB6eKLLHawUjR63tmVSC80ZCyKjz2
Wftd+NW1wLlZ3CUSc64Cu0T1LpRLx0zpsWc985ZtarN124VyF0EvGDOsNWd9hNw0N8Tm75Kjzcaa
/fEnm1c1wOMxl0LyG77fyRYIDsPgmZ6+g8VWUJa879cxmt/oVu/RUEelvHf4ke1lVIzCnjVbQbqg
sv8/APllqXzmQNRBmBQHPG/xn8VDLdRTBsr3ycKXgoo5y6K+t3PL+z1tO7MVbF/ixV8sUfclMWI8
3fbFvtaa/aoKqvSEAn+QfXOIAlKf7FVzvVtyYpjFvEJGx0RYcq0VR6PhsEeQkbpdY3fVcTbRGmPp
jA3jxgvge1xHZ/aAyT8rYahEJ+x5unu7LQgcjC+zXK+T26X94y/sDMmp1FF45AQWNCqKGAHmvRjM
O1OZ40aGZaVhoH8qTuO+PMcn2Qj6lNp5TE+mzVe88ZIlhnFU5w96/I1spah/2Fy+7soiPu1nqy64
CoPw3I2nh2a8hd6vycv21Uk/3vyhd+KM4HHaS4K7Y4C517MMg4Q8cI+UxgaO3UpX9T0S8GKzW6WX
e7EA8o8qzvVV2nNM56ia/4kTfGkS8pDqko1g0AD0SKv23iaEnfEwNiQ0g1YNtDIZTgMo83pdXXBn
YLHr9XU+Q6sF13zlQh7ranpiGZmX0Q+saLfRCQC2/lEcUlrTu4hdAm5zgn6Lr2FgD1Mtj2/OVlGt
As3/ta5zBbIn2Df3M+jcjrwHw9GZXmv6UzFmE//YNAsNAEcrYW+CAut2STVPdYZCYsa9hA6JItm6
eqG6DrGBa+uNKJ+Rhyt5CZ1Z9TzkdLLC9dmrlpihWLIY6b2+29WeR0mws6jnUCP4fl6qyAIugOjm
viEA9WYXpEsyN6NPj8eGwv7AJ/ELA4euq6wPvzTd7USW9IBDH9t2Lv04l+9n2F+pFbUpFIxmfU04
rA14Kj1SDOtBMXFKTCgyHN5JOAEVB470WEd89qPry9Ql6MsphQgr7VXn7NwpAYgNp3DxjEal14Sd
OJ9q7MrtUelA2Z6KS/0NiO6JjMzuvMUUkErj2mffp7Cs5pMsH2ffMsE4iEzFF3VBRvdBnJSRahiq
HE/+wyW/tnkneGH+Y5m7DHyWc/QrElw1Y2o1NXYkd+C55hW4ugD08bHElRGa49oQQ8/Ul9ZiK3yy
khgF0VpT79Req+EwZZLc4+dl1r9BC1WKA5PA5tAzpaNticsOwhmqHQv8r4t6q30riS3xlQCVnR/c
cu6aJ0bs28qc1eeEmyJtbFaDSyRj2wC/TQK3DztgApRJZutEgPylIbEM7WhjQ0gf+11fMdLgQdYe
P7u9ckC95/PYXOhF5Du6gtwY/xE4o6SCOJQ/LDZEb+xd17rquRvwnVwxMdMhN5FtikXTqRCns2Mw
V0nne8UIZv/+fgrmPAONI2b7EboUUB7LpXJeld6crbXNZgyt4ibMHap2ZmKrwtgmn5togxC407SJ
aa5eTf4qmb6f+CdLfVzKom/xJSx3wvtZ97nlkWK/cpPE+cI4RhhHR+7KD/OaHhsYKJTh19NdiQE8
jp1J95o0J29j4kMNm5OpMQVVsVn3aSHdLdaGx24IW4RkYVwXRxioRVjBp81eT2C7vGMqK0WwsClv
/uhNY66UAs6aedEMoSmufWhQ5lJvf9MGQbkk+6x6DDB7NtirqyRi2fT2JZKv02obbpk16MiR3Yj6
UbPaPhne5iiTug8TlQf5nQ3pfK4ceU1PX/q9prLXqG7IB2py0qQLSOSmfjiD1d4ftrGJQFiONQZ+
3b8g0SZSTSuzJJmuMkuyZSc1KiEMvGachGB6Od6EkdLXOMBvdtgGh1oQZq5Be5vtJq0Yy8jN8yOI
MwpuDqlmct9MwW9m4azIUxGzKem7sKez6OHWeQXi0fXS2rHEK0h0kXrUmfGLuncxuHaMc9G2XFBk
s4Joe+A2ftQrM2vpGUoeAYeTgHMwqJaCnwqWucCQNFve23stC6ISiGn5AuFteUIbdcyvs52Q034c
ENgEqMofLbsl5LyQDwq8D2pPXFjjy6mHjHAhI18ICNEmDT+HdbjGv8mwwVRCpPciwipK7vhU1eGg
ZNkIkq6awjKgoA0hfhaVqkG4WyiAu+AD5C/KzGWm98+BDeG0173/fepo9cyMTjp6TXmLeKm1oR+c
6e9RYb/6JK0ZOqjy8rw0N1Lrb32DXCyzJ28MAGaR1t+gb4+GWuIsZXtTKI08FY1WgM/hWfSdaksQ
mvtcY253IeaNh2MWpoxl7L49hklubgq20cmg8n9q0Sydy84h4iAG69uLpNvRBZfqFsVJhUrbxWyJ
aMJA3cFK/Aw8I79P6hhhxTGxn/koryDnB8Ht1+Rr6M2i/tiGkM36sNTIacUqyujEYOz+m1fWRRi9
NmKzXefzNJGZmBjX0TbfrXz8qsGwoI5WrxLE7TycceA7LlYNyz1qHEltKZbhJ6tkXMlmsC/xUGXl
rlic2+zdXwcvRYFiTWBLWAreK9LVZx1qUNMQaSiyPbAu30zfcUDspl72yGzGUgZ4TAgWdMkDUL1x
6hR7j/DQMvwYyBCwYV6UZdic6mGm2cmyCyKTUgQk0iauslnXB+0c4r/3M4+t24Y+I6Vm98vnySwA
37AKWjH+Ep2FFUTJ+ZtxaY6klf1bcMDYLT0qIfYMfRifahYBAC6IbRmGzavYrS7M/xhLvKErxWXa
wLlqPUz0fIKJTgqaoClJsSL5Kcg3pDlvvhBMpYOKaR3su9b6+fXTNHecP51dFO831SG/2+2Uob0W
cIybTzVfa2Kse6Hj6cP3pKbp196t0g/M+LmCSf4JTXmGpQtWNQlgjkEqT6GqjVnmyVnJBgs5EqTi
E509Jw+eEZgQg7HrW5FM9qAwcX0Xe2VVUXfvPy0UPHCdpSHpdlkiIHOCyHQUCxzrj+iWNuJCqLWc
m/JslgJyFm5THXeBwzCaNEvpGORptC4kD0yZcENQiSsx46cSLnmQPOxB+tTz9M10jHN3mQkndhPT
l3mATGzWeEE3/xGDNttBS0TT5pwr3VAo9o7+q+4+yUAsXCt/76VrqDtevIKQMmckRE26mHCzzAZS
mgrb0FP8DpWjfveOmsXVPqPeFRvjsQFclj0gIPwrecHuff91beIm+zi+FeQ2Qr9uWemGgyhhuN0R
sQjqRyGKBygLKbwmt0LIK2aTlQ3QS3YjvEoWGFhnYzbXPpkjaZlTlRvi8H6NsZyQGOHeALJXOBZn
9eZQXchc74WbscCuZKSfXf+/eWYDsJOkQGRH2VV9BlwsOLDb1qcMYrwl4XzLVkjy7NBdDHtQsfSO
cAFvsQUdN3LzBlHQL6OsNUXUNE9DZBU3yDXhGpyvFn1tbr1jYeqhU3sIeqZoGl/V1AcQOkqZ5hj1
DYNBMcfgzkcaJeH04Od0L6mPnS4f5t4Ag/uMvwv4WDQnDQM+01/UHpizqGAnFHAyxDk5pJ7XUg9t
G6BzF3tBx+PrKQ4eyu0YxAau+Ko/7sp0gm5L/uK0fNkcA4xrAG22SeYu77J+LSJNOtRh6ibOC1rX
w7DG1EeDi+6bkQHmrJ/vaEVfvQjQ4RMITDspgy1yz51iMzaG6NYL+RwNAU7OA7eByBdsDmWuCCvC
/LlSQbcuA722+A3wMnDXrkipNNY0rcU1u6Cz2QyOSmMXAq5SXZsOSm9M/4oAeUdpsMgurPrWcju+
67JnwKwtr3jdRPQlrsYS227Y3mTkk/+pKO0CnDSJ9r6JK9exy5wTmN9uKucpV63wQuhkilUn0WJo
M0RQYpN2IxqDzuRIM2HEFmCJbp7EIIgSAEGBlvvq/3SOHiCmBaLOmPp9taAGTVcS67fwEmpibkhF
Mwd527O4XdOBhGnQ5PkuMFa+ZrMen7PEt6TFjAoynNh7nW0UzxOJW1ld9YnBqPLlLLavaaB1vdo1
iYmHG9oUnKKJCQRDumXJ8xrWi7A+RRHZN7Yr2Kh5/HyZ3d+rVplCyIdxgzZk2qLhh6IUF7bqFbvm
EjoOVdyCOdCNMpV8cW50RYy8Fpr5khH4lSXrclXlxXSimSKrDXpl/pnBi5N0rDutT2LyicaYqAZn
0rcVmBo6vHPhN24QbfOGyHZhrprKB9dO6CnrrSsiG2sgNRvg31ghn46s7oari7oXkbm6FOzkax2U
pS7hMw5ts1z7diOFukoP191u4uCwqXZ9pso/BwggrZmXRsan3MwSKg5SuvPEKhO7mwOcBvxC2+Yu
wHaOQuFAGZTQHuABOhYngRCRXe6kGkyrHZ7jHobtlwOJ6f2LWzmyabDnQnWskJgo/vQbYb5oVCEc
SPLTWhzu1bqh/Ey64YH7EoyyFVOn6jsGVeoL4tqBe9M0rBHhzNWgZc07WoutXeppLQb1Dt2zrwIU
yHG+E3uk4pp2yJ7kNAznG3sFapgh/XxAFLM3niNHXAXro2CUDNgPF5YixHBXblv3rCQXSuXxfHA6
vxX8R12zltcorjUWeIvo6hnxYE7jR0LAwUWGtbqav+bcJDACjX5qfMZXwsHe/4KJOLTiDmArxm01
2wlqOPdK4CE75KIo9/sY6udJ5CgJfq1mkBrlcCE7cLStHVSwV1/52eB03kk8EzkLKhIhQLB5EmvN
8Rd0/SzCCCXnlkJqeUI4qYeiCQdqmrJ1WV6ixnxBd/6Yuxat36l6UvlAUl3dspCDUwwkS+CA0pTD
HJH2fB26/aGs78G3S6QdFHtL8a3PWznxivxtqdYScS8KmBChyxUUMF+MvyZPfIZ9cVz4cw7yVf74
dgTn2Si0WaPxYbwjquDLmN1GiV+ZnR2on2CD4g6J+4cqJgwNKveMG6yWYkys8Tpy6rCYSMk7zYef
aHiSKbKCQ4NXbjeszaWKYmVBwcEV07vTHkYKALq32HOHD0Fmjrb34LvWj/Yz9gt+zFcgm2TGwsIu
QIf7ncCR12YyNejyJJMXF17ZYXfw1l2SluApl4/wZP/6vPtXgCftIsldU6cNcKd9WJfoJd945NUC
32Yk4nRvQ7AzVQd+EIKEyyGscc1RG+glT8ogAZ8vdhxGE7H/aYfnPK9MlkQKEWixEtd9C7khENfo
bpoVohRok0yKN942876IZ6FSFCXFuURJ2tGB9GT6G/oYl2vRzOoHSi3MvCYJFjfBuUaXZ1SR/Lwd
jj0pocBBru1ddHCHuCPY3l8ljfTH9LasHds4Md2ivrZ4j0K9EfqtrdZTzABxvQK/u4b1AIm4fb+I
9LsTySuvBKXvrzQa2xCZbnDDsafJufZn1+ClBcu8U9EPXSKCdfrmLdXiVp5WPj9iTO0W9I+8LFKG
4+6K6OBCZ/Jw9bLLi2PbPRRkdbZ4mXW+CByPaVhB/ZvlzzICDAUUerYv9ssZveUpO/sxVgpfv5eR
Hw9xNvSRiXGxygr3LmBCB57BYEsUfsilEEBsV8M3zUDCEMVo9hmKwRpREvHcyB4YOFkjZCQZ5Stn
lH+oobic8N+g8EIhvI4IgqPDQOvvBWRNDSWYjEhibgXwVt8YCU+SajmULcM2pcDMTapvpHW4LgHg
swPkIs0OudIqdW2sJa6/TbLOfotbDHRGwbuvy/jPxqElVwTtCVojDhhtLdJqfMZi23yGiki/Zl9p
qCQ08OU5gVppDY0zV0IRvxRNU6ZMHNNUkJU902l/9tXCBpIGaZ04LHgnYGNFm0YZA+8g9BDq7FYj
QtyE2qrWyh6/HdlVgbhcHIYayO7yzZ45ErHpixstYSodlRmJvmqJZ/DKooRFpHfBnSvsl6Keyj7I
eUVvSkJzqP4dnjcaWrpGUETraTblFagTYQddKFv6JiF2UxiZjd60PtJ1FoNBzZNOyI5ta41VLqTu
Uu9UF5Rb62HB0B2gtPpZx6doH3eiVCBroOE1XRNP/jAr5qY7/ITAc5VERvd+daoc6pY0Bvk9G4Si
U238u4w0WfnuY3n9seVrvePAQiWeroNhULnMAL38nLG3zLJm95LADDPiI7da68qIlMua2MLDWMdF
Q42JRU/qBGHTqGR10wlJS9jLTlluATAUBlLYgY9fQDTNL4I4yOG1J49+CGu/gqVHPy2WbGxdcZ7I
MqjROBozx22UOVpCrguO1OpFTQIG8oKEUmUIp1H9JvjIiIxaqzuCL1nQDKml1/FnnSuhMIDn8RAE
M3kHOy64/lGCnpGBryLNBLUlDoBOCykGq2nqeIpikNEcDJ+4Xv3NYkVLSfAc2pDgdnTeMYRYo7II
h+lkeT2P1e/9QtcLEc58UJaAPx5a8UiX6+Hpx1/rdX30kt5FrU/NGkIxPb4fDeHw8E7q7hbpDdSo
Rtkv8Fa2x5mj0EjY9YKzNX0g7mg6qxXbAMGmlB7+fChqDvvUCWv8HAq/7v+A68K45ttpOwnkW8fT
LIdPCZXUhM5io9mIxIVKCEF8SUhuDPcKEcKZ28c2AjZHZy57IoH7fEHu/oYASPUq4dtDazEwEtuB
4tMqMKHCtpoSXdXgV27KCOzQPETxABEvg+XLncwDP3B0yCcF6kbnF8Vy+20o1HV600RuM0tTwwJV
WZ3zoVJ+yCB8jLqFCVTn+d1/JPpqu+PAEljfgDJwQsJ57Ai8nstdz+2/skcFO+G3euir8u4pY8Ns
5EI9TdHYPVZ4PPd3/qDH0ssDE4LzrLsoXNqs6a6W6yv+Vp/NCNqm9gZUxsWAli4ANrEcVuI6/MCI
bN5wWuS5T+eqNu7/Ui6/9W8kaDprQ/1oA6oLjixORu8/EC8s7/MCdk7jH68J2obRweo4UCcFC96d
ktVNTqA1dmUxuvBaClk8u+kwba4mlMsCbGit2lGrNK66XkXvcANQsxz11uwFB/DQfb+Am4a2oXn2
nuxOtM4lqKyAl8Ls2g4b7jSDi40X5KBx7ALlKEuiS3HoDVEFU7LczPvvZ6bZK8K5wTv/N4eoAsbJ
XXHN3kcMsKo4gMOd/T3yT0vYB3iyVFrZ06co3duIn6/tCgzITgANcBM4C0gTInngY038b20segC9
oYwjP6WvTYOskXdUeI/REiLvJ765S6kQAGHXZux8fB2YCFN+LsD6Yo7yEV6hLnGXzanZ93cQJU9b
AErNKppV4PU95rQmp1SCcVcp4+v7ebPqJKKh3okllKxG0quxhTMHhW0CC8ycqNOBbMaaLWnjnDSp
UMDH4brSBEG+ucVObQUgLEuqEfQ2esx1yQ/+JKixOKtE8RGwzEwexzzN3GVrK6Ran3kFh6VQX2y9
SsSu+LD2S8fY3qqPgGxAPUV6JICApxcGaxM5/eE5diAMX4v4vvRiev8Ftwz8GtQ+psCTawgmHV9u
TtuEc4XmSQkh7aQ3q2uIiXYfsrB6rmj7nKABXscsLJe6MKplZyCycvUUhILocAzcE4e8+Wo9ZACm
vfq2IHTFHcsOTyn1qaK4wRkgVZxwDbmJ2MJNpa/Ij5mGpOsGEe9rp5wOXQ3OSUshA25GB9E1sKhS
CZCN7UQK45vAHnfrFCrXxVp0pDQBiUWeYCN3PF0WPXCzsYt6MMeLQWj2yyn7KunHD5IEZCDdRbag
vLPOLg1zJwGzJFoH5C3P8T7GY9+wIfB80V2W3zi99c7p2Pqm/tOw+z3PYrGp2liTxIHoem7a6YIm
V5Qpzzq1xF4IAcUYRbJKZYZFdyFESnJVRgi99ONypRqZpItvzvacPKSzDUEu+2Ugj0uFynCkCNJd
m2Xz2drlbOZGKWXkWWq/1tfj/5B7oyIvgTHMZur4M5WGAtnOWPtBUOa0N/3nu/CL5/nDbsdVKD+M
YhiCOadA6TBKmzOjobpESz4jSBj0MtJbt07Xz3PipxKrZWTvS3qHMj/Ezm67TvQ+HeJfPdVLYD4o
GL9xPLGT+3ELDJdwsyhYYpcCb4Vj6JHph9+0ZyYS+zterNaVcmlJx2kKs1pVbuaWZ2UW/3rsmiPM
QU6Z9VNBIwnGnwF8JwmdKymw0RaJic94TMBQH62a7fkmi335a41A8lalHvuipJjhqphAzr2G2EsH
U9OZoX/F/xuE9rYwsQLnVWI+mSOlP6Qae5eVd5C+X10OK0eCiata2YCfcjHlGe5ZADKdf6+Ph5Ts
LsjYjcV/ngyyPmsDt2yxdtoJVPco5Zyr2lyBFFJq6ikLRZXluoPEnZdTYWrjst1l3m6Z+wE7mrAO
VTlTq7ptOW2D/JPSnLnEBRn64EDlvfrTVyVCYZPPX1mzwx/EW28FGE78TA1XfLVoTCbNf5s6HOWr
kdyeoCUl4Ye3XwtUcDKUQRfEFSo/qXTKzdwPrDzRDjQynZuLISoPeVhp9HWhJSefyafCDYb1I8Le
1M+RxK0Gs3AW+n7IfrSiwguDNLdWZVMn9s1akwmuopoF5lJ0EqtCinSUEH4zh9Te9grXS0cKNsJI
6CBJiRjmgaJNpdfQ4A3dGolWublDCr831Ayf5RUl8r2TZNUzgifJQfHjREsG0ukTn2znqBT2RJ3t
u81qJdvuCIQIoW3llG5t49oE+Iri7KNNckjP5laq4s4pVwSB9AjTwqOf+5tVT0YM30U0ycJLzU/u
n0vVPUGK1UVHKVuvHr9zHeY6wIaql4oUAy3ZygiFmPyvgnWeL4gqhd6K86n5vh8AhwETnQZb6dWF
HS4cZi7/QQNasAUExHNk8MEDiPMIAHJPhp0cVsOiW7iKCmUyE7r0+nxx0oD9bw+UchUKFs7jQvwg
IKEZP8wHEUZ4DOmTtSDfl0xab+85rnxX4p8Rsxq4xEnKPPDA1ahympPSNEbrlCW5l9ksnAKproCz
rzoBzwkp9zpNuIazCTtvn3N/fEEUWIucGTT4LzHBhQlIGx31uZC3IOZkWC4er5sQIh/ALv8AxrXY
+tXoKa3wOxybHhug2chGhZltHwcI7bGtW12xN0Nr+CPr77qLyTZAJUQ3FK5l90fgOrfB/udlMgFw
1bQ5C1NxYCK2pvtNzW5GqWPp0zrJkteMDkbc9Kb0p9Siwi6hPpf+C/DYYM5+c3mxt0Wn0QhKZPVi
t51U95GRcKndhehURuwoOS1ThMl+fj9W5JD1tf7p99lUgKSZywcucGw76B3neG4VDQVFpr/eRInp
JNLW5Xlk9SlveeDQCbH9z6i4JAg9PQAjbWFquvCl//2RgFungCGL54cFFXvMGhAwWWM0UdU0kfIN
ApBA4r79odDO6GT0Dkewdd1mZmU8T9nNE146yH08TKV8B+YBcWd0YU1SDWeLVecayS3NzX5wyM0O
7gTBGf6SO3FcN3FWjLTqq55XZIh+3uScnxElfChkBthdov/ueXY7/z8MDKeh9vkn0iMSxSGW4Oxu
2ZMfUAKYbGfG/3Lpkw5/oXCYaPxG8voAMhx2bWiCPWIR7V7SXypsp7LPlokATdqMnRDBL3HryjlD
lohVBqu6OvRQMPck2iNhm8maPFgt6ytdxp5qVw9/M5EFqGk14w8WMbPaHFsNkVJA/UUgTYxB+323
+HC/BhSnTGila7D3rc0a4ZeeTRaF35VeJlZcpH5V+qjhTJL4bFHffOZ9pxEaBMadMhvsfCix+UjH
RxvVSnI5MqKfFmEaAd0ImwtcfnMM7hzJNDkcMYisOPIfCTf3jBbMVsRPK3XU2HncwGP/MrxP8tQU
QiYuUD9ODzjMzjeFcMT7XML8ZMdRj8QboWgbyoJUtyK81hPmkl/FaD/ePnkEjQw6Quq9wSSFnY58
KlE+3rjWhVQwpDBtzoHBgogzQStPCWGMvqeRHY2rY9n2mtbRDijOgAJMNVGyNCLObn/XwGC87F1L
SESCJYY8m/yq+5VC8yu4nc4hKt5RsVvjHALUIjGw55douOXh5PdCtsLdI4YWInSlgJlMFy9Hcrpc
SofEhQlLDMWWIIQQvMVA8ZhqBJzMmkqPqOmSBgGRzy5i3ZVhbnDFeW6FlCrSu2a/NlmNX5Se4xDK
6crK6kwud26X6Bfu9I5kBvEXSRK9rpOd9fXFpFh2nnjvItjcw2ZhjZEcxhfNZ6GQXqQM22Kccv7+
DA0RTEaFulTYmSvjCStBjMS0gfaXV6LlDAvoH3pHfnzDmI/D6XgDtf8DdkvCIlv5oeO+wCoPqk1+
9A1LxBCTmLfl/OT0H5Ea1okWSQtsScGok6fj006NiGEGfloIGlrgN3mCuPjJgeNOmmJKL1E1lyzq
z/g9sb5r21e53srbhsZz5omOwAl8F7jBfn1RTr4+uaVvftjZQ5B255f81U+YNG/sMfUXukwZvoBy
H2Sz2Uw5pEnONVwJBrUhb/yThOMSOSjaM3ptl/A6eTaOTXjhMb6zFnVd9VG9VzKw2xWgCR5cD2r0
Gr+i0yGJMAjRM7df59X6yAxHCVyxiWvkpqdKUS2o2d81gh+h7Ocb+ARcmj8YDFNm7GuKC33xnYs8
8jI3LaepPeTuZr7s9U+Oa+bjK8+3bt8ltGM3U5OhiQ9j6FHCtkroSukb874aHl1Kayw69lJqZGY8
dnQaFta71Ed0OYFfps7bq1KQ0GG5uXse8qIDPAvnL5ltHlhIo4mWQBwYDnFolczvl8Y8CPEgsoTU
QV5o9p8ndPvBjTpTQoc1uzXVtL+pc3BtMDTRYKVQfznXt5ooBwCalPlQYCz44srkf5EipTOVA4xA
jG8HuQEjr2D7hbiu3xCpX+7uOJ+I85utu+RDp+qoQmMghDOI+QUCC5ncBSh8mrHF99yWXRgU7zUI
BUplHouJJil2SxEk0R4kTjS8Fntk+hsjuU+U03pRF5iFilWN3sSeUMqKWrTfnXFixB3JREiIp19w
0V+GX3vI7vL9bbs6byc6cEzr9g9zGfMrGOT7poKnuRUdjOLo1oE7Dp7alGjUFJiD7NGHU07FeCod
v+gZGo820e1PMO0fb2QIc7O2GNUYb8sg7rZmoHidz48kgR4Qp+8FGfo1BGcD3z9yiyR3MhAWc7ZG
HjybbiX9ghYs81pkz1FLurBteQscorOzvREfj42kJ0ubWANmNRrDMp3ECNbfq4Xzv8cMPmtbfSQx
efOqCBieH+eNC1vH+Thyno7a+JS14XDpqf+6UQ8m8yOVjsNJiVLix2VHHd0fpwKZCbv1Vtz957x4
SqmwW6PIh7Kq77HAibWAxYZi9cgKxhzOCK5wOKDZUIoUhVB3D7nF0S9CM9/sSDBpujgRASbTH+dk
GjndXpvye0XhRBPhW2qcvDvWG6/Dc5e0gZgTlui2yBTbyCMQHjHRv7pSBMoX5HnS+RiVPfWzSa3O
haG5XUOR8bhuvNMDNCPQTRINXiSdcPjti6boXp24TGh5f7eqh8kHV+Urch2kFGGV/wp16IPvPQxN
olua0XmfJbpDhiLZMdzZgt5DxojMoYbwyzdx34JEMIXfad3TQaey6bnAPwilLB8GkyBatBKnPVUi
g57gZ3sjOvQVAHcc1HmIkyRktZgMTLfunyQX+9zxLwLvwAVWO0pKizx7QKSf9s7La/Y7Qi2/VFAY
0kqxk7Pjr+NHvq7I7MO08vBu+bt9Q062D6ekoQlley9Tw+fSKFFrl+vQrg1Q3vtQbmG9SxwU0F/E
9rgDnu65e2mRWWjQuXmsyX2HQ03DZ9raT/Aac3LrscsT+PydEDvAX+kDf65R3OeKkoeOh+XvRQ46
QJw8bOpUcwmwTqikIUmh/hgbCWZAgpEKhYcwva/SkPhgRJnfOTaQQdBMj8vntbUn95mxTxlG/NL/
ZNOV0jVDxlbrVBNwqgo6OEkDe5N1+hW75lhmt0jZtLniDMxuXiPckCMsbEicsm4iih8g/l28kJma
nMzR+KiS5ZLcQzq0zsTUcwJp8TS6WrOdSMTOaG3gTIk241KttsqH9K9wwktNWt7gm3wtin2n9Ey1
ukeWAnhPbc/2py+Ve3M7Ip5ELVaU9zB/0SKyTJv6mQvpWh5CQJoWRsQiDThRFq+ERIyj/+NKZIVs
ncWjN+QHmmei29gm4Lt8SHa4Bx+tL4zyfCzxdnCGJFcIkLBWLGorI8h/iaGgXMXpUjNWDOuza20C
psHDManRa5qIf4vuCy/9hM0ziK5tjaXPC5pbC7+vMj0G2nmPA28BjcLHhAErWbF2pIA8oVEnME1s
SNOruyhAmfyVYIT4u1qg5C6eQyv29Pu3jaskHY61zoVMOz1Mvp7CLTd6t8Bm/TgzLCUmcFJeonKX
+qKAmBEEbVpSI/K6neqodzU0K9VuZ1QzXIoXMZb+6/Cgwb8goUjfiSUbxnr8+GOEhm/krGzM+IO1
KNX1cc++HlQI3cQdtBWLxWgyLPNY0zE/YtO0yZhc1YIcbtO3U8bUgEJJtk5hRDRLoXK8XqQUSicI
edbUfDDdo3XbKmhXUjXnisIjPIICrIh4KTO0euMof2+cwzw22ifXUqmm8M+xepZGAroHYbum4HFW
mAAFtyX/cYT8jFxHpIOHu90nf7HeVf7f7vseUYF4W5Jk4A8YL8daavDUxOYUrb8i9n7zckc2z1wH
9lAQmrdsMsx/i1z0guCGHKWtVvKp/G15joBH63H9X6YvooQWbRIo/NvpVxlyAFYFdiA4FeUx9D91
H+r0ZR9pC70ezl8gLJU2ezMpnvXdKUKYsc+/iaTsMbgTqgO1ac7gcDH/hJJubR6xHlZdoPZarMge
mGRO5LMib8b3JTry3u1XNYpfDkW6+Qp5ZAwneJFb2gPity5Ke3aPHN3AysxFZBMXQFyes9Pzb4KN
n3xdP/rV7lpzYH3Jry1KUFANGEod3y1mhAMcJrWan50y+upXdY/1n+JpUR8Bo5rtPpeWBvbVCYfr
eaWKsqzP1uTELNqzsykkdfiQPlAAOETv28FwBVQPPIIqTywldjBuwFbZJQHINxdk+eTqM5BOqAST
48QQBM0znB+l+2TddTlNAPdZx/QwALSBvjQea7rc4JvmDHbf4xI8ziNdb+ZSmPxkSwdgWE/XbWpF
Ncbg8YMULqmaXjIMxtiJcFzf6P45f+71Ey4o0u8tE7w+c1xwdBYinIEZGwtJs9P0C7AOLHGDw932
qwlrv2hvnxNbZQtFKKBi09ClAwUAsWrHqZxDDSgQ4d07MD8BOa/3OWHSqx/euxEGZii8Po/0j9Ty
oEqtJpxEH8e0YeOzDLx39dqUAQpHFcjssXC+19ISGii14kfuEKtXfvcgWy7570wOo/4oszDR06zC
+oaxCc9wq4+aTZZyFEyI5eEtRaiJ7/eW0xAHZSfq1n1e/aJkoWmsBEZwSTgn0I9j9HO86s4ncCvF
D6ovPOn/lwmcCIXy5MvLCv0DO+Mb6ZSuyPP5Wh32rAAWVnMEk3wdDSC9VeWK+tZ+qjCaZO4WdUse
6dt+PGOhZstYduqqfKnHXLvvq2jBDeD/h75IGnTeelhQnc+Ui2BthMhb6x+eZ5au3H1lyRbI8SDw
iXogUCxZUhTjF/MLvAwS7qcpzSh7WIp6dnq0bChV2V8OPHQYIqyfzAjTYItRL8oA/3aCYu1lw+QC
uQNkkqnrpRLK5M4NECSas/I51vvshJ994kr9UgPi2NsxlaJB1QreJALXROEdMZhdDQjD1yLEgvAU
xSu44aUkQ8W3qhX+iysNRVGy8lQhGfssCoaczLYUYZsrc5JCTdtH94gJ4KA7Xvi084m1Al/uH+t6
aC++84zFsOo7n4dH+d828yBdpSaUHsMUL6kDOiI7spOsiW8mWe8L5S3RVJgnmWN9/5Z3/HZYC7e5
QyaYLMzbI/Irov392+kHnVOwOBFp6RDzXB63DfhMnrAV8ieZgELKF1k4gTue8t6/5WIY+opEuzkP
vA31v/O68fgoIRN0kyIurd0Ga+Hy9/OgwKLOO19loWx5Hg0OkD36JLbVrya8M9s301BhU8N+7e9C
tFDqY3nvnx6OIAF6xKbT5Uh2pyNX3QcfpiDy8/qWejbzx2THDBl2rvPXkTvV/2Lq0tUlg0cuBP+3
adsxe6Z4qL0SEPsmEgpN9b7se5yGHS7q3A3XR8KoT+wkojDGwppBsF3WouzWUyfBnll+BxVQIDas
a9oWPhKsKOkSHxYeX/MBsoYzVhkQyeQZKKG+9ETgFrMjqIpkm3bQEO7vnkOISw3LlSQztLlvkxCM
rUS4Lvyi2Qhg7s51ipS7k0VXtq8MUymZhR6jrFJJsu8J+a6avRSurKL7hJTEEMTSHJUqJkice50d
ATF5Zd68xK3c7elkGKM4KZU+or92jRLjIg6bjJuABq3T7pyy+xmrRk8TnFuTJw7rRDP1G23jnJde
cmtIns2AddCOgCxCkug/42fyexq2VdJO+nttsf/PeDu2JeWSF0Wia2xnt1B3+28mcEzUBP2EvtU1
Vq/fk2VPduJNkSTXBHx0bmYJ4qJU7mCYcRrFk95R8+teIkqUnBDASRnN8U90ZWo2izntCHnPHtEQ
8iV+iWtq8qZpQkSeU4BEJlD4hlym3xapVoYFVG5sckKWp1hlTl9rRBD7Kn0aITAMEQI0l80imW+P
wxCDEgpgVGFnI4Z1qx2WUbiEeAq1xfPWKokOnvd6kklubySxP+Sam57D38Mz7TnOpv2+PmHfhdKG
GvGfC0g8JF2e7ZgEsYgViX0HhfOyZ/DgsP6x6fzV9RrBGD3HhVpF9salOB1RN+0TCbq9h1AMg70R
dLwFaW7HWaKMI8CkKvezZSbtGj3/3NRPGBaKK7SxqSyJwM6xJ9FAjCEGzS1+m5FCidoatF5Egt4j
3FTDBqyLlSODctylQXgH6D8A9eV3R9dqEBDu18HgWXY96AYeIqAZwtYJUVynxfI1wNvIfyA0y3P/
tY18UPW03HbB0gjDU8HFk1ILt/PsshPQMyhp/lWiovf5swFrPIq2fFMa85fB9T8oULNBUzQu1OPB
/xN/cweWskydj8xqPnL2bEJFSdv5AIPmbgqDpPoe2CbqYyjPqlXDe84jh/nVAPAhAn1Deu/JhlA2
hhqj63ai+99SMowZM7lOiLRO769W31i/Qxh8QbUidHdqiNLlLDEKhXerkc4dJJemlkMfLDlyb215
H1QAl38zQA8qCdshsx6alyTxvtbMpaUTAbMrDJzI0vupOU2kvwVjqbvca6fF9QKtDyCXredXi3zU
VV/qkgN/JHTrlDpQTcgAU1nHMhJrv2A+3upJvxb6cpzJk+V1HI78ZbMhv1GwHq5B7qUM59OjS02l
ajY6ns6Zaanwp9xVXduLuyKNUzPNekTVNnRhx7+yN4vjgGJAovo9kWwlS7m8xZi1rjBCJSHPwCYW
fk8mQZcZRd+0XahyXu+Ugl2mnhr8Lzt+1xbgQZ7E9YZaachZ36lVCc6oxDPwNy2OOKrbMXBi1B1g
gs9xgvEY2HDdadgOqcmkvMh/2WcWN4OQUk7e4NLzzaLkMVOd5XzVioh5VzDV5I5PKoeVv6XgNW+b
OXUnXAODecm+OM4hAE52qIACeHCkSDsblsxl0kXPuUmd6Co2L95jfWX7d92esYpL/kL5XjuZGe41
u3GcqqzEZM/E1e6zBIyrGx7rI4egVccQxrLS+BlZ0c7bcd82qJ05HPHDK6BJtzA2uT3L9i0nPxSV
QaZr+9B2GSPsGVkn86IQicEaEi97ZyJsOOain0I+DZf5Pug5gpPazX9fPl93KvmNBI3bET76jGZW
7YwhI3FqGrknM5FSapoL/hwCXZwlro3aPJJEHchbPcMIOtyGdKFdhHu/QEupCJxuJLbipJYAbVVN
Xg9cC+Nyrerhhq/30U/1BQ1aGvdKqgUO+wfkVgl/NvVCnYh4ExokPeukh09teVcfNT5R54WksG4h
lLDQymz4kxSMxrvHzihdH59UtRRMGSEtEhm+lZd50xRPwlSjsE3LvT241S46gNXBdvtxsbdiM8+t
3JUezMvsxd9yyGJKTPUp5gHjkkKA76rmeOgTIPbNSvX0nNqH9jGnWl3MHxsGcPo7AscGsJRZ2wwb
GJUoO84Y6nROChRrNGqEdPg7NQBmQnD/JUY/wwBJ0cVwuu7TXjs74x59xWkktNpVbNR/NW0JGaSN
xB2oV9VEXlBSOQ276C8a76s09uzcJkQOyG7T1h2xCroXfFLNo8uZfQleQel4uc9vWfC+UUf41qaA
vfZH7aAcqJDfg04wghqyj03ko6n2k/4YMtjnlUWgsYAPOFZNKm2ScNGzNR2JfcdDKjssUu9hy1Jo
6cCm6ypdCNlLYj+rDxynRFr3x4YHr+Q+vQ5swR9f2DX0bXCcsMpFcn/5ds9Zsu5kODvZkC5PTI4W
f481iZwXfXzA/hfe2gUv7ythLducExIXwXLVWUUDNP3b0RHwCaWmIbMDuULgGZiYbuec8ljFQyGH
s1pAkjfqMld5UwKBINvIRYNH1MrGQYGDplCfnHhbWKsh+M1tIMevdM7uLKBZZyGM8y1kB/8wBE+m
ZVha2OzCkeOydTfNnKOizffK8yNJsz8jtHSluejwtt48+DEHHPCqwF11Ab4lDuumFRFLqR2warWW
W+k5y0+zBPI/nSta9SChffU91ILPRTE3K6qd6ybsFH7TV9O/M9gpsI/bnScisTR+I4CQiiLShitU
C8K8cel+qBI2/jiHSysrujhdtwzlWsGhsSlDzQ9G7KxPo2Ougq/IiTtrK/Ie+gSCI8yRGNy2DLNG
m60eCBjBDDmBfvTfR7/9j6BJrNk+Jv/OgMvYjnLfYpf4DSn2xtctyON4tPX/1sNE1wbbczQIh7qQ
ax0GxT2oajUKXktVa/ug1AiAhd78rOOCfbDYmWtKrqFcEDEU6QbvYFBbS67npWQ/qROtVmSWMls6
sqAt6r0j9PIZOqPtRLSQUE6cDiRL8DFNtEKGavpJ4SgkvR94DPS3d6lncqJ6Ptu52SNSf0Xkalsm
VeDANRNU0D/DlZ7ROalptgBJB1nueglYLUdbDLtnHl1ntNnLP5aBti3tnEF51W331pX11Mxlo1OH
K5oqYIUSolF6HWGixIQjaTrDmYZkKZRuWparyp2EaIMqmoBcwxzvq+zcgVhPf+i+hX5W0BHn0NKF
WCzIe5o/aR7FekfC+mS55efvuEF0yTlDfW3FanICoTQeXda3abQMwnOzlKLMKAzjeA8NJmDeWBdq
Er+b9/YgYMyUsfcU7qqWE/+BbSUrIoFNVKVFKJrNdoRyHoENIHqTf3rDHahr+3r2NGtinGLmJ7Fe
y60jVe8ZpHbFeaH/Tx4WZRE9tTwetxVzp+/bZWZZOZdgJOzTa8g+4VFfL7DNtrG4ySqJxm6dm/27
04Q0QdhazFrD8LyGqarbfLhXVR1zodXRTgtpeHg18NTkyq4iezo/JMUZldWs0eftA55Hx+tz976B
2fHaHHK9KAsOGDKT3oQFUxKrw3IlH5gn2kICF9KamOcAaNuD4zqpLtKgCuGD1m9IVcfTIw2bMxFx
xqDZtgLM+4D3xd3Q9gJ3jtR4pN/TVHCKiAgQrGFfTq1BAqTvX14oLJB3POzAMEpT35CC6/Vl4cBV
XeLEYhAp7omEfS8up7xdmfJwHPLeLXnGxcv6M6/aLxGn3xDzkgBlptU0Lica/14rrS9j4LetAFGQ
l+JOISc2txItf71kQO5GKuV4bRRgfa0fp7zUSEOjR7m4xQUinOqSZwvbEEbL4UtkI6g5R89N//XI
0eAOhYxOCDBughkKDH8N4of4ZjxzC7TPiFMwiXhazGP+OUm5phhqkZ0Wp3CoRFuAlqTEDAQQBeE6
NNH7U0tj28wYhL4oUsxm2uK00msslWq8OgkbSEot/Qx7paoCtv/J9p6Fmw4aaL1yMm/CcBSXwxQT
P8gLz1nhrSuieKDYVjT4kz3hHGUlbqXL2GCPr//Rk1A0qPYhyRHgGjZxjdYqMwNqG9WD0TXKQ8XC
e2SUhuL+GW7jZmCURJefHh0Ak7UD1Db0BIRoLhh0zYnsVNwcLzsL1yDgHf0xnIp7V6FlOt8B6Ol9
iGf2A4voT5NBtC8ePeYsL987MZf2chpoSe8ULl0AgEV67zgbpUW8nnSKSZD50oQwnqwc7rtNRR9d
H0VlpQ6XKC24W1EHQtVygVxbZB67ZoDECFnAgcL/tebyXdVJinbC0QdiLvKGZhVKbyqu10SSL7ni
yVp6XSr5kAmJExLHqHkV6IJB1MFbuyx+qH7rFUCpsLWuMBEUaH6yti8NBCLgsrks4l+q6GfyJZuT
3OZgEQCOc3GbftbqMlCC7am+jSJXM2rC+hq6hROTmwdrGNsyMFMC9D61jo4pnQ673abX/iV74lhU
m7eR55o/CWYDHHoYX43lTa405I/codrFk8O1BRl5nWtWCus/7MBrOUvIze80lHKS6GGB3ux6Sx3a
S91eVUlmrqviJ3HmB1VYAjj8BIhjY2OEOp6Bq/fgwbY52TxRRfJkvmkplQfw8IdZeEMMp8+m5Al1
YdTk7UTrlTd3fcB6h5laSW2o2IQD0kOfb83KsopWEDrxDRHTIqC+hEM41Ou2DKv1pdYXy/16v/r7
HuuAXD5Gm18bgknEHu1dg53jMDX5pqqxXSyhbHN54ltx2hp4RdXPZetQoWzn/LD8dJbd06y/FPAZ
wDGCSNNI/fjKOltQtal5Sm9ROd+wlltrtijpN3CcGGzEINH9k56asOZXDCfABXR3tC2TFavCwLOZ
cSv0EGAXMyE/kRxSRU/njoUnIL5sWivF/5/3Q9PtgWCnDsikL460iDJnT0dgE4wjUZZbpXqwFhwk
x0S8JvYp/8p13+c/Cjq0Pn25dWGj4lNwB8ISvvyw09yGeW79F1iIjmnCflB6yhKts6i+sCcO6xio
EcEUKMtaz3sovTe/kIF//02EpOlNzfpse8RI0B/M844pRD7LxQRv9m9HYfeCZZfFY+uB3gVkhxfs
36txWKPNz0JL82Pf2/wlgUu2yHbpDwpgmHuxZQIpSSopgSjlix8MjlH51CCZfJef9I4mnPCS86E/
imCAr06oqIwHPkWBidQACNmFjDE43FpEjmJwJhcXWK1u7VOQPjtivcdxQ9wtE23gJQW7y1JJ/Ei3
BaX7V85pOjbdALEm7wcNSLCIbO7JEmNrD8ONXrDY3pmUqmbPM3S9+53u1ko6eXPyWFbAsy9mrdwD
ltD4O+HrkmstRhaNIrVbDcpxOsHmb8JyU7FOIH/iFKPdmB/M6p/MB1eXNReqtepGlbivNFUTD5MB
T70y4t71A+/aZ8ipOdbaPVP/o0M/yaCSVIulXqdPKC8W4a6d/G/+SVeqCYhd792b2t1CkrnYOHwa
qpnBsYKPyUAfZBLhjhkebt+iLYew3S3+0LtR2olykpmdZk0mVq0wa4B6GmQlxJ+Sra3ctxY/n2FS
097Vz2JUBBnap+TP9EG9/AHOFzTNnbU2oVphfmRYrew+y1HLSuj8fQswaV/qAguNy9WxRZ7cQB+i
9B8VCVeK5l1dRfP3Ocqllc5orXuh37nc8JmFc9wZ4NcPZgXmxvS7Bj/yfR1hf4SoYqIIwFd9CzGU
zwa9zcuc5EeQmqqP8063CAI7tMHArtYJlPt6jViGbC47AnXxWLY00pLmQwInyIFPmG30xleD7CaN
gKzsU5az27mXvbqTIQoxspip9rPT0OIc8mWIhKRejSomnZmDenfkRGmTrxFjs2JNbOZqc6QGvSYE
OhIWmbMBJ3LrIU09a+VzK0Hd+qTWvLaTOuHAPJu+TMUE/n29pY0hu+rvWipmtggPfvMLR/fX9lGo
REKLlIFLblWzDASmt+fKhbsY6w7Ea3Z1EOp1s2rKOjiQQW3zXbbxwewPRbckGNDbf21YoGvxVpEz
7Ffgc/jyEivMBeJt+gJiYseNmpRlBRDgVNGZPjY9oThKZVWiMVAD7yOC8O/1v4ezDqoTsCxy0H4d
F1/CNTBwAkv61aKhZI4v8czxxayVlq9Xpl64TThrtTyebHEAgwrZdel/x0J2q/J46AS44ARjxXw5
h4VFEqb1AKo1DINrXdhh6xQGh1CrYxSBmc0BMPd90dIoTV8dkXTfD5jBaYbbvccdwnmEOdPAFc8s
9sE5rWK7boSjyz/AUBOKKS4yAMRI0P7dCvj63BKllb933SM/lX1DG7/y8PI/BoW3iPqvei9NE5Cf
DuPlZpAiK/nknj54li3ZC/XA/p8sKME0FyfHKOmRnkGzfZSBkmg6gcJbmWXoCWxPH8DKyRTDZs/M
oDjQPlrBhglSJXzczWVQW2zf5OeM96a9zyvriFAMML1jpdVShYYckPsaWQISB8OSsU5/oP1Q8tlx
R46j4uFRtFbWb9fdFd/+grOE/lAS3SjwAJkavpz8AP0o8JSNEOEHoqkIWBb/pWLtGyjVTua59puF
70OpVE9pYbbV55Sdrqb/awq6/sJ7bAj4oGOu8egSrIrznnXouC2SEGf4+DFiQNHTMrzvlE75pCDX
no8vJvoNVCq9Dn4ghBNs2JM92wUUJC/Cgmzs3ASj52kJ6fdoDaQDI6li/inqQmQZ7MktcJtNUsEw
5zEESgOq6kNzfZViH8p+BHUergBuhYSefRJPSc8Z9EAlT8sfrFIT+1/NXMJugRY5516AInESFZGh
CtBNj0/2aMS4RikAH2tmvoCudq216TpZJfyNLT5hxySLNQjX77WaxGdXgV05mQGE76aeaqJ9jMzg
W5ujZCA4MsDb5vNPJxHPluXhBbJTQuYbE2nBitDZzXnrzuJoKuu01vSiA8M4QpdTEPpXzkx6llWl
se/ULmsgQtqmS5q+v0wQcsmyorctuPSURC4v9KtMrRhkZofqrp2+lM2grM76OTQTQGHB+5tX9s2G
pKcKnwrjo1Fvwm38OBGMU1/klBFRqLTE3qXb0JWn1rP5VSP/IJd6lLBJurhdyP8up6BX1BTifyJp
fBhkvJrkt+HbU7LyGcnOy5W0YA/2xflVP1Rk33KKSlyiYh9qLcTZJgIeaD8UgdH4FNe1+k23r7C+
UE8uBsu5TfmnhinFaKeKeQN1QLZo9Ql1rAvTm8r4pQcKIDIrjLedAvGgrk2FvrZbRZQRx/Q50Xj5
LlhfHeoNH0UicAImrT0MWXtyJyZ8+bMmUMCSyubErNHYfIux4Aol8QFoixchA//q8MBAmSgXyCHw
YI+chQNjtHnjj3xbP0rcHUOFu/drpOswNF8QfFcw/YOVlv7KWLKrHoXCh6H0Jnr7k4v84e5aYkwF
Fn/4dcnCjwvNpSKl/QdRSC52RDGKxckXekXUS3Ydw9wmmz8nrHwbdMw4s3dzWYiFp9FQnTpnw4NX
XUoOLX3ecMDzeHEWwqJZgdgVp5rrcgTx1CnKGYuma9otU46wErFFnkalI5x7hEmauaa6Aa2Xk+sN
tpiEkKmxZp1bX7Oet9/PzT3fda+Hq8Rxt7A9u96akQj00JkyTQaXKZl+KMQ+OmOlWawslikApKim
b+fDQm2iM9jRR4wxrI76Tx/G3CvQt82rTsUJ04Drav6m3mwWhiK+DjwoOGzZ4LSW7LnhyuulBxdy
AnucLoIAKK9ByTEC6xrZ/9rU1kkmRbZln5PArGxE0Ey4X8CE76J2ThUSZuvnREAXDIS+zWQLufba
iP5HtiCC51Naxn/5IVtzXzw95gzwYWSZl230AH8Ptx80t6fPbu3juAZul6MagNUz1jc/dhvLBeNf
DltQhXa2F4VQbuvUIasJ9DDRHnII5V3IF6zPmnwRmzTtevs2uBVYbbCTfSFchcgOyv7OSwlj6gEg
kSGJpKDnWttIdPnybiLUgpk4HG+CZ1qZlo6yo4r1JovMZnE2k4QUMq+14Lt5wsEMm0jnhzEVzqUp
091pibA8riGzd5VBNvZb7gUZ8kY4XnuW5WI350J3RFKDSGlBuNCbP/SbrGHy1fPiTvUxXd00QhXo
bfK2b8ywYtKTK0XQ8W97yOE3TLKdkQU/5NBmferVGKNbI2hOcRgDIXCMgXoD8hhKT/OScuQrg5Fe
3R1DdfGKlU749mpqGsnouc16P77icKn06xl1A1KyRg90it4QGLq3AuGKZo7lM1x57gkEljW/kjYG
Bdoc92SE6uijnalQm9vPvhfQx5CENI8SKViY0xXBHI9SD4hmmPTGWxPKWkDtXgsBfZKPiGadZRZ2
dsZQBa1AlQ/4MMMgxp8g0YyGdcFYuodzvboUSV+Iz4D2qCoNBsoIZaGt08IPjBBNTzffeUZ4SIz4
Om3NHAqv/uXebi9jI0M7y3DlnEzWXhI6RIlvD7xoL0P9Tywym1RjeIvtPpel1knzkKZTnpCmr3Wg
13ArtHfe+om0R6Oro3BKHUv+ma2XDeWGrstnMMK2abcduvlq0JImnRE9reVfynnUYZEND78xeGoK
2LV86JPDAtxilFuLCLondalFsauI2TksHVBdQFNU1Eq2akSwlxoFAzoXaaKrlPIh6MtF3r8BCxa2
ILvp/mhl1NGoMOp9eWeEPLFr4aNzT0TeMglmZ+n4TIMX/RLfZDf03LsFh600gNS59vjP3lK/4zbX
J0n0jfUCIJfRKlTDfkV91f8ZPpK9cTjQ8prtdKs7ik9BqGlCfIPnk071Id2nEcDeimaul3CarQXY
s7vj1XkeHQQQkOoKEZTzQX+bbY11YvXRU8i5LgoWALnM1HrFaxXtwEc/QoN7SpXBUn24rfpa39/b
SYv+T3k9hWq8QYs8Uakq2GMKGMbyMjmwH2XPi3TqhkpCjm2FvcK94kWb/D2idGiuQ3Ku3KVtgiSS
cUkBOdnSaz7JaIMbaNBoGqz4BhiJZ591MjPXps4Dv1us5ackvtkZJLpy2SNGGFskKrYQb8H7xm0Y
QwTX3+TCFlcEnKEMkUAtlAtFkbQmoFaKfJXq55u9yuLe2EEpYGISvX9SSbjxoBK02OadsZKvnx7M
JQjEELmWCl8OAAkemeYHveJS7q98VHUxUIbM+OQ+vBk0k3V9iY4+rBJNB0qQDA9HkFNg0K8aR83R
A8MJTGuq3TUb5coYct1lrpicsl+Gx3LhQXXYmV99FLeReO/v/NDZDwpOsi5XtIPC4+pRzomT4ZIE
oq0bLQ/pNxqRpuEFivaH1XgE1ZanDn/HQWDi+u7zVvr233WWhUQhbD650anBzUX0lGHhkxlaJdiY
Q0DSmATRz2/9jAuJdOj4lF+hkYGgDVRDonulnXrIt54DFRMp6mb8OhkVDJ7ko5a509I4qQksoFqO
ZtrxbvIWPWoDrzfGv+XxUlfo3+SsbqD00eCrATl1GJ3Odw6tnfC+91HBxdsGOBfJ20Zduim/Kn7t
oqUq86opGvOcmC6gjNjfczoR6kipmNQGt2BjFZqaIuVZjbHG5M0ndRkIuJ05gQm8y+bSzUGHIaLo
KTSSChRgh1v1Nw3UMU+ZmUG09b1q6nrDTx9X6R01fFKRW4/iuaKEntfWtM9QlPAOPmdzihxTrNFX
3pxOfsFxZuYE+6g5N0LC6qxOc2REUGtTOu8nKr+httgTpdK0tDw24j6WxyiHnUvV5MS93dSWxR8D
BSU33qnFiyuUyDIMFTrmFdUmVsd0rUaJu63zjripHSHIGrewHCh2ut50vD6FS6IoUtgDk+V40lkp
E7rJbg2yv2aDsFWuN+X1LAhKJaiVdXJXEIS6lNu1NOmUrP88D61w+pt0OUzM/FPYIdnp6w2Zx+C1
ywoaVawpc9cCqpZfwEQA7uZMpA+vdpC0GtRunBrlCWwNHPFA0Xrx1zqCNSs5zc/o3D63upnPL65U
74N0W48x3tBtZrr0KV6vFBwhpzMRGDkKywrHcDI+ED1UYkzV7ux+aAp06k5p3PBX8AuSatYCxmr2
p9DtqqRttn8mFSn2sdOOxxAlZWTHX/BKd4an+92Tl3dOe2KfaAwgoQ0cXgQ3zXc18ui1K42KSiJT
6sfJ1dhUYE518lDkW24g3rWWA8FgwLjNOfOxLth9gwMg4YcxUDp/VvzGr3Z+qTYiIlLAw8rV0vCG
w72ox5P90JMwAsakGeNrn3IqZq16lz21MoP8X6ZfwpxfBHzdWfPgYS2VuFyqS/D3hMlDDFcb47Kh
PX9KefFUAgxEH3wEzuVPDUB3rCIw7ZUPT1W25ZTkG6H7wu9GKl7arUyDzGQ18t/k0AEGT658P+pp
l421uV+DA11sAyLkXyzXOcJawzfNQXkhvV4Q6MDHklOuJLKlDFGTr38LDh6MiEgbTiCpEg8v2OUc
yU3Trt9UdxzsoWBCWhzWueV6GsZVjarnuo4wDQIhm7h4HmIQzx9kUy0skEQCYIJJTxIrtYS8z/7X
EqA7o7ISZMtYxYFS47UkQbVImcdI3LKSCr3JYZgX+3yySDRuxPx5zLTqGX4HxW6Tf4b68bfIwhDh
ShunRNUIgx/KboT3kThTF+6ibc4MXN5M22+jINxfNMmg4WJfIkyRsRRob0Xag241deo2WlafV4IH
+Dy4m4NLF2eVdGsbqRlJLjlNLCwv/h4ffOI4O9ep5lS7Ftc5Km7MS79AAOK+4bKagfkjfhuyecEz
qV2ZKe+BKZbl0+mqCO1L0XyEsAWCO+qTrym3KkYzB8e/stN/X/gq+Q9tRU/2mIfIYC9d0gA7RpKU
HOHqoO7/mtE0wJTn11w4AkVNmOg/lcfM6oUTTn+4QjoxZe7EiHKLeEDkhCvb4HT+hObloBXEf9rG
DbbCi8QKTcUsGar30kSAcKIxV2KOilIDRcHFinoO+d9NieiXtlT+pK2TfN6kjAu4OwG4jpc8s3xr
ll71ZlrxEKCqZLlweob/GedjKSudtDY0++bRc8EFixZUBPKsq1ZjqSjGhqZb9rK+ZoBNLebyM469
U+WlWLrs+RQpmV/s9InXMBsiTsqBaRLbTf08sFSKfLe58PvsyTOHlfe3PRSYla5xrwoSVmk4xI2X
Og2/bCrSRI/cgjYlYJHqaNJ4CSsRPeGV3NIM7JxaMeptGMcOQdCQgjJ3+dCoOR/xBDpAB23vMxF6
fp0DlKfbPYVrlsFFcWAc8CPA3+gZCoA2oK5SW+i4XAT3bp7INXEXzRHAAh81Gv7+CZb1QcOlLtqC
cos8cZCKEtw2dqzTwiK+Lskz0fGvCnf4f+AAw5SknkxgJ0BXAraiYMg36t4QzpN98O8qbSISCYAH
VjLmVKInf6qaPSre7gvCCmIReKr4O8pD5uofP707sgVdeZPv95c1V1Y3GaycG2s8sQYm5v18/FKA
feX4+LKon44/PQsMufD7QA2kgLkkCre7jnUArdA6FX2tRTacdVbU4KiUep/ImAttiAzXnHctqAhg
nbYlYPga2U3rT2l+09rLFQTSJxhUVTXoFnsKSsWOTO3qrhtKhdmpihCTu/roS5TKT7rjojs9Yd/x
B5OZd+gPK3l1d+2qjWxd9pW2KE5dA9FF5tVZVJoVy6VpG17I22aBqegicg3XrZHt14dNHW0dtOzv
JRtA0/98yKGw9Dhc77mvdJ2I01PxWskxCKe1Lb1lbHt+tZ+um2u8ASq99F7gHkpqVj2mamSqGSIS
AfsFBMiElDuk/zZGy6q3ecwV+0TIWgWCufXy8ZNfeESB7u95wJpLclwHcNebvQDOwpZx85gk+riJ
EOkS9L74nSrAMxxn91A77avslQarIe1cihvwcyCiI5aHDAr6Ucm9/wsqaaDqJV7JofNf0otRlcNU
CYVLMnfhN8uEee0Gytu7mvuUIUdhjvH5AvlJ0LiMwqVWNKS1MIdsv3DZ+NhU1CXpTZAYkYf7cSPF
TTS9/ftGkV6qoSaSKefE+ww6FBU9YdVt/d494/0LdP4By+SAN2IadWoNFWPgfrnKl+3nnMJt8QIC
eHIri+o8myFcrU6vMLPywZLbRJ+dzyWGx72q5JaKLvOB8yolj/B323UbiYLJRxJbAlhmfWSWIDJp
3Ts0C3LhfVEX//km39Gdm25h19nt0Bd+LmX5Lfy6vUYcdUUHlzvnk3MqW/v/UI7CaqiBt+1PFgeC
ZSnYs9oyMFyDpzz8FC6P3AO6+QBmXEcDMvNEManzuGCnsYUp3vDGR0L9dyU+ZKoaozy/CLRRUapi
hW0A9amE8O5C45r4qR9pGmdhZ2loYRPL35DHVBYKtjl6LFhV49td2XnjrKEP6qolOwuzw/QUBUeX
Pl0l/47gajZHR4zOHUOwYICQkX+6jqcd6fuHInTpr+AwTjLkzcksxgR4CReUsi+F8tVuq82yl5eR
N6Q409FYlMMfXzKWWnfmkxDSDNqvhJJ14kXak+FJ4m9PRmefXdr2x2DXBrUHmfPIlB0ZbmJxF7mK
QctmFSZDwRr6c9xGO3EU+f4Sw1ibplsiEPKH9x7Ve476Vlvtx7VcS+7bMLDrrbHo12t/M2E8c2J3
82AwI92d7/GbSLhMzu66so1q0LNwb18E9ccStbfZQkcESbjFF8QrXy1G0pwSH9O8I/ibjojvKvxl
VcEkJ5PkZFTX3WxnzGqnOiq9Flj4MqklI7Bo0zJcwyxKDxO6mpNLNERVkdffC05fP0ke7QfqtGym
AfrK1y5zFHZVjXJDpBmZ4f0FHblftoRf1fmEFebidEyH8KXc/OyweZJq8cHaxyBfhS9z006gdcfa
PNIrvSguvxSMnjntAfISD0xA2MNJ5LxnbM+HvOmS7zDnCt7OogYeTd+InOb0mmorzlKr5b9x967e
DQTB84IzkJYhNUWnpu3+leON3G7yJGk6ex9M3pbLG2FMQDh07FTwzcrgW17ATXehSApGwz2lwx7+
J28R9mDKZJjHtRytlWviEuwbh8i+koClrCv7eMXY1YOlqi+P1nCgwbMSTiq5qPdRw9alQnX8CXAu
upBj2ZFof5Ie9gfulcnq2iTOc82JJWebkFW40TBCVdLFvlY+US2fJt/4LzXinqJIKzufSudRkK0K
Jh2Uo7InBFkEMN4Tm8qtu/9NLTbJYYCDlnSxgSpTzFbcBE3lAznMcT1jFR4wrHucaLLfETHs0FAP
TDdf/QbI6vheulRpkINRcVF+8YgXdWus1OlAsHkBZ3Fwo2AM2IOLKj7eAbA6YOwzq7v15wioh4i3
cRFhkW/+iUb4ouklaKkzlieelYX7AwV+RV7rl1oxxWnwZPbwI9JKDFBiEF4AosXOitR/wyt6EL72
LJNwas52Aa8zmJN9D8QnNz2I5FPEi36i/8lb+xQVkJkzFt+0Qep6/zDAipwtARgzPTCUaHQHhrOR
jVr1YAk4wDoxmg0oPweSd6rg5Z4nHA59HEevfiGD4U5pt9F/NR+VeOxbcYM73uVJ6erzp3gr50G5
dEYLcp97rJ/BO1kcQB+cU8gYhip4vs5jB5th1PbVJ/8w2g9BNWvKluXw3TFVhXRbYRFsKKR5EuUr
DUmbO4xs60zxN2+uUDilznthF1LI2uyIrXZNiBrRgNfa78F3rCb21fyprwPo5AKjHbPDu4PkbjRv
uOfRt3hLT4lwllCdgfWGjvD7EfYs8yw2lnSyLE2d3iZ7hLRKpxOkT/uEMO+maaPEyrI4TM8gVigJ
do2C5IsH558eIOfWqkGgCouqOhToBM3df6zAL73Yd3cRziL9qRSVpRgp8spBMwfuHTWgRN4iovtw
9TMZdQitCml3lDJ9M4A3QEAe3kBdcpmNca453wVQybR/R2EqaARIooOkn907TGoKUmR588JU9rYw
eeyalM0tHZtMsrT1W90WVRiHEy+U/1mEcSvsNPkCGasXsXweQNu14HNxNqD1BIMa1UtIv2MsXIxc
fAgWQtw/vyRdxyPc81wSIqC74Y5vAq6URhcXEXiRTrqxYVmESRmKU1PzVIcuQZ3u9yUYto9cOmtj
i/XYziyqv9iqMD7zaP4rPk35gAIo1V9Q7K4VyvOozcruY+dww3IQjIH74IL1+T21wGe2i1dnRUCS
Rf7cDKWk+Qe0A7qINygahOAHXgwEQnTAlz/Oi0scJ1EkTMB1KhmRDU0cqPXHQS///YFW2PURyd7L
Ydkezahxbnu14gpZM06dYoSGqbNSFSaaGB7IO6/LSwvXVObarR4ZkhnnJGxotrJ0Gg35Oa3UIT2y
9ZhEVz2WvWokAl29mRV7F6jCdIJ3a5J9nJ1Zx5BLRYIKXcYCH8QMgw9dSKiAAi6sOmLT2+ZqVQjF
R0xEGiUH3RzppZM0q06PmuW+nvJ1uF5TNhBqcYQZn16WOMsUqCqOJACJCKDGjkazKc44gKVSKt1T
0+BNAedeFLi5n9RkqM/hKPJYu7FbfzoZOXzyEmb9OSUl9e3uzdMopZ2BjihiWtX0+a/nRM4lneRD
Vvfd20ph7d9HDC3oa8QARfTbgg9gIgVuhGzmRIM+q3Khx1BYY8ek0CY+NC1uaNWEz5+fh6auQ04A
C6jHCMLVShX7zD3XwcCM3+tyzsBmw1DihD8/hX1R9QQy4ztUiWffcQti8UnrDE4LDOuOnpqO17Y9
z0JnmRsQJD+OujTDymePUzntB80H2il/aCh8As51h1p/qcakeCR8GnjvLIZOgiYqBrFA/f6xnz59
cBGP2RDoFFd9dCQMnK1XTeB8O66weoOItxNoDkGM9/gegWEvrzgTLYX8llKq3tJvLX01fVe4mbsZ
hLs4N4AR0VtozGSjUg87ZX6zkCSwDMGZSUuzWxJX8oX5vbAyVNIHPYaUobrWmpCYWpxUQHQSsvnS
2o5vtvTV+1ASF6SGRjXvRVJJO3jXzML+Qxn5qgsl5HAkIVyecQdpaZ5gUqH4v9o/edl3jp7UDeEq
kdNwY7QD+8JgQnGBrtwQZ1iJfCcpCJCHVkcxPLZlRx39CNP2u24X9bJJt4YYGnCTWe8/XO+qW/Ut
HvPEEgv8nzASY/IJbRxMLtmUdQjfGvt9COmb0BIbv/RWq+qCv2eGyAUvxQE/m9MxdN2hHoHX6ogX
RybG7SbLM5BrL6lM6ROerNNO4BHcB/AxGJhU6X/p/5QvQ8Fl9glk4oUcfwZJ19cfdPLQ8EPE9NiG
qTihKsL0KaGbgrQl2HhB5NUXl3oH1V0jxaIuWnacsjj98NmvOt3jNA5P1iZInW+vMefR04KCSsWB
nOBa6pPzKRsXtzw9ljpNvNKrIhdGQFeUzOLv7ECpaYtSEuLo+v1XAdUoAilt24if6GNAnfhZ+oCT
BNzBvyWIQwBQfiUg/32jsU4Jj3Fmq8X6AhU0OF6UvcAZzMHc0X8tK9S1spvcuAE+bMhAr8vM71TL
s39VviamvBNuJLdFTmqoctu4Qt+5dyOm319+Vnx41QjDm6xgxpJdnje6RcBu9HuZB0+qzyz6yyk/
pxiCwKVZKTZ+5uhiuqP4DgWUAbX1ntbTT0l+6Pkx8Bl1/A7ydsSXLTtbmO12X91Bsi+2cCdsIA62
IgwjsW6IPxY5nlIlCVcs/xzSt5vM8eMRJrBSPAUjEwtOdN6gmrxHe/2m413Tut4XxxX0In5Brb5B
acblvyiY04IYCAJr9c82QhiWmaW4YdLl/Fq/Y6HHtGJDWAvc6oOFxGCFuFvAvQjXqBd+BEcjZz7W
3Ua9RvNGo8ZZ/t0vlGLPIaqM2QDepZJr+Rpawfo/0b0FrzUwOQLkPlmMdsHy58eWDdP/orXYLH+n
bdA1Hnevs2dqNT26bkEhIIcCTUxbfnqEw+B0uBnLRzGPTNUrbS4rTl2tcsfSj67q5C3sPsKNpLw7
s51GTtB0V2Xb0pOXjbBUdtNDgVSy4hTX1+5SSjwFq+YzdaqNKJ5PLK2BlcVXpg7viIkzRhT5FPWU
jDG2172vPXr+gvrShK3V0nxspQnepuyBBriBqjTMFHJguwBSizacKgVeCQ6QNWYdNPo4RvBtfqus
xVjn7Dtbgf5pdvXHandrLYhfIYhypzhst2hoSMY8URk/S0MKB+QSWPUjEiAPFZ21HDcs8vkQrvzt
33c6XDoJuhW0yn4/Vm3QDPlFJ+CT7p1E8zpCeT0BI7XbJQCJAa2onkqtMinot9ySGx/4B8zqCNoR
i4i18e0rfFVLvFblyLakMF6XNGn7CHzaKyMpaJXYDtOqzIT2wEN8pgZpd+MmTECTBtMIhh9LLQrW
0YVFY6/HQWguoPAQsrzvjXMCg+gJJ0Q5zAtKVdBGmgLUcC+KZj9Y4ADFuaeSh21RzElwLWX3G9Oq
+YNJ7yLKsasvxC9zTl+VVLohTLSMwEqHE71PqXnT0hqfK9HsYX8Aq4XhHtqOgaGwSaRrP+ZKzDXr
i7pKJsITN1+9d2lgR+tMcaplIH1hr3kX6fZ9ofWZRqsjlGe0OtPrq2ei611uIGwiDBDhm/OflBTq
VJY/n0JdVmFEc+QhB9LF0FgafiC1xPu13YNS6jN5v3ZZANeemSsIZJN66jrsBfcRIq9MgHx4QGI6
3dXPeRh8UZV90DernQYPoelS+WG88MsbpttxmryjV+RHiK0xKpUtT5Fqs0IKSsT2GelbhD66bbhI
SBulXssxILPJ1cmaFMd60ToP8OCvPlVRo9KbbApjMPib3uvMIiGGiyCn/IwnlYgH4boDhxTSBpHq
ZKxqJXw/aKfLPPfDHMGhF69f/dJee2COLmrb71uVctku13qMH3J0vUAOJD2KmuNRLmNlvP7PQSxH
7Ve2+DqidQr5UmVH0W394emF8Fw/S1YMtIxrAJriCAy5VaNpEJLRhb6k9/Xxsk4LrQBS8Dzj2egE
5pAr51UZqkHtnU3shxE3Ai5Lux5x86DMHyl5CH7uKOkwiwyYdTFEU4+EKDAkVnTjKHAIFu9enfgW
2EUFqlIEb4GIdSW8RAvHLpSsjnmVP7mnl0gyUHx2qauL5RkVRrrduj24Bc0ekZo98PPjg1u2kZiY
pYkulco2rNIbsa4BkBJ+aeNXhvGwvALtNgaz8ppcaO+eHGwqwrPWJ3Y7IywilsZXKtS7bbcKQK+F
q54HDdfvtknS2VczRylLE5omQZCjtz9cHJH/ypjjGTz1ishuB0exU+VPtepZGETfMyt3nS2db6ou
IHvMrGRr+V8VK3XQ/XVV3dvgVWdLQJq4gI/oKWB/conOws/ugI2DMysXWJv0dIZao8Tpfi8m8gCK
WvmcRuS3JFMtVMy+dZOcZlNnkRs97iN85pMOGq35AcxS3YnkDwCWMKmGDwlr9hoy1H3F/T7me1rZ
YFcHuglcEyQoksWDXXTuotDs+Oa9YoIun21knmaxek1b3KomTe67PSaqMydQmA8O9RXtUFeBlkWG
oypqRQOP5K+puB/bpm8RRkscsQNVCH1pHqZpGjYUBQxPK4bIBN+4Jel6Y48R28+HqmQzfavXHFsM
pXNgw0t6xlh1WF3LrqCs69cWOb7StASCf/nmaxBCGxuVS5e0baO71VjFoUFiTbsHgFlPyQ9qEkdf
O5h3Mz39GTTjrepTDyxIh9/J2o+74g1+7JHJjKV0nCpCQ41dxwuO4FCzDIBKZXjQp02k13gS1hn2
RUmhRdWd/wquhieXCp3u8LA6zXCnXxTGjv5Z1PapxrsHRnyrz98Z9UpRTIXYz21bw9/i7GLO3Qo3
9xb3ZnPY99V5TO5JGhP1Ezn8+3qJszNnh7bd6TMJbOzzG+qysbQBrn4pIBbY73LTMBV/fY9u/0xR
lSr4PapR5IV1k2fe7yLlo0qzPdaT9+3AAh5H85YRLBY6tYwfvJwQbMl/5zo8QDP2aWMW4ZVfHITE
9j7aLUkejLEay6in8vD1SBffJXMmvhP+krQSQygAlTAqHt/53dELx1zQC/+I67yIM67Nzj/l3Tas
z6hBdiXIzY1ZpwjgT1Zz3GOUUeSQAeFo6Q+nXRK1sg7m3kV/Yx8OpSNfR0o9ei45FFNR8ZSNCpjz
RHJj3+kHPATAC33lcpMZq/bwWeIN/uixhAQdoEHz3yLOq4IU2H/Q8V2Ia+UEKGUHsK2jNPSs5Pqr
/PvUL6/kqkrBRvJ9/CTNzINJytee/u2cXfJiLrhsDzq5IEFyuNb8mDxCrkq2u28M8Ff0BtKFzYax
gCFjlS5KEILZkl/1r5NRALINLtGrfTZ9wJdLE0FLxFUXleb4L38DslOcqwD5LrxeB5OegK/QB3Bm
QF9FyMMQALpKXLHifE1/faqK/Rk4LgXzOMbWRyWT0XboVmo0au2oFuhWsu1fDg8praWMYKvFRmzJ
yGO6nP4d5F6TQI24rk4OVOo9eN8X0pwR4p7n3fGrXbVXvx7z0pDsu0S0A6HSfL8aTnbk0oNpiDWp
b+cywmGgRdlPLBW3lryi2OWQVnjIwlSbuovxn+rn1Lsh1NTFmoRt4blwk7hWElaoWdSkiAVvL0qR
4Kj00ReT/9bV626cDXAFf/5bPrWM6HCoqmeM8KHChzbb3KvmXqBtsFB90vE9lazMZBq+xt1HqPG8
4CZIX42XlStmnAuRQM0MOyDwSR9nlgMQvbkda0F7Imlj6zjtYQCJK2DDVNCY7N9i2XzVV/KmzxIz
QjwB4ze3oVTMUvWU8/oRaq8Z5DAlIUTEAGpclt2g1peOiNeYfQBUxbg8RK2JSDy4E5/keQMT5AnP
B8YnpOM0y2Nj4YrhRNNJftOy8A8Uag0mgHjZIN7pS4khLV0TeIvVlOfAZ/TTDD/NetKpEN1Ur7p/
E7pZ3wM4G1LWFWvJfmUq0AarK+/7QwHu2D3mKtCUKt1tE4oOR481l/llw/kW/RTfuHpx6mRd7BdQ
qVbMDWee9EQBjKj2BrfdX0F4klPB4gMzpc4ze0M1zEpuUZQHFd2LyPRCyWBvgJzFxFJkcL+qoPMP
uzeCKwBcTLvi8invveLIqgozkP6KxjTVuRwWYSWtVswpM7yui3ITdGyRMW36RRZxMjScxcaB2R8Q
C1hPA3151GsZpCQ/jiYIuxhiM49UP5ivPC2gtJJ6Me2aHwi6sbwuJh+aauBo0oJfxeYDjz475+Ct
hswZ5K7dQTzCgiqr1yowqmfibAgY41as9C1QTg0eywJwaJHYUMFBjMNsaWBAo2HhScPC/Tq4FiU1
k2otpRnMTBAcDEVBos0RZzFRdnWeSnWje9OV4ZE4DhmVcxOTut47Amj8ySzLhuKzK3z7igm9iCRk
FOA1QcoDZWQIzlAcmmPCTI9y2uNvwP4uT1S1tkFHvd2vqnDRi/78LyatS3El9f008+UgClZZ8Szz
UTNG1No+wBGmAswT0a/feJ/tErpfj3GnDrrLhxFdMflQSIctUhu0bzqPOzPyAqFhhHKqQETTY68s
ueGq3tr4UiSwBLh3n2ANWpljWTf7bOWEyLE+9vR48adFriFspQ1erx4wDMEsO0xStUhpa93yJu6Y
QEVePhjPbw1vtxC8SGhaJjidko7BeAv0WOXQBecL3sNex6IbGL2hCVOQu68aiZZ7nKU7vj5MmY3Y
Fw/4wNjgZoldTr8E4iqJIBJ5sFvnKA7G+SPV448cFztI3PRiJlhq7cbSAZTq07knP4ge8wngWOLu
fp1jtmzQiVLJ4+Nr5urMCG4YopxJhfB5GGZ+wBatruQzmTXOuHzoVTZf3Krbw0alWDu34vFVD7ZG
+BT2rNTY1iLbrF4ryVSFSMuCRJx1RT39T7hSzmPqHQCuzls4xKGIB0J8m9XfnKyP2rquw8J5PkVi
oiAbxkdK4ofXUB/8Ayw4ByinBrUWoo88fHM4E2ViYM36z9D/k8/cyUIOMTHZTh06CJbUyI6U9PCO
clvwiBLCxKXx2jjBCQEzyy69/5vYJZxa/agHg5bTZyLLmu9l4MWwLQW36vhwRpuf1vZjrG8ETzUs
gNxa+78Ctu/wAsZkfyasqpcQCHQL2Dk74R4TrS/xOw8M6sJlL6yabyjj7KmLm8VUOnbVzjuasIvD
DqWP095bRbDkEQer2A+ImQ+nj6FQEY2vbxz2fMVMNbncplLcO+35ZGQE7NqT/Qq079X/BWIJvGKn
urXYppIia5Zxy1Q5xs3po/IIsBFkq5Hq6/nxUCdkKHBhiwOW4rMWP9RqAm5GeyLHz7gywEmjRkhH
00vbq4DKB5yVBCO1W77b4YFxC1W3xaoVf4ee2NW3odnB1kRiS4oZvOFZOVhjG6ZqfFISuiC6Fptq
oiDeU7jnF3nKesWbGR6h1eLEr6qYwzbPEitVXjqD/We6d8iCpI82oOqEeD7US91kfd0vAsh/uct6
saZLwWiBwwvvpp83mBgGytnAEwE2EQvqfm25PlmbpyRtfVTen5EQq3zMPtB5DAFRHcBQFclaQ0xe
AnbiAy/rExnDa8KJwjjGWd/pys5kBGQeeVIjxbuvcWCdVkfwrIfqfa14HEZiGCTmajTfoATuwybO
92XkahqcAJOxtajjO9X00v8NLQNhge/dLrQwB9XSs8zBVmpCz5P19/nIjf0Ko4dOfZo9HwIAGAt1
UZ5gOsrNDgqcurYlE4CV6TxPmAlHmyqaVlkXqLwCVsuQkH8FaxYNFbj8qCCuw+lQFMvRfpJm8sxA
ZxSdHuLD+WfJ7hDl3/D9n7xMSUNNl/6UxFYlm6AS92fjdeYNhAb1JGtvNP1GziZQD2XLWJDhyIj2
PN5pjW/YWgZoQC1YCI3fhMd9zQ4Nf10OV8r/+07a9WsyyO6w55JuRMIv4ZFKbf3gOj8TeipSy5dn
tkhl3TY/1R93kq6cmhbQIkXUFc/c38bI88P672ZLFMOaNk+n1/EzINSl4kpuVyX91z2aSK7SdRBd
fZirS19lakvZfglBqvFZLHVcxEQFIaOzid4iqQRT2CwN0kvXOR2ktrRtLZFUcYYxm7OFTwststa8
MnEKk7HKWtajXNFafi9SYXJfPbbtb9DXYckWAnPsnYtpof6eE2NsRYho5qyI2jtqn4kVFNaJopkE
Rsy75PDVRwNmwv19a+256IODTuipVNLzuEtsq/sS2k/r7SwnCAcn3Oz+muC2Z/qHnwTiTzE6jbGR
YBW4XNgdPDsoChYGCXDjqLzSYpvQ8/fAw8NKNJ4lTpXIl8oh5Gg+cWDn3N7aNmxS8UI3VSV3P+ZF
TScDZN5pTSDel5gw5Hxy5WC4FgZeBXXrlbA6y8yhL8RrYSY8jOyYIlYcHvxJQGqISivggdqbBVtn
60PdA+J4sDeupaUSEmIGrBm9qyFZZr+srVKr9kCxHz4voT8PFkbCPc/fkrvKYQWYBJoGw9WjPTMe
A/X2OlLXpbZVqpt3rEjXGEafDLAucLqcjbjdC7Kkmn47XWAnUXkB9e+A4iUcs2yfwqsevass3YxU
2nGB2jQ4Yq1GCBens25AY1yu/2sejFmSigpn1IgUKcRxuMQS5cEHfLKs7LXhgiKYv82LBeCpLz6P
xiS0cPf2S+4PDwvmyb0l1yv54uj/WyLs/Kp38z3UMX+AcaPvvfjK7hFAtH52uLK5rfOoD7JZW5nU
zPwDMvEhzVXI/s4BB8EU+90LnT3F46I43wSvtDzlptt/X6t/DhKicvbAmljGAKhCd1KkqxDWj6B+
37jKxoGQ5X5WX6IeozWoxoB86tPz6z1SXjuurHlbL7eMJB8DIyw6Sx5khA/D6fy9VyzUcJfOQIpP
c0VSTF0GbXfeoEgWCG7bP67deAhRMSOubKSNGcd0x7IgrkGyaw9SKPPUJdeyOSrVClhDb3jyLiU1
91ZghrcKWi9lXRhu+tj5Aqwebp5N7z3lm/785SITZDUxxf77jtpaJCQ9dQElaMpYIAXyQ2js14Ua
pKomJVoD6Pl5+ahDGe8JylQXSFWGY/6XxLfuNK9gARNPjPm0RPtq5iwhX+vX/r1VMnvKoGwnJRoX
CiQ5jTi6vJn7FAN3btsjlqkY5frWxkOmkpvvTuubQYzvbZ9prKzfbqLc3WgheV/vhzkAmY3AaDEo
DjKEYLD255lzO1HyGHL+oLgLulGWe+0A1Ucwoq2yWFTSfBODJ1xnNGlaISgDwSYtPVQ+LMw12EZR
rTt19Ih3ounh1mMWcbyg9605mtQMbiAIQ605NrAJmYegectQn9MWqQyXtxgqpNnDf1g+lt/Qo/su
YD20FqJCyULi7GyiqMAssqdwk/sersbPCZzDc2ulY0umsUZee4o9DSDlRubgI7LUnsjViaj6jUH+
h75r+W9JZzU741/sumTZT2Key++gc592j8kfu7MYVDy7FNtVzbFIHRey45zQKNAIKG0ZGMIj1t4c
3YRCTF1UvpehD8GMcNpnGcinNblpAtp65ZHJMCsWm5ZC130WtRcJj9QDG00QTHigiTMQ2cu2RO4U
MdzD3xEEprdJDqYjEee4yKFeQYnkuIe0u1LJRDaZGdcKOhsuN0/u9zvNBUTvNZGWPA9ukvIl5Ft6
9X0myVL3E1i6jT1MR03+WZkSmdVSzC7n4VCL3u6LZcnUVfPSoXJAtrqdqCLWGUhGzOcowMNR1U9i
1bve2phpm2nTYI3vV1XCXBbt5U3yA0WzMpxYkijJt5VgdZA/hZQBOKuK4veRe32a2iiBEmaQwlJl
/xRLrEGvEqKN3ynnyPMGeqgLXDCssbnbmOZQz4/DFZrHe4hdoMdDcDoidhXJhWl3Wm9/dcSwV9XW
1KobhuqTdoq5kvkoRBh5h38SSs7k6gCvmqDcihFMCWwwp0Xt6Y2BCW3gXZ+ONMXOttv0UkKd0iMc
AADsC7lACSLtF5H9CSPDRP0LWFIIW0Xti1fUjvaeDxhAcmSEEduyXo6TBa/ItGa4fwQrJ66QEJLZ
CKZpL+6Os/EK7eTgplyItMVCAYvIhXR341X43Svm4YlOpNXwz2bJ8MW4Ki/95M13j9FVvgyK+14H
OcITXAsS1ezmgxfbE7ldL/IqQklt0UdWNn8Xyxly8ZorAc3n8Bhz5d8I307kEp1QWSr8tGkVtyCa
k0mzYVJO1WTMZg4tzY9xaZHXOA8u+5qx3SdbEbl2VaAu+glzueH7b/EW2k3VBGiIhD58rxLrgo2x
pruI7BqHFgpqtZ6ueVSb7DjzF9z9oo73y+s3SZjNCwNd7kjgO2ZZcNaEZGVxNIUWjJSvHD/hGeP2
kSyrFIrq1xqRm4D2Y8JeOwew2bO06wZr0BWFERjXp5XI0zQBcrSAzErIOutouMp6TcBnR9VuD+Ig
BkTuxclkXLi0zX8dYw4+ImU3iyNct8CDR+IbjV6QeFu1bJX23On8KBn46Z7MQXELU0CsoR52q2Vd
olbZpJcPjv5+dhVI7HB1BuWlqtqUADipeIWYwY2EnIzB5JoxPNagNiZW72KLJdVP2g3KUHHmxmNl
vSZ8Q9l/AdrdhB45BXNOIMIkdq/eYbHT2IhCu92a2YScuBtHVUTh0yncIbbUuZt4wamHTyjfLoAE
5fIxej/cQ06RnSA+sezelKx9Ima8vjfGiohXVnbMnpQLsxgTXOhWziFWNJf7Mv/ZICRWLqEdh65B
XUh4lhghmPUKJ2VVYM4U9s5TEwi30cymZa2eUK89KSYrUfBj7cJSfckNfyap5+d1BXZw4w5hOXzj
bKiK6GaEn3rrANSnZJUqqjbPzA5iM/G2adOgyN4HgMdim1qxbmNsFJoTZ/OcFMXiRcSoG9jXrHx3
Lv8prs94lqcpvTC1zqb/8BMEPyLK6+/sfRnZdKc7rVGwOPGBuaq9OXPz5E/qU8ImnagseMUhKSLd
PikyB5znpZpomP3hGt6YVOWEwRMWEP+qr4WJA+VwceiTLP2SSKDb59Ns49uyczM9TBn9QTgp3y5S
RHGWhAkKF5PBF3/2+f7iWZiRhyXG9t/TYC0uuWF4vAaagXblpg9/E4AdAFFAElGbg21tAE/JIxsR
Geky3Rtyisc+3dwK3FmQsiGoSMb2p2dziij81wIgrJtnyPVvWfwBCWuxT6ZvE0QIpiby2hJwvXYS
aspovrCfQlRb5yhBuG04cR0+5UGrnsldCDYDKVlgynjaU/l7ouL/MuXK0e70CQDqLU+SdPUQQH7S
vWdWiYNhspURVYWKwdIANYQgR5K/FpnGCljkh53Spp6EwqPo3cjnS+3mN9PyoW4jjeraxblaCVCF
7m6puDRTcyjQUCjU4RvOKo0USPGXjO2EDm3/duE2XTGAoj9u+R1hYG+y3fXlAP4zGMx68Gnl2Fsq
VK2FPKVjB3ZWSQiBX/abp5srnLFnruCnht82ehaajA51h6HOr+JQ1BM1wtYDHP2KAOGQPvhTA+xX
CInyKJPK/mZWFHJnIsEDaOnBLJ9g9R7LL+Tao9MQ6h8RSmHpXwl3Gl1pVk+TtpAL88ovG4pdoRIE
YWPx/oNexSTCOa4UnvqKuZ+w61VMe1dym8jP+qnkaBq3rh/styjcWLUaHv81AAQS7W6PUwKr0bIR
8crAvSaTXMtxvd5rjeZ73Al2hydjVsXlH4qLUt1fK3B8m+gA7MyCXLTQKG7mogjiBx7IJMqIcaL9
3pS7ippmpb0k98kjgclPR2MBzfhAylsn+hmaCkN17jW4s5F9L9B3Aqxs7oHpf2ySVkB47QlzA8B7
HgYztjQAVHQtwjQhOUPPrXDfAcYmWxX9Sc0F2AULZe1nKZgvDjE6huyvu2NW68r55suZatKkZ5Oq
dFIg++0nQ5ZoX49xyktdm678UxvCy4EfJk296e4KMTmzdF2iclqMPg0+6or9TnK2s68cNLjAVrgK
wybE+eesYgOa3TCCLTdfKr9qTEWhETnLTYvfqFwKSEXkAEd3ZaTktei23rmkGqbzDs3qJj2Q6lZi
0rFB5eHnKGgxMSEDjR/SGKngcg5fS1KKRq59yD/DZvtyENY2j3rMroa+C1RimUBllpnWYTbACeEb
4DOWDUovf1HEyBpvXRtj2rn+AluX2unADYmZA6Qc2Mzz4b9JMu02A4eV8hwam/SUgxUAspIuEeeb
2MEszU/+Hse9kqCNnVo5lygNBceU0xCKJ6wDrHX5YDnHdySxhGn5X1z8r46L7C9Fxuse3ESIO659
dbopK09+d/xQI4kffWMddjv2Yh7MPUoqNo1IobdoS0A8ll8zx8CEiNJMBk0oI/EvaS5bsgj2BZuX
CtmYFvn8qJ4xbnfk1AKk1vZH3geqKiSYUvcUwES/Lp9qkE5szqGm8MuSHqXA/ai0XLgwgs0HMFcK
4l9fDC+0HM1Ht+XWEr762MWZClKQbZGronHcNDj9gIvEUdrTVZDVXwWpHGwxAMBmc+xm8sYi2UIV
ON/BBAAFdPoiGj8jz0oCCQyMtaeYW4hnuqw9+oOCvsGTObdh6TK9UgkRO2arVrMXeERAzXa9BDGa
orXnF+55/Wwq7bxyQOUotieMyN04CC8jV37vLPdJzRdi1yelkz2gpd5jzF8teGT11TvQGDIGhsHR
OxlEeKyMTt9qmwWwf5QJI9nST9wyjvOtvjc3nH83jh9WF4awTWIJhAaroiwgAvIAmoEeBeQNh54U
SW1JJqt/3sE2g0CMWi+eQ8KHtoZgTtFd9RYfBsLpk6dnGOUAHqR6u/8KX64/lWwEEq800s5QLM/Z
prZbxWE9e8523xVfdgfznDOqyFJfXjqPH0zn2rIhQUvEgPAwmJpoU1m7Deqh3dNscUvs82BxpTAT
jQUOELWc+eIUPH6izOKTXI9yFd1SQBZX8jvc1pWCUoAjKteo8oTyhfa1jHi95dTri/JLN6E/lp7m
bFz93bkLR5JjHGlIznvsKfDuJzJLSo34qjqGyNUDXeEltdWhi1vqHjCDeUn+42Qozs++k8B/oJLQ
L20HqJWYiIrZdp5aXCDwyXOWVXd3p5QYLCmTXOV+R7Q4vA8Awo1msDcMQVoPNcPB4tmgMCGEVZHp
S8mG2ufsl/63RDu/3zOQdniYR1UJFET25z+FkXTMK0W36AzC0VUCj1b6RJMdQ0cDB7aYP2ngZngS
LdfhbhdnStUrjZectUystq3ZiZPpJcWDbske76nJpq70HLO0OHor8q9nzJ2zYvSvDR4z3FJW9fsb
H12WzTql4bZ7cOkYPlDla7KJYLlkOQ6OhDPrez29jNTPW+j+81Y0PYTHb2gXh5GJhtELf1iFxi+p
85Gi7Re1iIduB7bP9axLlCVXORlzI0+rm0/xGPyDwESUwUNz/tpHs4kyTaLRjVyFIRPjM4D6zfx2
mA+p9SNtgvkiKbm3okMIoHuNVMyca/vxm7HMLQfIyG8hTNIPB+jJsqo+0r/6xIp11JniFp4sgzBM
z0atwZnrf5fW0nIk1Ytvg1OK/zsTjIY0fe8sRfaPsrd0JQwzYYJPMdKfl7nWpgY2kjDcR5Ccg7bB
VEs3ZoiRZsq+oPaL+NwsBcYpOaOddPe8bQVDURDCv5DH0vYCr23NtNX8t1KTiQ2M4ArTPzNHxkl7
TL+zxYu9AwSgiAgvrpS2bUftJLf19Pdpw5FxEscM8LZOkBfh64sc5h5KTRoJmv9sfBWQDk6Nf+9O
rSaoYxPp9mVrzRfIQvhqOfuC57uhF4EfTwydNYe4ZRPujejiWhNrlXvDlUoZgP610Om8xRHjSwK/
1IPnQaa273/1iE567S2S5KC2jxTPkujIpjRcCSt2BDSjqW8MkSYF6tctHQGjdy/vo2kVxfRD3YTI
LU+eXcj8C2clijAQcNBQyi3otww4WLXaZqMwxkRFdoWv5r2Q0o4KxUnDGCkZRnvaqaNqrUmGUy8g
DL3fC1AXqyyBJIGfRnk0giHDza+K07lBzh71bigHPHW+3/5bveb2y6vFgzK6m+Oik+e5g3HtxgII
SCV5Plu4ifIeOI3Oj0fYNTikVIKbr29Qg/fvDjTzXwTigTlAdT/b2tFcSUjmzb8a6n0jKgujIYYz
q7BgBimRaHWp6h/XUzQLHxkIiVTUmV/O2moKJXICBmaZ8rdGDIriK4RMq9TkHLgDYjeq8whsagMH
6TgVOdV6oNeUIA6BBcTIB6akZhDU4E5RpOCNWM/1DbeH8ES91C6jwT94uQwMxlupOGhdlBFMuU6M
GryHtd5O0tPRrwgdhLPdHRPF1UweC4t6f5VZxQTI27ZheR3yknz4x7N7bazxB6nAbRzbNh7Udpxd
ERuTARjXDEdS2FRbFrMQwj4gIqJ28hM/9XjzJKrMFKa52B7XcHBsw2KvQgYcM5m9KX9ST8AIh++L
NDg69cH5rTQLG/rSnNrh3oWYeAq6KIe4AljcuzN0DC1wer+p4gtrEV2X86vhsKZKz/pZxSvook4w
jPJ20A3Y/aPpuaoMNe12edQftjYZgS9uFsh+QLvfRLhsRhCiffeQxs6wqGJyx0dqM1a3CI05r/qY
FhjfWv8QOngGh/TGTMROynPSvatzG6cm8uvYS6UDskc8l5er9yOma/fhLz7U2TX507BDXcKeNN6o
GLmh5TWX+pjGF4ehEyuWTv9cd7tgwzao+0ehUr+z5129GfeGLr3YeeR6VgnuakJB/JDpDxeRMT6B
dBoorw8FHLfl3S0FX0+h/VlGg95XbFX2ZEBnNiSxMMRUss2N8VY9KUpUgie9KXMrvjyjn8QDIjTN
dIPCY8I0x/65AkTdkldL6lTjpXgq4JJrKr6HYZLIdXgpKU03J/tXvR6v31oXBnqc+Go7elHRZ/MS
6W5+frN+RKwaVxUsCcuBWYEF4QQknBdK37N2DWL7lP6pW127S41yxONCUHy6PGw6C4CK1PKhcHr8
vOrqAjorQniJHp6L72YUVoOl2KjNLgsPY9BwVYbh3H+TY4bAe3n9KeUs6WuhBro2aW81zhE+7l+E
MbJzUY0LPQ7h7s0yc5c4kXPdkx8UrOzllrgnFW3Jsl4qYHF1N/YVN1j2EN0+vzvamQ7eVApXsrMI
zz4H5yPD3/GRyT7gverq57PBiqqcOk9zq4lgC2uQ7Is+VA4zO0eqLPwC2d10eb8IO4yfcY4WmTG+
Cigs/xbSc/g4f1y2uKN2kVlywvQmX+M3vklCnShXXIzpa5tgN1Tyg6Pvd3QS7e4gfWC7Kc+BSA+Q
BUt1282+y4d9zzDk//y8JT4IrGbNgqiIuc33IU60GatXVF31KQ7HaNCOn+QhwAehzkLYVP7JXGQY
uFky+9Sa8WHrYHzCcZBwBS+wqhnkiZhc6qLmfmUYNvOLFKyIRBRXEut1f48dw6jaEj6BS4o691i5
oa9Mq4kmC/jYNkB5rgbvuB93svKhFPylevlouDSg7qTmokIV4//L+i4YeOLhQ8hbZLt24g/YwgqY
BaREsvs5m1R5N8Eni44jvPoIl58Rm6fYvaY3Ezfb3EvM6Fc2xmCUlxwgTECw6Waz4KTIXO7KBO02
JO/OkbkIvYp5rgJP6TBLXVbKAluh0ScZpu83VxgpYn7faCKIJLao2aPj8MaTbpKivaczisgQK8wA
n5ypMM1A2gnz+8pC9wgfyVa+vl6oM6pHRk4ZXq+8spVvyNM4V3aB9ANuRt8e80lPcPOZOi+tMhNG
JVx0UkcGeVy7Advn6+DsNlN7CiWnDMcZNvLOhd5E2y5yB7ocj16x8TwR/8yG+f7lv7/yjryBIj0h
0RXk+uACyLJMzguoJyrmbDXGDl5Ww/ZkcbThcVOdMZZGS6nO+SFt9aOGDd1/50TQ1OAGtyVrYMhL
tVeyBotnSTi3BV0ShmpyO+hWeKymWvuLtjFDUg0chWa9iEx5WR1U+JJ0rm6B5PiEVYouf3Gkk6bb
XSUOY1DhU8a6vLWZFS4M/8Or9MbuPJpW+lM0PVz1GMJ5eT15k84MrgGnScMM17e9xs0qfBa5YJ1+
hVgYycZ0nZQuwivW2mo6JY+rNsr8+t3Du5qEP1XA2yb+DotwL2GUt5PyLBAHqLzkEqNPD+gdjLpi
h0p9jhBsVUdtzIKZ+eG9KWcuzGEDmxj58DaPRMMUEV4PWVZfhEEUr9O3PfpY/u2qsorDR+DfsyAN
BAMRHJ22HXDWJMKpoukzwjvhfGrjc1qF/49YBXGTJxxDT/LGmX5kfLi4QgM1xNy5whxwL/5AF2tr
TM4lolFxmb5ofLRRJkVRli8+UgcHkBk6er806o9Nf7JBjd28eRTIA45hCOZa/GCrHOeuH42v58Fe
cICZi0EYY3FmrxU5sAKiaiqbNY6AlAyAKSbiJ6FFhO5h2aHFNOCLZTKbrYViIxQ7omhaSRvTFqRe
MBURjziS+CyK6q42CboiNRFPpp+uD6XKBQGSdhCIkrkDMrhts0eqnSPzPx0Fd8kfMI+9Hfp7a0jV
ui9Mrb0Rk61rFpoJrUJ2nsvrJEckuQdJF+h65oZulCaZ6HvHhmSyEfQelyyQ5q+OqbT4olql+Cib
eOe1Hs5jZGHQI7NBRzS/Fng4YRKiCTPT+JMPYhp4sEGcZK+A//uInrfSFUT90xEjyQ0NRWC10PbL
4wz3hT67Fwl2uvd0ojiJ2Aneb3mOeEsSy3cobonnS6xWFEjIw3wc/kOmm8PkjxHVfTrjOfPzZjIl
dJ8OP3Z3H7+oLnmR1+YdxaqkSTGlwM2qmyRiSMUBwllNCt+F7zHiYxAclln6192tYzkv4oHrbcEN
qMheasbn95iPcP2CkDiatEAT89PtQ6mi3dP8SSoQ0rmS5HwMgIASpljz/5wiOrf+FLhMy6sMO3bB
Sa4XnhrNBghPcXT+CTS9UGdVhjEvsTNu9FughkEvUmWJzcpZpsDNLXNbRHVzDgSnEeeGC/y7ER1q
lvtoXMnVBOTsKUK9RQ9DymPnPR/e3emgefHYZqZHjXv0qkvmm4jl0KmnZDXQ5Dc6nqiFtpdqCxC9
3ckJv4205DF53c9yMkXNYH1+qh40Ag1zQfCwPMWZsB6KiwBvDsiGGQ3yeyy4XEHrst3COXlJzhdq
PzhLqgrJRnewwbmVCm/B+GmfhHsV5B0CxDM9A2Zi7KsAkr/qwrJfgHqAySCfcyyAJfzs/FQnmy8e
8jIVJqmWDao/ZvSPZUqFZZuVDUB4WhhW05RQpiiIpzj1gkTymy4/K7EDsXX8ZQp+B0h/QkUELirK
UqCRGCq12ekui8JeqozePZ3IiTXfcXh0FC+k4Ax/5u3EX6FxpWulmv747I8osaTsA8DItn2FtWC6
wOxDy86zXHzvWI7N53behquQAy7NJfkoMRJWk2nytKEJA4849zG4ALaxzrmxltx0heBv+02rcUfq
HXdw8x9bpYVHQOuUGSMtG49wRkrnWJcAwGUxiDp3/2sIcL1GX57MQXDxY7lkomwOxwXEPAgfevEk
nzKlrkFX47wL+ltYRe9EiUYCERj/6TOpiDSQQoeaM1B2o7ALuH/mbT79SSqGkI8QY73JWF5rpypU
Ls6ykcfEjZBpkWs9YWGZ2x7UfivfDN5nBmuzNikVPBO0+BmqhT+ne1rDyuGfZl7jVWxMRiaHzMYs
9AfQ61DoNyirWKapHS+0IGLBE+PGpR5w3Xt3qedDbybUo8XxnswHnFVg7uyRiD3bQNPR7szTFqyO
oEKXGZihzWbFArbPtFALS3tg+tIGuEppqXSdCDqZp9JbNb6XdqM7LtlCVcexLcWZhaqVaQBk/MKU
6/7x3H8iHBkQM4ZSgnLH3XgWQVTj8tpEPHJWD7eU2/GWGoMMil5PckV0eiGOWaHSjeYNha+Oi/gR
fy+Tu+fyKlREI7Qr2yu0ntJsjyilzJgdEohJ8he2uVmaI/hQD8iIcWsHV3xW7IwtnyzDNmiMf8Iv
pvX3NiAUTECaQ2hCZrKSUfrLtS6PEQGT5ClOk0n0LX5z5x1V5RttS2TYTT6+rtfHjueLwrIe9UV5
DgfzcxeAC96qhMRO8mEwxjlMGnt1RJ2vlWTJzxSJwUcMcvXp41R/V6Xz7uzTxGNJba0KfFWsfNtc
2sa3g9PzQ+NvfdE6VGvZo0EkqNdCAOd0BP1zOt/bIrYumKdlSlLnIuxb0FFBFhNdJFnOjImyunhv
64RQvTHeZWp9PPND+Uo6rwYs6e/HUiCoSYy+RFFvWpSlWNCWh1cHWom40oxkyxbDTxNeDjL7xZd7
06WIEuRlMA4tn8I/hUej2wDnku2I6pbAXh6kQUZOHkmgN3rflU4KQSSC3TTrpajZJYIxWgFAd76/
cdWUlkUgBycEvRdSonBG/oZYRwuWb5IpRrQ++5ARaVN9ycTa3RPDQQ+O5d6C2+yB1kZkECu6KOtu
11ADqDcu2BY06DiL2jmuMTpJk+Q4D1Epcz8EeLtYNavrxoCMYX9XVanHZghdPURfnII9peAke92Y
l5TLDjjudDu1H9kZFIuvOxiRU43PmaTshZznJehmKUzo/m/ThNchkWRX+bskIsIRIs5r+5BnbPti
LKEC8AMuTR7SIhBPzsc5Q2nntP1HMQ0Q4OxKZZmlgj0r77JZ5plJq+xZ7uKqxc8IfkiojzomZ/mM
lzXiZKFSi7gFrVzUscPUDsPdKQVg0WU/qWRhdEqYyVUwEoaADOf4/UBEzbcGWfQCweZ4WidLFLOM
DyFHoGTlmIUUul8jyhcn4+C+Gp1FCQF3Fvj/ofi6XJd+rIEiTUgrke3nFCKmr2+hPuEjiIDijDDB
56aNTGm0gkPLLJIPti6VitL/BhBesVbh+xzVcf6oRnSStkSEfAx6VATFF9iQotTLuc7fK/3vuSxP
ljogHps7O9gUE0qoOcwnlAoQSE4hcelBzJwM8X5RV8Mp4I0pwYctmmMrXbM9CiEaSI6Lm9Gv/zXT
WoAKYotTKCqGyUTCuxj7X87B+sZKLcuCPb36OgrnXZyEFS7NLmrWKdL+4VRvV6PKJVc/iGZ+7dNE
1b85tZVYvs+W5PYjbfCdNoUPWJ4E8ieg90p22ikJl6WFpKr0vAXdWoNJIBtPz5jeP8cQSj6Iud3W
JCaA+fNTZ0+96RqMuKhUVy5elTRzfSswhnD1snuKYruGRqliTanYJfG0xJug0iI8MZmSSZFRgwQg
3C1ve7I0P+ruzohp1yKJPWuv7n6wmXMDnNMrOaplz6sxbTj5GGQ0/SVigttaX5EwUrEg+Kn42C/v
Tyhe1Kj4TI3hOhltVJSRpNSnoolaEyEtMbtU5G0l1RtRv+gyqMfaaL23YxGrwHS9x7bQhGEseiQW
ZOuCutSvjY23k/8LJ26sdmAC//ohxVN+dSSaevWnO3dWZHDklFPU+Q62CqsdM/GUeZDBzSeZnzjs
LplqWrtSOK4Y7MvIr3kNN1i9tlVLEbqcQZBc7+8oH6gSHEniMOO+9m/8YCSjVeLVjPeUxdPHXQl9
LuoJ3VBV91ZKTDf4w3K4LmMxD0qUwRxqjpMTsbHoUI1EMDYekl0Uyq+zqEN4sei4f6xaNXuOzsU1
wZkNlLPhKfmgVG9CgbEIRcPzUoXu+1eDXuEXq6mljWAbrqjKJB9OlzQHK2/ljWxxBCndEjUbdRoQ
7vVocvwb1JCRWWJ3JWanLnK0wQIUga4e82o14y17sGIlspTjPtSN0FqKrS0R0XA5wgxwsTjrMhfm
6ZwRUqJzUgz8BLeNpOr8C1rxjitgtKtxvPV0ZKqASy9CQsu3PeV0t2hYZgOY4fZ63IWCdznmhwVL
aio2t0G0xNT1OAtNzCY0/jlxZt0so+5HsR3mgt69456wl/LJ288BE4SQTRBx04QqXqgu7ckfjJZd
c9oAojoY4Bei/kfCp35Kd/l6Gih80N5QVjSEk6MWPiBGnhGLb41sYa2s1uQ1AZ2W/g4TnTDe4yxj
pOD+iSPkvrP4166lwojKzRB1yLPRO0k2ykaVlKF2NtOs9UgT9ni09eZNVQZ798m6TL+D6SPPpitX
FLwbDbCTF9WY4hmUJPw+tr+vRye6uK82aWpCd2uApreArZnffZuGMk50we+fVFOEmix43CWk5nUE
aWTjbXR8IWh1NXnw8K6p8/tFdRQc25RcCuIwd1zaEbQ534rKVN51i5YVAK7me9ChGGFCh6/NK8YV
nNDsmoDiHRd+NFmjL0ilR07PqxknnVsalkSbbu6r9yRsFn2/TeyQzEPmXGb9vTou09PuVL0bbYMY
nf7w02yKOugybYsPGOid+Vs2uGdjeoEEawbxcZMn9qAVKwyyoR9ArRm912qHkckB+4sg6M27aFxz
zHqZqBvsOYjNTi/VVgOvg+uQjbY3sJjnooRhQ+7XU4KhKzIM6F1n0twSv8voUwDQGRl3h8+RIqLV
2vAo16JnWNH9ALAXD33ksaEAkNn4M0Qc+u5VIXZ9IKHPYjS5Gnw4toOJ4CFjiZVtksh4Tfxi9LBB
8LTqFl+sZsQ9awOiMYgI9HC3o8AB3xaYbPV8N/OMQ6swwgk+Rt8lg5audIeOkmBo13zf8azQujoy
v/rnZQEc8fMcG68wIZwJpmxbmTYS22q8BV/GwHzceAJsgNUoGh54oKSEFS91SuuM/z4oX2meC4sx
lfD0hb7gfPFXmumBq1Wocso9VLfsvNIr0qrDf8EV4Ia6GfeusyG0YCDSQq0U/QIKsSTPb9HHK/V+
Eteak97R1dAF17R3DQwDeAqX8JnV5d6+HYS6fbs6wYcAVj9rU1fNgUBrQZwj/3JnAaAZXESKYNDM
uL/AqcffFxjFKW4cXqDaJcNmhH3q1Ul/MgZyVO5VmMqUncBaogQKpSciIE6KyVif9jHYuUowIPF/
h0LbRtyg5Pm1B0OwaHRXRWCXGvDSyKSW8Iq8I41Htvfv9iw+P4oPaYvpOsghIUR0IYBjyaruq6vQ
MZjWywWPj7OFk7EnOdwICOyRLLqGoqxXUnEgmbmdB/L2Kk42QeaVXd1dObbuDLnSALnYr0iFreXZ
tEGAYWGW1vQoEY0G0l4Qd4Z8AgKIHJWJrilbcEXnuPbY7bfOOjaAFLxuZQ6J9Pq7NeTBQKd3IBAa
GSbyptf7gDg019g7oqCIOgdMq58b9kjfbCU3kuGTfMIhqObP/5hu+VoRA5PZHOEhBf0MfkpOV5yM
rJse67cVVPfjQckjz9qQ5gu67sjP7ZBdQe6L/C3UPyGI6dSGjnzA+5ExOHgh6oeVbmGEY2Cc0FED
t+AAgT6Rzib5nVR7jtgvfIOpWXDo17Y2ptST4IkZbNoMuduqHFJLiaX+gY5I66O7GXeOr+JeK1t6
+do7qUk2UELRyU2/MHzyaXvB8D5QObm+CsszX9PI8QIYX+k9O3ypzhBB7laLflQQNvrjC5SKf/Qt
l3Kv9LYBTOkHJ+pFLYYxiBZCCxkDZArdFAS+zM6oce8ndjlLbsiH8x8oL69Di8X0MK7AzFHgl5Nr
fKLBuTX1iJxYHrbFhiCPoA/skp8axPUA6/jKE4t+FubW+2qZ2v84kny7UWJQ3KMAaKd9qKBsdvhT
1uUulOhSX9JrSTyKwLzymmxem6cYjFkHisfelOzqAezkSisoK4enHE5heBRMFYUI/IOeUIsYfFJ4
ny0geVUsZFWiLAma4UCNdqcQuiygrLqyJB/bJiBGAn9ZQ7SfxSeHYY1pJ42NM+pdAbFKW5n+DGYb
c7jz6b7sBpVEsQa2QTDE94o+lE/EniyQQtaF6+jsONGCYCIg31Xk7ywdWDcQH9mQrJxpFLdC/5ee
vSTQMcEfxqjpzCIdmgpu6ordewooLyCyN2yzU2qPwIKJTbQqLFUxVlcRSUaWTE5hDElbWHhDa/oV
ew6iax8ec3MhQXn/xGHuK+MLKLw+qNY+Wn79h8sHV17Dne5zBi1sAKrmBiTYZUDewUPyIsri1XEm
T58xAPFNuU4wrscRuYFC4bZNam1RkjQHMiLVhcAV3VJodwLH644eHpkm9U9IDmA2aPJkrSayv+gE
vg39zFm2i6TImpsYbPfEpCH8YAdxBbGN8hyrsoHiXbePeYsV/AOS5uxv0ZQctBAQDNl4lpKoPwXX
d0Iramg7pRfsGQ3HvEC+FrP7aSXaVPaLruBfsywxrzL67GoVDT60HTkWqGjK3hkeJ4lCkm5b3o//
ce2WhxEI8UW1xcZdK/owk/PLMoGbHSLMEL3C5fPLGCIVbrb3ROq5X+xZSoV4h92UTHncUN6zMI02
tegIxH5w4U6cpUlvbOyogeZ1pQuhdZose999gSJKeELiT03rev0p1M7fOlj3905HYsEwdS3VOOWP
n/LXTW5ivHYjImLPe8buGDMg7ICTuX1M/B1aMk7HuiwS8U3A5LsKmYfuI96AyWPhNgyazphXWhJ3
TfhchmST+KpkRk5xzePwO72YXqD5sXGaKiwVsX3JnmrgYL2sf9NYUCRH5IxG/8fdPgz3IpAi/ltZ
AC1XmC4Zacp6P1ChaXf2TJNz+1PDFJJQLBvGfUPfVhNYgOVQCI6z/PFCaiEZcke8zO7619nL96nD
/OnUKFCdlwKGSI2w3UCBXlC9uzXEc+DtKZiK4gQmvfLomao7JtWxXC0T0TrrQZSwxI9m12O1sX4s
BHCHyfulnKbHIhp2PvWR1z0qhbPTg2C6gsx7rk0lFco0bEYEeABpwWO4a9AGwbl08Uy6ml20fM2h
e+2adNDhMAjVu11EH9XOzLkzCDoScS/010Jg2l2GtluElHJbVB3yrrQNLNowT/GSWRW/BwUynH5p
XjMhrVSIiJJ1d/BiJZGbyPRzaeJA+L8RuLCURh/Fvv//npGnW3fAVF44okXvvW4HCUM7GWkL7eUS
PMIw1iNaBZp13iG+Yfh7Dg+IjHAYMnnaklN2sJcxyzQnmir3RfbG+cfnhoJnpUuHOi92HBwjNPJR
9PRKRXJxJLfspAUxNzUd+L9uVhFsB4pmmUL3jyNBNnlc8k7OOZmgWRucfZU7191ldOJMUoji3cnp
gIDBm+HHoxXZg7HARuzowa3pBBeFuco5wX9d68AYZZ2T49kOeb+MeFlwzfCniqonaqGEHee9RAAB
I+aGm9IdvxSR5AIT1es+F5eMxmVyMaBCJkrLrNNPZPHduvRtRzxydYPM3wtsJ9FKp2vOXsty8PTl
H0Z1DOsou0lcz/CmWA4Pd7syNSQL/AmK+7Wa+NI1iAxFgfaFa1pVfr+0B+tkltXBkoT84r3DD9N9
YeZRtWeM/LWHCJK5ZrLJFELodDLSXTwSBLyI8zA5EZIi+tKDe3cQkSPhr5ZrimJ0p71cl9uJcDKo
iongVYrDEE97bMS0WPWk+IixUel0nS7vgByVTd9SFcElrnTgUL+wZEsNMsjaxx9P86/xEW1FLzvB
IZpXBrNKgTstOzMkSeXThhUfmnnazNf0e9jqic7/ajoWBwWAp+4zgfhCG3OYbo4yJfYmVz50xxjZ
2jMkoB83dbJIJWPBlRYTDHKamxjmYmBTDtdFRbmkYekkKR6jXEi4rvw8UrnPkIRl4F5DfEX9N5Tk
DM5Ymm4DCwXSx1kZlb+xFKzG51pb+Hh+HFJArBFpXKiKweK2HBufm0bGcAUAGxCrkTpTQr9Ntgvb
7JV7xkc8TzQ5pwRpjN/8/Q32sH9jJ3LBILrS5xWnxpDjdeVZeaVj2FactWCmeL1zLtkcTzK2r7Rf
DnMeiDl/FF8stKsYP0vMmnSgAnqUdXqeSVb0+1o81bHvCQ86oCBYzPGt93WZGXqSAooN8drUNHuH
Yl716tJzVU/QrGeozBkRVDGzpu6c9USAPrz7fGCFWmRTrUvuapBRPVuoS93/tjS/dGCWVRS4xu3G
z7s1WaJuKsABek5pELwMQBfLbqIU/jmhJBv0PLj+dtakNrtgsgPzcCBaQwdov51jjKJTfMEPv85z
dwKGgilv75bX8Gn6jhW7U4WUgJYMKrzqReYlGDOmsikFxDcnGhQ4yokk9KVMAHFv40KKFzFK+Tls
KOH8LT+Ss6gn+klks14AZgAT4nce3/getxoeR/9YADHevCwOo2JDwYzXeEEOA+zAl4nJ7V+/nG1c
vaB7v2zLUYHDYQlERf93hlXmkwruoPv8nDTPpxvlIa+Z+9FRWu2xKsVQYA8NICvpAhOwt0uchufL
Y065v5RGRi1gDqOKzJ656CcvG5SfPedZ0+R+PaYQMH11mLqub5aYEoCJVPgxdY9z/a/DJ/J7RQ4m
ZvV2tA7HBgMZsfwoSZLUw1hZf5T6WWZ7tGLOZLmN5v10Ue0VI+HqTcGvV6J9bGttFjksv8rB61je
/9X2Ah5ZW3nVFXj6whukZZuyyc156OwrFU0Zanca6i1hKBWs/erHLTZY/JuPBKOMd3xVH4MtebMM
XG0jRq0Or7LAJ57PIjmKc1vCLx3KneJhP3f/mvbO58S+3fXmnY/EWWd+xOdSknyh6sw3ofoBoG/X
QbyaL7WwsTgCCN6rRxmjvdaOJrBCwVS0BIE2gcEgInWaroogno/mTnSm61g0LfGhz8RElQP8+thT
oPUQq/O1GDbWZh+wGqvyfh9r2hWhiKPSoC+Ctzrh0h4sK8BGKpmxpZEascdywWpDkZtZKTrCUndO
5PmYUyA9c/ASuL2j5O1lGdP1gpVIIstroM+X4ZmjpB65+Qr9lmPI2aj1PyLIG4zWel1Ldw+61F+z
0rp17e31Yv1Wxi2HXfB/1O7F/s7AGel8REaOPsEI20iGchKwvZhpiSfO2fVWEWrvT8rmRXLZopFA
F/aMF20NrZ5/l8islqUqiGIEogUQs9atfbwVAsex+cN8/djIn7PJrLZVmSCNQNvo/38xaWgqMiDj
x423d4Cku+vgTwwjkuMeMExqNjZgqCuFcxqIgkbDR1GMIVV+0njZ8PdHiOhMkeY3hC58Mb2NUURS
qX1hkACaTyJtxD5rZwA7HQp+mC7BVt3WY+XcM/nEBEFDt3nYkKguy6mf5jI+/RyhekB/2iKRLQsS
rmbl3YTw1bkmyyHpYjHTe0CB7IhPdX+eNHNdfyI+hV6KrxCClepCnNN461JP9o/FiCF5Yp/LFfbi
xFBZPcKcFIUEfL7uKpCQuLHe90dkX+wNCiOZs15ATn3Y7y+UiMWPeTDoap9LgRWMBHIwkKrXBxlV
2U6X+vl/mVroXQ2PudVVm3X9Kdfy6rCoD7m1kP7hLcQVCqQ6rPqe2KI1dw7xjLfiFqwBdXam4T/U
QL4L0pOANQuYI8xjTHNTIKbt9aElT5ae9XCe92MANFxIQFHKTWVTNbnjDN/Wi0ZuRc4EMunOPHcG
ayljUFYy9zH3ZiGIt2PMXzFLFJ+XoxSU6j+Uv9iXH/3azsNiNS8yR7naYPtRxJNsFX3TRUl9Zzk1
pnXmnSK9EXqfp/sK7lBOleA/MCw5i5ORi5PUo4aWbrtJddWr+j/aEaLpnB46zGpymzfjQ7oC8QNh
GK7GKCQ9PvWOrwfipqdzabOObFziXA3pwV4RUX+axbUdUxecaB24IGVekDxMq/nGfyWeHDRTGsqk
Y3o52zj59yXavruCCxuUeii1hDEw4EHRDM59z9juV19HwaXHUZXsnywBeFnBaCHKetIS2O3+vcup
oSfvj2wnfg1e+kw4MhOVe8o2my9KhDHU58S+KXUmMLKidLi+DdQZdwUuIDPKmOLG7iSqdPJFFWS7
KBCbrRxbajeW+YT4+rvYn006aF8ANAqWrOsML4tl3JyVriLCtv7u56ZDz5Dfted2SqsC6JG3Wt/3
gBvqmsRy+Dyy96i9uRe4DvTjiXt/+QeidlV/FkpU/iaiLql2zIdrQ3MEPhuNIFfZhGhA4xHYf9kN
Cp2KGVlqDd4U3kBMIz9UXOIHb32ARHh9zZxKZJkSTqVH2Ck2H3QzXbPOsMptnxOoAQRx2FhEKv5i
IjaJhiAxuzlHUZf3iRadbYy7PiCQ0x24Zt6JIXjv32v+kvVvL+WCjsK56TnGBgSi5JMT097f12JI
UjE52Dhp32XvxCgkHDyf8IfoIij3ONvo/ULnpwKn/ECd+7Ki4i2gcZqrDQa0YS9SZJdT/m/yOeQd
shMifqnSaDd1VOQFus91J79ewN8uQw8NTO14J14SVjdRzucXG/+/zNLrhuwkbwcVkEpmoWPMHsZC
0a7UlKsfGWIWXiYd9p1T7HscbKb6/H6qrBH3yGZ2626ReeLuM6QBrtdQAwSpLaRaXOZ2taDBr5gk
mvncZ8ReAvNDBcUU1f/j5JkK082nxVAdlW1/nX69AWn31cTMRJ9bV+has5LswwWXqLaOQJ5XApj7
gX8t8LSp8NAZvIgg7Bsda8TJSx5F+O/qWDP/FARW5zl8ZbqvthZH4t++yd43cOmuZBVO/Xd+VAJ6
u4nq6A8c+SB+glc25u2dl/Jmeoz0AZMDNn/W1IbgwBLwryRZExqbro0YGsiwXFofPLZdmqyasIhP
+W4vjoI9W2HJo+llyK8RqqSsAtkLe/LEw96MNGpHOPjGndeVuI8ufH/gDpwWuyCCbX7PF82NKWpn
PZeuWo/l7UmhQoq6z/INt3cZh/M7B7KslE6IdTSvnZDA6mtoZ4uWIeGxC6zvJ3zrAGfK0Bl1TO06
VLfvf87xNECNbH18UE/X4Cv/+ASugDnTgeXmFQgMHuvjs7NQC10ITrlCh7IgWDX7pLU3IIiVDC3e
YQccWkPKQ7cT6Bf/MNM5HjgAaM1JL2DvXg/LPGLqgtTXX9tbZHar9wmjm/j3T0xQj6jF4uX3w1bS
dT1m2swCVRwZipWAi6OGWpqO3mbEV/I0Ra1PcbLvS1YBik1uMMC6CpdS/EOMzjFI8VVzohYSTFAF
Jx0KfzvfDC4DRPy7EDAd7xs9WkFMgmEtiYdB3Y76Rhe3G/Px+o89xy0w6c9OUJx+cc7zHT1JFgYx
05BoJ8DJi780VTQXvhTzwVJjRiaYeNixmIS1P17hwG/hsDNIkprIT7d/nCBPZJqqTXx4XPclcq7V
ANW3EVrh2FMKEkD0EWUbaRj+9HxDEeNpU0iqkZJgZE7nr/3Aja1l1mpZEh4wv3qzOEgwtRozcfZq
MtzncW4mVVN39i6nHq3UdTMNOBy5TQbu2aVLgB6R0IXFX783ntqAiIfXj/w3ZmlK7RHEtPHWlYGA
NWDRpk3UHRiGvEt04vx3nY4zxKmzgKuRzeYPc7YryfmvOfzZl13Fha/UWrsWHD4gqgqL56rqU55T
vXwqLV1NbPhJ76t2yphloLPsyPa5MF5Dxc8SW7pxqKdOuAW4yd3VBmFdCAjyw7L+OoLjUxJfYgGH
Pde9lEotyeSYXYl0d5eoO+tFRrAtx7ngh15FNQn3vn8aKBAkvCnjs+mC2DlR2Llfu12u6XRS+iJR
n7Lc7B/W05OdM7n6U5x4FWjOxclMYRN+pe368Gx6cvzDnXeuGNkm6OKm5uFgc5Db86m1tfI13gXY
jRpli69a8vstZLHik0Q6sJIHE3cu6jneeFb6O2Kta9Hyvu7lHV2RszFsEyb3gfQD79VKH0GOIpqp
kysqsZdiuVy/TSyUnropc89jbpOAiMJKXK6W5hOL03PWrjVKEmSXG6bWbJpDk3A5up2xYNwKaqsl
JwjPfIaiQna2RozSn2F6m6HGMZW0eV/pXvxyStjq365Aq8ZYzkD/ue+JiA8UTgyVbMJhpyelYKez
JiK7fk2E96Gq5nK+IYkRRv8e3dU+tsQU6d2Njp9gTlqxMG80JFF1kSrntZ3QepCKwD0YjkfHCsGO
6Z2GztIEAkvYtUaHQ0dCS6j696jjIfiGwaS1OX0f03naGuTzifab0ErFQVg7qgI0vyN/wHsfHpH+
d62in04HmDRntkacEMDzWbJBOFYWrJGGIQ39kGKPfGlyDqPljDvK7XqpGTn+hq46Z/qP9ze9uZ1K
pi2UtUNOw38e6NMIeNZA2HXyBWacqxH9p3Th7ukQPuRarQbw5nksZgKPhFsrkuPU8q53gtrykM0N
hNWycjoO1Mvk0rA/pSQO/U/zZjFIPIAdVJuKQ+1KmkcDksGETZNgqhrv4MWqlzSnZGK9WpGTl8JU
U2zEgr2YID+ownI0hO7pJQpHqW4FgX6UEcMzZKNNT1wh758xcB6CTssSDsXLRFbj8jlscsawABoP
qdNH+Xg7xzIYPIXklXT5dvH4Q8581py/Cbk+zyi6Z12sVm/wCLnsOq1Y0+4y+/taNTk9lpNWZRiY
zhgj7912u068+427TDWsPYwxnaOYYWA1tCmHB9guM4jGN+o36MSCV+//mgNbMyyJ/3UhN4O4B8/r
5OrnOlqJC5jjw7l8L6GWG0R1pcQ55Dib3N19DWtewuGWoAdWUkKBodBel7pzYzadGlgqGHtOvx1b
1ri15Bj01vl9/huAdzv03nWpSaIzzAfndu8900BllN+HkP0mtaLNKTzHgEpkr2J4va/1cphv7/Nc
qPgA3lx6vzlQixtcH8PhwpQaTqfYQCIF1q/zomi64qwPHmqOL8nS2cmIxvyxPVPq3UhAOAfpOR/H
i08J6Pq5tyxNFKw3XZgGw9rCKgHiYrNoVr7fipbXXIE5U196OH2AwiRR45KeQBBQYTB4O69ZycZ+
4GynugF62LPcPTZNQPYj7yqngPjok/AfBG+ljsrflo9Iryoi8bAyazNFbdM5nFoXH+7A6nDyIBGU
o3UiAsnsnuklLmtAw96VXi01y3IBnO8iKA2t/ZN5OlppOxv8lvTYo2l1ph4wXsx2u0GtW9hZcM3c
OFzdeYfVQanLlBxqhV66kK2goVqgi8RdK32LYSDmsiDQOUguXsPetudT+RYLOZvr7CnLIKp/0Pbd
qpFfqnlnwoCjEFfvEamtYLThwP94o+flolWbzHJLygS2Y4BABRfrolyxtMhPkgfHG/j6fyLkLevg
ApNCi1tdRm1LgyvxzaoonJo4GxKt5CAguMqc/6nV1crgzMEvop/N4vcHUVN+U1biYeJTJyfZBFF/
VRa+VXT/w73bVzBl2Lx0nPfT7o6rZAc+/BowNqazM0hdfYN3B7XQeOc/CSjPbsyKtWUzd+UQjYHt
l04L4mNs/FTrYUTgb0BfuUyEKE8Bc8YyB2BBck9zEPZwIkWaHSSXUb2pus1lz2W1GAJ0lLLiYaD0
tzDFp35yOyCY/k6kX+opU9mOXsMGKzMW64NJPr24fvaQyiBHj/y6yxWJSNyeoRVpArWRJetbytSp
F/ukwekBtfpkb9w8+ZcxpR+TUGVPtXYsx4oDxWpLhdmr8TXNkzghLeOSl01woPDisx38KkRGe2sA
3fh2jhB2j9O9yjNA2pnTpxUKqHfKhZnJzd1tGOcMr3ljJBgoUfVfv2wNUfVX12xO5uJXYKikZxXF
2q9+/UqxyLxo025IwU/V53hkkAjK54vxTkP2LJsnJUFLazmyUwjw4m6FAHU/qreVmAR7qVu0cnm2
z5RapYD4w27+ctzvia14qWjr5j/Nc1O/kkVz6b+c3PeDLBxyPP9+5iArAdUY6UXnC8LN6trnFaT9
0mOpUpSoTSFT/3PdJmBXlEvHOsZ5ko/O+dhHq4bDwiWw0WP2NtDsIxXr/VkB7Y2eWsaZcGbczSNZ
7hjR9W63zjHk+sE0dYVj3+IVS4Rt158PYUzaT+dTAvt3/2/r0KIU8U3j0AK2i7/zy1m8wmjOIBJQ
UbTPki/KFSDsfhnjqtV08mBP31PR137B5tF7yJqYmCm2CRKMS74Wsx/we5y7dbZGJdKocBWRs/JR
uNjSDS0enrP+8NzVsRgruC60fLvX36QONTwciJxvVaclsqOTlHFlrXNeEoCp/oGjykjHCPWvD/tB
lywk3QwkjLz8dhBmW2QylV/KA4Yk/B/Iakvdk3Ij5vK8wtGLnge89EfTCjc726kGIB7NzUQ0gF61
Pb1BMOCuwtbVyi9UnYI5XtdPrEMZqvE+YCN/Id9mPBS2uDrqcugAlFiYs3oBZhZq7iMkTMwkkpCb
RcLtni5EQK09FLPrUzLFXi2XGYPamo9pvCrAepXwxSpiPYA6uUB1cM7iNljyx/+gAEvEcA+VKso0
JyZGGcnIYv1V44yErKizDF2vbBcTmXDmlj48RB05QKhzvGIbiA6h2kmWS2IW7xfDR2UFWp7oO4+u
byvBAtS8JryqdnDC74M1dGPT1y4CWtVjh26gqaI493ewEdlOLpviAplL1VvBOhFWvRU7OcfGlDqC
a8GuMc25cVgPmgwkkTBG2cueRjJOxfNVSyem/N2fkcQHXYM+zALnhfNmSLGSXp7iTYyZQ5FcJYnd
qaAv5+Mjn5naqzpUVD72eqn1DDOwAqRZt2dHlcSKfAT7A3QzSFlr7uoXdwKkB6Zcb8ghFMU8DHiu
G25ZLVoFXUIjD3ACObjfWR2KUi3Ep+EopL6bfiRyx6fa0r1KwPBoMG3jdOlkwyGWOP6hCRBWj98X
DKGWukFKYQEJORwXyThdNKd3+pJDLBpy1G1p6zCluoQlI24z1PclswVjRRsvTH49aSTnZHUkmpz8
qds9cz0YndDisPEydZDkfVtXfdOXvAFID0iu6Ye0pBSK1TdFNsdA5YmtSCnj2/T18GzTHm93mbUc
BMC/KguT9l0I/MziYEbbBZ3yxxUN40G/Hj37GX0XeWkN9EdqTZdwoEzOClz1Uq+kT/Zcw3Id1XSk
HOgxF8dPGFVYbFSWdjOk4KhZm4M4GtyGNrOaxOnUvbQcvUDe9b0FVlFPymFDYc7J9vOHiYdKDrqS
5XAaXm2MaiqjW2ugNO+3rDfcEcZdrhF1tdnMRsV+01eblj4ioZbDj7kAw1sirzVCCTNTtBTpEEu9
1vViNNhc04nvsDDn9HK4E2Wc4D7cd7783ojmkUb4d6e0vVMntfVYuh2kzeu0dlel76stdUGlZAtx
MQYbPdKBf5WsghilWF+iOIOFTdEJf4zLN94zGmMVGnZYLbQVkDZXbbDAYwgHwU3LpDaYY4P9/G38
NAB18sd/ymKzyuPdTmTGjSCDg09Rl/3aNBocFUzfoE4P8GjTdaBDZG1DcYUOPCpoFKMwNxKfXgH6
/j83rPTCDAYm7Zu5JsgInpSNn5KrwMHlYlrhZqbmE8vewm0xeTT/dwBXN3+b86tObBLJZQxo1FEl
Ml7vErvWvm//KMIBKPCjqrujoD2Gj19WkHMPhlOxFR0n+3bbWQQhPFg1pHef8nI+eZxy8ityU0iY
SHbkp84795gsS5s8d2qBN5fznY2fu2C0Iu9saTejzs2IJa6CMbL99LEd48fzDUqz177y7Pb96LtH
crOwK+cNZEEyvSSRVShXb2OS/BtnG1MOrmCcxxWghgTUwLzG0u9y0J6Rz6XyQEEsVn8nK75mfGcD
Xjn93C6Ef68ZNVl5Lf/z4upyBgqmD7K5sUPO6+pLHRvhcdoXiJQ/6+RE0M4K31VMZYuJmRUWnQhr
RnsBIUJ9It/RCmFx6SdviDtPAaqLQ7JD57hTPQKDZecfnWCSw18/rJdCYaAH2tjlSWRd0gEiKfba
gCypt8xoSzmP4vhQ+rfvIrRugdXMhPXHpURP2mgfl00yWV+zjQdkfV56S7QV0rVZ9MQIheH5o5vS
Ftpabf7FIrCvZFLTnwNWvATfqhmTMRKqU/5Tti+e5iQkWjehbzfnB6QAWX6yAb/LELAm9chbsQcz
0A95vAOUzz7FxmTIS14dt8nqth65izDKO190L87uLgtF92dyAwlUFESY8hm682C7n8xOfK5uKCDV
7EEtBR3laAXKklidSEtQsCOYWbsnwz/4vElVDOhNw3/RRSQpsC374KVApNQmohkSXGas7tGkKpn6
zaLRXAxzI6jSKCX95PL9neZBCQxwEGUtJhehZ8HxElEW6DOkApKToyubGgiDAc2UJzUwkE+fG4wt
D0pVZS70stfUPmDLAl2xOQXFYOJ8dRimX/nJ4shPcyB7OAToTt8HV5ckTPvJDyDiRlQWWzS1fQf0
1gj5IrKNcjK7/hu2q9+7aFv22qs0zbpjCVg2eO41oyTzpg5CDF/5FyLgMivq4ywcM3F90UqRMmNK
NPQ9Zw3G9lgfhgFSehL6E08TQPja0j29vp9cHyXb5os9pLEmPqvTZayW0wrAHMJ24M6eXJ2k34K/
HtKntZFDWfbJzq3/uRKO0GpnH8EISE3WXoUGnmNwBT5C3tKlGYW8Enqjzlb4uqOmuUgygyu9uigq
/2bovLNm8bsQQGX3Ya4ZNad1CM0bV5rx/zajCuW5jEhZnNa1xWc7ZLKQOX8y7Qz4V6wiskGa/iiE
flr1opGvuJuv/zzF+z3URP0OVQmoENvexKZykm9qscJAipUe3SL1ZEuymXdMGr0VvwutbDxoqi2/
O4mzta7IAibrrz0TeVfMtt877oPGvo+m7SJucgJYluL1NffFL7XrpCXwhOqur82iNpFiQ6Hu1U3Z
FK5vuUUWiKnNtIVtWL3X3RUuejomGkxYsd1QM+UVoheLpTuCR9tIIAzb9hvPVvPL1LEgI3C+1xT7
FrapaK4hWC/XUVjIoQjUjXukaB3db3QoVwh9L1tUhZTeHpJ5L66aCAHNKfgXdeWNNxSS0CjV+l9v
mMaJqdccvd+Mp7slJnsiG4Mrmi8Xpv7wpYgqiHLydvJOOJvYTu8P/vM30OQ0+/6jmqrXlHH6i6DP
4BeqaKOOpxKIFJ6YiiMK8TcTqLPy3DEFuh5xYlsxiQ7vybnlu7tH53bfhBtp27DeQ0Sknd7CUKX5
9JzyKMiiPG8nXHYAykkeUWupeG7gPnhpPn+D4ntwSbA0IVfkpmGYRsxQcWQWeePRVak078qYZGOA
q3sc0CfR7KMN0nYjrlnCsZNn2TSwijA0cabX04uqFTJI0Jhao8pfqSAO0eoKlftR+8bKf7xeV8Hs
XNGl/FvN6YbU+s0FcUiB+CmREtN8gv28N+JwfU5DdhtS6BDKQltyJspkCkl6v1b+MEeLYC9dB7sB
J68jKW7bNvWNMXuBe4/5b86m9Ou30sCmbhZVmNeTtJCOGw9rRS3VSSEtRx8iuxRCYZ13BzaoUDio
88U6PSnDmSE6XE/AShk1xetSP0Cwxl+wr50dt8sFSIe8yK7+HG9K+kyK/1DkYtsGlUI1uM5vLz8D
fHmhAbktz6zUdUruheQEJGaooly54R7gmcOdn+VJlOSKxKUMG1f7+uXodMC+DvhGiLltYFNfp/ly
Rat79Eh0nc3hrSwbpwr1O2q4mutWeogfdwLekHwv3IeUQNEE+IcfdQDnKyRusP6gBhhBgMz0aUmt
CtB0xkSssEA8/gQt9lk6FEKVfMnsUtA/DmKIaNHfBY+WrAdWrLX0s017pNGf+kHiojlbnNt/Uwie
jsfpH7l46Pp33m0xvv5rYdTr0G+sga8ua6H9843goM//vN5wuU3P6OO1pAhZMIX5Zw+ojdtjzASZ
yWajcOwitDpXMg9tkhAsjJECJtbASVLO5+fh8THlwealRuxfcffPAxVce8SazrfvZ52b8+1tL43l
+ybABb97EXNEDv2HY057x11rKsJW11BvXbvu/Xm/qMPpjfb0FJvpO956A34BtgCKvWipKp3ti5jk
YF7fkwIqG7uedEtaCNgFLGyf+U47vqd5XBxHcGqQX3W4lJqSb5vOZqaY6RJaLUai3x8Gh8rT7EUW
A6v3R4ySYi7CpTOdZ+szS91kmPMHPl7AuUSdu1SsKgpp0ftf5Ev+5hpGk9A0RLQFbSV+EEADDl4r
/6t/edU/0qKjWrHvGl80BSMcYwqfXYrjZ/YnFruw8xAa0eBFnPJTHWBXm/V43TdEmalXzSzesrNK
Uz5uuL+BinB70P7WepfouWlPGYR0kaGxpAbCDY1qNbPAlE3V9Wb6yJyMva+4d4tIUwXr8YWn8smh
5PeC4sOFE5AhCbMcGhLP+NyhxAuBvnK4SbK54FNLVA0tu41mR8nKyeEYjpNkziUm1hsTE15eVYmN
IdPimXjOxx48CltIyTt7BOWkAfnkzBgCtQBUv/UcPex3K4CdQz3FNBmqPhMNsoJyuRYnNGPC4h9N
Y9P/ApBni/QGmnu45FeMiNh90juq8bL64Ux/q6UjLni4w3Z6K89u5V4Np4/qGsTeQ/lC7+jheX32
MPwa74HvG0642X1MHCDb8zoG7+geJACvEK/hDEhljWBDyhpF1baVPsd29TLpnwNA1o6G1efn4SYP
fc5/AXNrhb5WKVjReeEh8r6JAvblaP3o1jWmyPSTpjlAsT3kfV5W07NAfRkvog+0dB5EwAyT+RYM
k2dR5aj8Nzw/IrObApiX9dJTgpVpg3WqiRtVqdypvAk2oT9n7KTDPJ9yYhHFaRT41Inqp+EiMuFX
vy9sViKSnxKDOC8iKv3JcgBXunasKnH3X6EoOAGx1uBbtDCFRqdPETl+yhNDa2x9ButvwJmMdJ00
h9N0WvhjaFPmzEhj3u5yaKcZ5dxgOiUTAMJJIlmoMeZyarYHQA7mnsd24x0wn8tno7H6Xnipo6Pq
bPvOvsznNuqWW7/3M85gkdvNG32RQYwqE9zhR4qAGdYmy1oFwf5qHlH5XF41ljxyre8YG5vqK9rU
KeQxduRtxEzf777JCDABOJ3XjlBSo5vxYekfhhA2BFjBkfk66D3S1wqyC2KVtQxZxRS6tZN4LXz8
eifnYTyMiADw782vzJP0vvn016DZyiDaZNpijZH8kr/q/WQHf2k6uHHI1LvljpAreVCHntEX5YpZ
a9mUEWhMwDcFzXkifGGKmX8yir/BYgVKYIXP8HhCNY6EgXBX1XVvvzDPxaZ156A9Hea34DFpUuoH
iIYnxVqubOz+Ac9SV1PzQgfc+usuv7wGQLVJqDFyPIj6OsSlkZhere7WAvtlYwHwSHm1CWNQXd4N
QZCA4SV7VO1ll0cxykn9L8dgpqPVXDU9O30NX93xm+829BSX8Vr9eQNukjd7BnhhpBd8xv9DKCBJ
guAaXyXjDqYu/SjEdm0qPYmGTh33rb7it7VgkWRFslVaAOEqooLUei0QDUdljcsfMlxDcmu49Eq1
Fkdtj2roi9AMo2069NaQ2ju4uyVY236si2042tfo9P37rhfAiVKkpfEF7w5FbWXKsmjBTIf8vsoU
k4lKiAXGScCiyXpjmiccIq+/4/JISwZaiZOAXEAeq+m6Z6LcKW1QaYlgQ26EiFGRr77VhXxZ+NC4
hE27TYzOu4oH8L54iN5vJvNsiQiXpNAJAgdXmIrcZsTbeiGC+f76201xyqZl/H+cD58yKe3sU9nN
JN3kKvmMBGB2rFPR6AhGbJ8PY20By8wfXe5gxQntcuZM5wWxi5xbbD3zSlzukGKVVBh7tHi2tGcc
VGN42C8feuWTjHD8GlmW6i1W+cfUdXOo1cYkcSTCInuxke/UHgkodqouyM/11uMJF5ND3xJpSGXh
bw9LVzDhBXbWpI+JRuNVsoK9K8hnpVtOgKJ8uFE3cblKMvm6t0w9n81um5NEreh3hyyWFNynRib8
ABJjQmMyifEw+8IYoojBB6NN07Xql6cjNYDLAbKLAO3RV98tiQffX6A7WeTrdqxG12jxbS+K9GiH
FtijrkdDba3Xz2hZeZObTu9gVlKSDGaXqEtlgNYryPVujxNZjhRTyGiZ/B8t7xor4TRjTxJIn6oJ
EQypskx1EtJCSuQHAY+0Grw3bmOi+UQh97FYWE6SU4Hsd4qs3CyVotDi//hID41e2RlwQ0Sh8XpU
T1dPOkBwqqBn7OVmau6EgXARBaNtEx7O7R6m99iRf/rbed2Q5XNHAfkq2O1EsdImmaSA+sYSviJe
r1pYnh97by7gFBXwDGj55x04bHBiCjLSnlKnkyrwThxzG8yyOjxMnDa20dEhWlffmewMH3IeG5BH
Wik+M2Gq8kXbhlCVV6LOc9LDqsPkZ6iTxK+JQbwKCznoVCW95RZt1uOxFmvPf6Mgm9xDo+XLSGfl
WUBybSGXIT5m0q4pVry/1ihjbiD+CPD9wKRtOb+RdBwblDWEMLGwcRjcGGoaVupuprZ/N8NkJjW/
R3kQq9KGqmLlwFs9NMX9C7SWP7xFrpk3AbSFRrf0bIZWiq1K/dZVSvzkcqJho8Pc9AokJfv34gL1
hJ7zhZ+zylbtDK6nEn3v+JplZXxcmPYX5pe4grZK7V20Xic/eL1yO0GE7d7hkQ4hbHQV1cA9IPtN
mYOSMj73Ja4aeeaODW0wlw1I9TojNhlpDbLFzBK/Oxup1db3hU9K8HFe0DcHva21NWkFKkg9jfUc
RdfxtB5W3q33fGPrrMrleXUtziUy//N30HAfCQaoo8+OwS5FEW1Tt6D89LmHR8m4BRWxZVugqZmL
ugK36RoDOJ9ubM9hKKb00tPR9pBk1tJIqN/VLJGWMtUShB1FwcvEeXJl8/o0aybC4dwqJ9oqbF0b
Fsna9oCcWr1UyrknUM2lhvsVoPwCy4KbWUIEqgcibVDyLIia38+6D2ql9zmKbHIVg1lAyLbjzjM8
UMFP1K3YGiDh8tot0SDOSFkVtewAO9CmNIYR/k5AzKlemC2zcEdDHCUbAAuLR/4PfkYx9eQkZa6D
4GJ5Xp194Qkl6jm5AlYA7MOHTKRNzotitFxyu2PBth/51rjEcykwXvJnpIx8Tv8/3htY6kOAxMIB
K0OOZttQi/yCdwgZlb8YKHEKbFV6zJKwhEfQDN0mAgua93gtO6y2fAT29neJClyDA51qQb6hnPs1
W47JTLKwFKZL12IrAGOj63P9cH1SOWzUAoeGndHwW6ukwy9s5An/9QzP+2qs5tncUyrjJc6CWyx4
jepqZqBx3qefv40ItNaySGgYsbrBgwrwxZs80KEMrjDCUiyA8nJ4kfz53faA3LUsTfs2Geyn2ILj
wVmxS5NS0O1cFpkWPX94HP/Oi2cuPSXJBnDY0BSkkkNDhOVgFTaSiMLu5Hu+zWLyXCZi9vJL+uOg
YmJ4qATb/AHiT9mTug/Njgr2UAbhW3EUVTlZLmNXPM+w8tDIji6ez2R21SU1jrzULSwXnjAWb+VJ
Jqo4IUzd72JUl9yPc/1gi2GzuNhMcbpM56AanH+lXFZ0cXm9KAp/wRK/L08PabFVhJfeByVXWaAv
ehJjvNQGSGtepnGRTAUMxp18wDwoHn1JSc/WS3yDAboeQa38E/op54dCJjvV1zYm2jZz9tHsbrTJ
O638pN1fDAUamQnux3IEiBQC2F2JSgOlsGLskhyGfS2UXtYwsFAzqtm4k1iSzwb3qfRdt6vPXcRd
KnFMMpNp/I+uVgPtBsxZTnqWA4BQDy2ljhRSVmHgue6W9rdVpJ/FiH0Wws2sjlqBI2SolGmzajUE
5oBne3ptY/+mKA7mYw3UEaHLKy+cIWDswFVQmZ6H0EXqvmEdQ5yoiLeeX/izWpw6rGIZuHz3Tc1k
V8YHieKzowg/HDtNwuiqMp+idJI4ta7f6G5QDYxIM92a4JAdogjO6sTZEHF1YDPAW3mnxkjGGRAn
+WQkad44JY+QTX5EMVd0vIQymt9V7zL4dAUD7NB2+ls1o04C+1WkwvYckf4scxYWX2WYkZWXqYR6
onqBC3HT9N815mDhgJYxOVAbpC5z1Sr4JQfcVwU3cl9KE0V7wQcEdfRDX/d1e/4AQl/3guRlOq+q
/Ej6FL89ZSuQPx5XY/fjzYE7i8MykxauGFW+jkNW3+pnGZsPlF8v22P8XP5/pSjMKuKvgD1INE+4
QL+zllXGv8sVYAak8wPkTyoVZaz+3jWWbLRbVT7q1o/RZivB9BddG4LNuo4RfBJSNZnTEugmdFw3
kSBVD47ZvnGt0AIp2JYQHSPqq/m+FtnoK+ajZLmIe0g18nysjBZPZeJSCCtcliBjjBZc1iQZxqKi
kihtA1HzyYJoaK60gFThpjr2l4SuCh1Bhldu4xpKessUJToF/GCHImF0SgG28/vZVXMSREbIXHjV
qn/QFxoCxluQU5zncVb6S2Z6lAU/3AqqNFD70FYzw8cAykY+YWUe0MT6whnR0wLZl9ymtNGQGB+i
nLj1k6v9Ye27yi1ktciNCSenrthsuYcVeZPTo8fte43yw5QkhqiaOY2C3ce56NoujEDPJyr68BlV
9isfoz6onTCAOTq3Rco6Of51orzv+yQy7t5gZwQBqHCLEISHJVyqzYmTUqm/vO2BVtYdmGnruQtz
LOdbOvFrhne29KMPhOS+NNqTZZqRbE15M+gGheevJvet2C4SO2m1zhu13pTN4LPqF6AOeTTk23lx
cYqoysJEvpgjziWFohXH30a/Tsm9Ly+vFZZB/Rv+E1qLRJzjy7OznnjUvjHZErvvJ/DAx2KEFeP6
wL8sPChGCykH3oP+y3vKNYsCxIFSOdc32fd5LFwJhujbG/Hjq4Im1eUDe/+7Rh+ZtJ/Pv0V9QIaT
wi8Fi+64IS3bwRMlB5ly+cRDgQL+Rz5rYsKcwugW80EhrnObProFhH7WjcchLSDQ2yhpA0rlPK9/
QCs/tWnu5cECW3ZOKvVrSiVsI4sQ+K7yc/rYfUcRqFHsjhc7FH+l6fP6z5fm9Bh2PPgfFjVdhb1C
SK8PZYGGEH8r817MMSsfa5p6ev0zpCJtnNA4QmD7hCvPP9SDynwL7p4SPpYg1nlbGZ6+OsB9reKc
Q1+mjVFmbE2yvk/cffrtEoKL2BiUEKhj/DmXPMhzGLTX20zkpIcJwwhwZtdI5RkPBKCo37ibZyxa
pkhXuQoetlJTvnvjdk3lZh6ZCkUknk4A9i/K4sxLbCvpIKp69Toq5y5x0NBLzVNRW+FKBukkRLgz
7CbVr6HSnhETk72dcIlv6jxGcJuM+DwIotsmoZnU4zS8qGu2uOh/TCSW1rrKVqTkpsrp92X0KCPP
2WEUAfzjV+dYky+aIbu0gCy11IdBY0OCSXmyNJo7sK26wq6BsH7vIhgkqkQb3FxIyI0e4TYIiTg9
v3mE0usjdVzJp8+bSs40rEbzvRWZ0i+xC58hhPaXxUXdcqhp7sKrH2b3XS5vjMS0tWYaizRMchxl
+ZZHORxbW1+MFKkbFVFZt0YFhP0ZzviMohRUTWE0/f05F0BW1D4zZGHYg9+s0p2d8IbsjkO4VkCI
X44d+JGCkwuqaJH1Bs9CQYTJLw5QPAn9HfvJgc0yuG2MlXhtloTLigKg4tjMvs0FZI/A7ieS8TUb
Yxw7BAjAh1/Sh+hr6U/4kH0Md/WSy1GqX5hbMXvcEET5XmYj2WhZJmfwmSOYUYQ+IuGbFDRnakCO
nhHY2CXRgo0BwgdMwG6mugUnt0IrZQePwAsTPNrcjuXTtIB8/hPnPTZk8RP34IyoZ8Xno9VHcQik
4UuJab+OM0H+1704txQjNMnN80DUngLBqZlH7AEALiEeA2xJPrp/wyxt9hBpNloqHpZjWyG0KMWf
ivC2JlP5qY3LVvpJ7LUCnOHh5JJR4FJz0L7MvmLa5VN8/SqwyaB08xTxlotEaCq2xYkSHbd0UA1X
2arSganhMbAR2GuIUnlh6AGTD2HhyAMjXumz3+6Cjfwk6ek6w2IKfXG43EDkkn59oUK05gmo/xtQ
cQGPiJJWF2DMIH5l6NA/nOAYKwP2CJ+1vnoc7iFIEDlz1ZghQLDNY6FORyYdAu+4PnM8A73Rxj+r
cHuguKyv3l6r5fMhrn2+axB5cs/mdEmLek2HEpf45WTPRlSPKNu1My8y+S7Uowc9+3oBHIpRGL8y
SQwmh3hxPCcoS+M7OxvijusHYj3go3943skxvrpU2gSB4g4QfWXF9iEpGnQL501mxtTUdOL3tIZr
38YKtMVjWnz8r9XPf5Kx60m26NVck5aWp7qgG3usF0kHBuJcUxbVJJUOEnW6+uTjawed7QBcvkHd
VaBeyeWKrmi+V/8FjwTUhyntFZe2GjMyirUnplHplQcmZGwiXB0/LyGi0r76ATaS2ajKcBsk7sY9
isitTbe2GJ3QQUF9qoNWpEX58tM9SlUgVgUoS2/OZHk/RoAP6PzuvSrrZRVY6a7nus/aj1taDsNV
4IeWJvkDFizmTbmVZAp7k617fU8N2QLm93sVGifZSgMvdz77gcWn0xhn+zilbFppEYy8gtOJOgSx
ZGDmzpeFLVDeAJ8pPRE5d7yxWm7gGWs2dsX+Ummwez8hEhoNBXsHme7WRaKyjQQNE0HtStzNxII0
He8FP9r/Rp2Cq7tAIc5JfZ7Z5d0AVDMSFGVOiPSpmNDmn4TFhxqpUZZHfDVeXF5UaE89gZNEvXGn
770qL2Y+a+RLZ/e2ZIphxLGpk/+3DqHljbmWmWATE+yaK11mnWS0igTE6Hm2im5qNLNavC8R0y+X
Haf7DbQSHKk/BurrngYcSk3zgBa+8iXG5/pjZr8x8tsNQ0w/LSQos2BZnLR8boSRYnrzOxBn0oSH
ebwV6BiRzAsO8c1aYtAkSu11PrXKjw2mtaBqFf8C8IUKIVcKEYKtLLlExwQaQ9O57JGjci7fe561
AsVswom9D7R3/gBPIbLPFH89XjQD7y7PwqdrOxIjF2idZQPPYX0wo7ydutjE3W+BWuoYM/EGzO+P
o+WRAfExVO81ilAF4yqy7lvdjhCsxr4Er1Zy9VS5m0GYHGMjvHO0taF7OF0/40BHTLW6Ajy29LTH
kv8e7bRnqgw6xXajxGW5dPEKGEGVuGrsNI8cr9SAxBAq5z48qw7yTIA9LSFN87RRRzm+6IxDwNcI
aHhyn632R3OD5bKabDNFWWlN0o4iussDgupc5UX8BLgAUfcnBgtNJpOSzgzlRZA5+c2DBxiconwn
c/sV4lTqm9KFKjelRGAWKyssf5Rqgx3UvIomImbOV5zwwDZu3Q4iJb7+GRFvKjzPVX0ynOrnzx02
qq3mNqnE1HNmb6pgmzhMBeRxyjEUIddUhosjmVW9j/b7CGTdQVz0uO1spAXsEQn70y3rEWB56sbU
Z0tLLyJId+lC2QvzGxdhe+SpdarZGMJ4fEUFfXs4DuOF9aO+v09d/+Xcd/15jOvp28SJ92kdxmuc
D+WxlUgQLBms0z3+gkiGG4f5r79jhho1CwqUG6nf0GG3XTbLg6UmcOcpEpxG5Xtibb4F/Klecudm
enC/jZ0JLDOUlEpTjjY69rbAHo6RNsoTvscxp5sSof82vwrHpS4OLuT8Y8jxJF6WPi7cqR7xpvt7
d8g7g2X0WZfSJnIx2679iaBo63ofEFTjYeQSxFRPCtEz/pxRxlPMtI2tiHlIQfuFlAtlBid/59Dr
O0AvwVoPiwc/Q1jVQPhhZX3fPkAtn6qlxa6p6TT69vbz58lLZ0lBJz1QSLiLn+qPt5L9iUIdv4cM
g1a8QStspj3ejumGFrbeW1z/58prwJbbyUmDvLU0a+IXOGeW9N4O7Uc6VYK8jAmoP+1aQYYYq4pg
3sWCBwJ0M8mG3RISGr91i1odW/H3nV3OnX/V/vFZ18Fz43RKk4OO8JNvi0HYZHL4VvqMeucryDnQ
FFoUGWs4jRnsHgmHyOGGJEAwuN9xZtsbmAy47oLJ8FyVK6lZgstmUNfpI+uedyl9sYlIc151wJ5f
FaXDkr8gbqsQuUCm38ezpreC45O+NhHXuj/0z7MiFWEWHlQwgr1Cc8xoasc5qvISS7KhCkb5LUnH
MunZWO0scNKFv/bKxXYSMgf5CcY3yqW3sGOwTVkgzsSCC9r5VCU4BNojtg5p6qVo8EhNt32dF0du
AW2r7Ldmo/aMrHFrUe+YtTF0Sy/tnbs4FA7JS7IAkOUKOWd5/LILkjK/UGIkUQnvRjTQ7LJiRxDX
2myJIO3K0EglUoBR4bbDQE7pRoujjB3vzh/+xgT+53O+/dthSyZcBinRRIFTZm9uC40n2im47RRB
H1k5hvQUDo2H5iyPxGjeCBz5dZ2bg7Pt3J8lCHc2UoJYxjDEGYkswLRjdjhd2CWVs3WgseaBB1Qv
VUw0fBqxiK0p9kXmwXP1EAX44lMrw8CnYj4kOuMHkJepihccqg05IwiB9IQ0HjRAHDwfBdTzO6ff
vH/2mRwHWudV1P41TjPvHNn+eR+5XIe0eL8GABnBAkafeQtg9n+2ztC7nYkFt+m1MpehNfBVaeDK
CsGn45CXJZ4AOnzX36TZfaNHvhcJb14DBBE4HQvBanvPlJcDSLTOzXpBS3g4ZpS/4/QygJKoVqKt
RqEtqoydCwE3TYYpaKu9kWfmUMFA1VQDmUDuX6OR57fUGQ95fMOT3LblYZA65JcalJFiv2mHpiti
OPsIPG1guy6/d6LXTWQuO7iCFfPMh8fhL/IBBoFG8c9hdL4TineDMSGQyixhHx1NYtrwHIOHWhWi
5Q7RoQgbFfBy7mJ8OcCWl5UTH4ugsV/BO7+jdXiE9nuE+mlS1T+0ifV32Q5F2Xv5H0ZIdfT4q8CU
1XeyOE8ggpwXbdf652K7RSbX3Nmj93tgXUxF+sntZBuHnQzKVBHUINaUn4i1yNtHwRubJV2XKBez
XE4pbEy631FldlxAnFbYhdItCZbe/jQEezi2b5iSsLOzLdiZKOb7D+I4yKWBaAsz9S8hLcORwpC8
5z1uEZTOBdYXDXVt6ieq2o9HCnv5TVyLG29e/keQdx043jcbtFA2NNRPbgBW6xVRHUcy95YigJFb
DPd74djO1HiqruM84VLj5ZVhwB9H4twK4E5xv0NeNbt7kiu93+S61D+a/MIBfq8HuIVZGWCXSFHK
Ll8wt0pbRHXO0yiFdWZsEtJgEhcugZ8xVHGq+NljlwD7KlopDQz+svITS8EAHZ6lYM2FVTh1Yf4D
w2XsKQZhV+pPcsiVB7l7+PeXsS4kWGleurFN/Lq+G0NWlh21mE6nOdmYgW2Bp9T0C6VPq30VSsAL
L9jLilxuCNBYoyBwak4ZB9B5CanysKBoDeEHeaPcepuR7ZupGtShBhWUOsPUqsCTXUnvglJo6RU/
+T+1hHoqQLiJhqsv/QtG3udu6kORnWsYoy0cMB3PZYOigrT6ZrUd/i+5syjOaJxVYPnJMNKXtSsK
jsy7Dkfs8YYSYt2nxVW/yxIsG8fODRCMnbXbk/h6YEbY0GwVULsd+aG3wR4wxqecUi2UsW+EETWl
xkxTsgJuJBbWFnrSSN+jGM08HwfiVy59GgjFnlLpDZ9qecWdT3OcfyVVDRG39ZVal7g0MEsJt2Gn
szeMTLzsxi59ojPunNGQTKZZdcxqCc65J1xFCfjATWpevJympYJlnlxuk6b+Xz/GKbZEN2btg8us
CTUXIYx0yV6rO2A7+lpWAwdRcMejfIsgKgV0FPeLA6LMkEn0KrbseGh0We0Mvu5PXeUMzblVT2sg
BSKiOAnbcdgwtKJxdQfwdAUeBRT4qNutsJzdENjuuGNPsysTgPIx5WChRG0QG5nEFqVNIgKstytm
maya5k/ZCr5rGIHSLU6GL8Lxvv3rSvPmPyFCBSkotug1Tk9unhJx7Kgz2AGiFu8GtexCb+gRK2Jv
Vi7O+YeL4601dRz/eZJOQ2Puv6zZH7U5hXk2P/YScFo9V+ik+q8OarhxyANW292YyMHEZBoROJRL
jbGbSZ6SliM8T8EO+KQHZ1UmARS22UN6e+zY9AiquUEr1Vpkf6zNDTSOlxPwIjnCYc8375+TSVqN
v8RbkJzOTAFhdj255G0kpJtDZMiAFAX5Fj/z9hNnGOPlPewfOWRfe8JhfRDU4dqYlsglcWUKmbbN
aGKSNRobvkB/0a0BUR57c39V5rDiezlwXHZj6AKO1IPVkgUSculgLlj3QAtculEFAqyv0novyj4G
uKx8GeK2C97EB6gqZXsvYtlWrT1Lp8V6zMbSSuL3J3cW7N29ESSbBdWt6RapMKwU7rjRQUzo7tLJ
Gu2gdE571Yjr5kJPgRnLiDbAzZA09liRa8R2qHjz1c7C/sqhXWZ8AfK5mlPXOBxS/xv527h4Y232
NO6IDfm/JenY3gAfwtGeQ/Esp0foAYuvIW4knsYdWypgt+QEnvXSym0/QBliEFZw7cDJRymppOM+
zStAPncy55f7lKotT5i4ucG074qTmV0uz50ChnyJfo54O5wtMH197SSpOaxD0CVEnOrwelWYj5gS
bPuHhReAIbOlqRd12Roz0l3f0dPpcjD1dMRHLFPeh3H/TlLKNKpJnSLFONI19/B1Pjc4ZkwRDoyg
yGi72CF2Vq+bCVoNWaNJl1Sr0qQC/lgMxo2n6CulwmZrxC2/HxvJU5WovKjbyLwafisVeA9TkrkC
gTk8fwy+mGve4Y6LD/OZmb+R+PSCyws16hSET60ntChNbXpNlWVLUZhwoOxUW9hQMSaAZyD7KX2H
5uJ50QWRKEUg5CQRkBbB/K+y7i3P+PJjx+yYdAqbfVoy7zHGwBJs9btle8wM2+bYnB0rp3fU/w5B
G+GRk3/b0JyczJy8JTm6OhuZ6ksM+o3xQTAgpzCUGK6ezB8VlcLkBZ42Er4lJXBuctJV7IALsyRr
kWdfH9J+T+NVY7+DXVe+1Cjp94r9lxpq0QSetT8+DZ4hd6wvX7kTK2HdujpfzZKTbVqeiESRhd8a
I6PDgaeEXd4FhEyuDt0lZTOA2LEAyX05BSPBQzgfsHWlMsB/JSJX0VIITgzsctOTjXYkCe6TVonw
m+2Ldgg4cPOh8ogsOFTG6Zc9e6VY5obQSnGnCCEBcdVKmDgsSi7sJliKbQK2IS2GfOwGQHBvwh7g
zxgHZvJMxsb++BvK5QWQvPhk5duSyLSyMmh8BhUnTjanIbQCx5EKQ0udIHrtbpSm6lCXPJwCBhj+
CiJF1fLaniZ2F9CrMOAkEOdOhP1ayfvr3PX2BXIt3aOaEq2Idy4f3DwszosUSd1sJ6yvBWwCHMml
0c2Ux8rMxHaITa1wcS74mTKvycnFoDd6siZuUk91PyK+hd1hdaTWHHz8CUeuO989OdhJk4ufGOIz
yqqGuNAb/HwRXzSoGbAuHYBApmdWw1RBCQHDZfOBNlNJyAYtTD3gtFQT720Q58RhhiB3mOy0Z9Yi
+1fdSFj8Sv7RgId5FppqypW3r6lMv8KHC2thvTyNNUD8/cKV5mv/3no5QWZw6eistGq1HqkiTs2p
3JAgMEXrivc3MnWyZ/cW9IjZpF5Lf3a8ujZ/6nud7LLYkK+5RHQBdvJ5651ZoJUelazUBqktZtlX
z0b6PZhS1mHGv42g6TS1dbBR71epJiYqp4qMQVZcIBnlS69VCAAIEyxwFyS3BzhczUC2CdBmt1h9
s/JfNDorvRwFvRV0+UBgGPPDUS+kkm6chP1s1gni7tUk7s21QTkPBQUXRLmDp1RjqIZjvkyYPdyl
YhHOOTRxKBKZ/A4gRdbGUq7Y1EqJ0FQ3JEPC8Sxtw2RzL4DLSSwadbTilc/02AxA2UBoueiFE/O7
kagfEv60ygvEZzq3rJpJfpA9VkSedRqaE5JAHzX+duYEzrW/rucqg2E+QJiFF7+uOuQ8LkVT7T2K
HeRyHvQKw2DctvzAhS0ljRDTKreVhyiAeqG4+ac8zcEtwlB8YIQy6HN0HuFTom8WoZjqEYsOwLyF
IUrhbeqV4TSd3NS3p6YtkJrHdxtkZN32UIV9ZvozaYFUwkOEfRxgQiEXn709opMsz6wrRIP9MyYm
6YTVCsL5XruAvXsLcBV5i5JeUBeBY+KZeXepBEdjq0VBT3A0/a6x6C/RrDTfxScVhqscncUpOaIB
4tthGgxuler6W2k4IWex+9g1yBYaKNf8O3F/P79kRF0RtsLQA8UyeOzvX0E+n4ZBetnuMuS+vNXw
YaNHIHE5NR/Z+jXId0/SgO0T6N428y2wfxTyZI6gP0ZakYw4qpApxUZyrZ/gYxppSYeZ392jKgzN
Osz8dNo+/MGF04pAYAWK1yqVtikGwfY8k9LiYcc0yJGaJoqkMahqGgmbszedl6r1cFw058wjt5JC
VIQ87shNw4dtiYlzzcv6mXuwilL/91Px3uwwmbvIvH/aMmL3Jnasj6WIUYF6V6Fja+b/9GKejJ+o
VxmAP4IqPl9bMUyZdtIbNkO4LqrP6J701yKWx4xQXMt3WIZ5rRl2bmFAWa2mDkzgUQYEJZYbDIa1
/f2KKI8JqnlWasj8vO3qNV7Pnbi/gKnZO/CGWhDS6WbGzQOIMSACNewRwrHB79e2LiNQ5w/XzlG6
yWS//BwcWjmcILrTnKxkaiq9g9CHJ+VTt/Y2VnI10GTgegT/nkfwidhLl2uWp+8906l8BbsB7Ahz
TuuwKAHsgjbRvB8ouEPNW0/fRl5kULC+Imm8qH1brV9W56CiiWtNwVFQQPSqkDHbCci+TWZ6wwf+
HrT0A6CcVpYtl9LEmWCOXrQljpUMETTUKRCPNZcYECwgkORUpwqWH/zBbLwZ9/pHHlBXoag/M/34
n1O9Y8HNoClJRGK1hCcaNYsJNUDPIfty1GSTqyazZnTb9ae7c01CJthOlmV1E6DNTDqTNLCX7kAi
zCQXN4WfUj+MY3wyHK8ihbim9BScGv/CrgZ2S0zROBKAkeULjNxoTgQ2psAKX3eQz/9BGcCGG1eh
Z1klrdGLTfWQi2JiN5wQDaAe+gJghrKB7FOLv+V5w6T9sIVSfYT6pL9LLBaRm50hKLRCQ28DPlXD
cv7+x0nMP134yiX0BpSVcTxoH9FS6saeaWRH7mxKisuTg3H1DH2LYXMhrSJaKJEivYwZaXIrU5Fl
XGvZKMtQqqAAEDXO3Xa7xmLcEWVZkCC81KU/RKrNbfX1a8SJZUUZaImyZHdS7sng+lKif5F67OEG
J6IwKjP0vEdhqyrCRoAMVAjkMHMy5Iw4KvVlKX6cbcQtiW+nAXrsLl5/Sr+1QIaaAIZxit3OBU47
iAbueEeQcs+h5yNA2Xgtk4P/oBXeP0d1Pv01fMSG3GsqIFlOoTGJdwaBBc6HFOZVpoa2cpBZP6Gt
iAkJxdiEoDRYPGwSsEJduwlStFgwDEZ/SdJTfmWgPzSsSHovjjexGNYvmNlJ/WA3jo3pjmuAXM5l
U+HmygysidHa7H6bCiSBTiCDQHGXuwywBi+KfBTqQW9rxXU4K9kknonJ58UINX9vMTNIMkKhsl5o
H3eIt/0LS+o1c05GJTyRUVS08iYeMMFxbom4lbfaExgwbdmWdnnCZvVDArNWImr157qMSsjrKObS
roz4cu2qw0LvGb1/kz/TyYSPhAy2ennrMdOR8HpbY235XkC+bJtkqNno1X682XBGhRJTeNPA8Xqx
EGJzc0Hc3YsaNae8XhxX99iNDAzWYwxziwwXqqd6CSch54krL1gKX9pshob6nO3b/y1jy7tRf5B8
KxW3KyUXBN+bts1jF6AQuyMuAlk9lBt9yB1X4cwIyN72DobRugv+s8Rlvi4b3M0tgHlqfyHsFxtR
G45U0xEaU8zDiJuGdObWSkTFUvzZ27F4q+UkW11cnlqRp4UAC0o2r5TfVRfvPLLWmM/6QSQNXqnl
QGWZMxYRlDgW8+TL0bcPCibxH5CttUHXbs40QEgZFeUe1zn3nvi7HatVPFU/x1MoJyVN9i2SLOhz
Dp5X7FazASEXNdvO+Ah6eKQ1tRMgJxrIYY3XEijtJEcyX2bJ/n9V5E0iAEX431tCo+90HPYzMPU7
5e2JuZdujIIlOJmgM6q0SSynDIuOOf6IlfS/zpLgQK1d5NSqqCODRHPcCQGK2OtUh1VtodkkXssp
mpB+VF7pwKlXarVmrGFBEL/2QSv7dirfH6p6zqrQv6nofqY+YnNPFDyIg+8bUFMyAPV2PAOIyF7U
e3SdSlQ46PF6a5HxEixmvugmhWyybRjwE8FSA9aDVeFXZcyNe7+1XEY3AY73Vdyy02YKWCQGaT4v
mjs+24MiWz9vhXg6Z6+F6DCofM3DRZYQhoPJRllxMbzaZ22leXJFnTE0mCZFb8czKV2DrS+kl+EM
1a6QJg9rQWWRgP02cuji+gvgcVYnUMfxMONbwSAKBG+uR1OVhVLak4Pz2WqASmkYxZ2joTjt0OWH
7QaE6xvrP57wpEIBnL9jf4Lgpb5wWTp6SaWti2R5h2MxAVF1SdueeauFyE0/HIeftiIotE5sC54Y
1UFN+VvXKwhEg+Qcx69/OiXqeHY577enI+Fz3fzsDDk1p2clu5qkQ484SpDY/wBEqKccj+yQtEo7
1TpJsZORAjsXre8luon4Hkk/gfIth05lxv83HTN1meNl3yfBaWAn2AxOSatFklDT4qmrUGxFRe8Q
bv67Ng34B0Drir7GhGVOu44Drnn7+Kgn0KfpnCAXNGTSPHdg5GXEQL9ddV2HGFP1EXsCDbE8nFjk
A2z6qAJTA5urgI+dqk/wISY3NZutxCiYovFB+AOwhOcsybVNJHh7WuHhvsJg1pmmnJ+JD46wmOqY
29vIbmkGdNVPD3jngT2XZhZR7/30uJm3FsqR4UMeWZlMu+qRICXfvzc5od9ZGnF8vqRC0yfVnsy6
885QJ/DQFVON0HXwSlf9cLQUtJYn8BDCxI3tow7+4bnFjHrz59YHfJQKd7+nFEiGJlZBAu9qRTiS
oHZgWigdkRi776fMiTx3ZefGfCVL0vbQk9Oh/IE/UtotqA+gq1T3/dS9Ud2Tn7oc1eVbUytwB+08
bgcTp1QxfECxMV4FFIFQdGhimNhG1gRPvp24EBK3QgNZ1mP4bVt3EYBay9T74TpqXYmyEt0P6VCf
Z7FbW3v40nMSDfP/eOgCsw1R9NDuVOQ5vtVnyBTGeVmrwcmqf9AAEJjbQI344mnrmcbZOZqV9mb9
MwDm2FoSNHijDl7ueckMZcCkMuxmXIhuT6yIKUVdOMyFLqkN1QWGSTCgZdsyjFBr9g05P30MoHRu
ynrPko87m94lHolVBk/E6mK1oFhyIm+sfZMf2FiyO1vSkzaVS6OvHRHD51Ui1klgYOaLtceSktT0
uB4eQBibHKa0Jxb54jlBp/P7oY8Y8uQ9O/BkpHpG1eUu2hH/Wghn3X9IHwWSuMNAxvIbpTUr3S6a
kQfUxPR2tklg4gNpnPDuwc/vILr5aRCDid2pA7PIln1SRyzMvd6dYceZ6jSChm7XoJvYq25AaD+i
xcytl0dMswGrPwd2/FKydCAfYIMyRmN4GgCp36IiFYaTkf34EcpYiauEV9/Hoszda2VK9fbPXsFh
GIdflRIDunVk4toKiVKcNwfk9Oeok+pULIS46goGNjw8A40wnr654MyQJ2B0NBIXFP7Yte/9FPKT
bE3LckcwsHBGr7FwhPceRI82pHWr4c4WcQJOr7V5Og/B0N8GouWZMffQFq6lw7CwTMXAUuE/15TH
N7iV5FIDIzo6f1Ih0JreXI7j5vuovWBh5aYiHXPj015yPCckGRRunKeYn2iNLsmGg19M+AGPphCx
2wLbSH+Cay3YnZ8xrc61zKlyJEcZ0cx4GzRLLDc9AjrjmJVyiXnwEMrCodxEiMA2JL8GuEXbUFSX
Tp14aM8z0feLaKoreWERKyXboSWbTuLSc7of7aekXu7Q59o3q1EOM1ibaeypKhru0Su3fqRFJn6L
nQ7j5UTLRudkVUcgMkuMs0BNRIb1ExrU9H+mUhbaTNfnoXMtsm0jaaFUO+wY0ZijvK/HJ88k0Wmi
uxSujTF3Qz0WXGxERCkC9iYPtmKrx9RJhaR3tgsKKVEfPY46D2vDmYfd943AeuT+B0wUE0w/4Rhm
TzHSFIgpJwh68t4Jq1z8J4O0+gCEzl99pCOKf4agwOzZy34PZBmy4JpebvgITV1LIr5rMSFz7Dea
X1l8P3XwMhsQdi46t4SrzjP7JzXqIdhb8S7l90wxdJBw+U7cxHdUZ/+AgRU4FafJc3lzLoTBQM54
P3+X0V5KPyhRccEaM231f7fBHA8ED4EqAWxSmANWvvCDQQsYlEPDxDZ5//X1W9KJN2yHJHhGPttr
lzIqvZNvMYjdUOSxidFP2HZYoGy/f4KR84pIphw0OZ76Ua557klpYmqwTxMuQfKV+I3QBlhVGNlh
84wY4uBC9rKsnwh5fGR00fo4EueGld4gSqVbPde5BuiGGRah1GtkIEtp2GAj/TdQu901rdgGGGJw
eL4S/k+iba2BTzUJs95o1KrM7C9x5xUp5McFyFrvXjfJ806sMswpg2+JiWyAN7sjykV3Aqnkb6R/
akcp2YWAz33cBjcNTqEGsER0ZtMDfeK7KSrxa3Bt17e9JoIrZITYgk1hKQ7BUFJ2K42ItwP8S1En
LTVWgmFxmjQ1aBkP2Gn145MVHl+e8hgtBIMVC8YLZ/E97d0jJf4/Ezegvd7XxWuScRMaB0IjLPzk
3JMk0d6qOkSxjlNTPIXle5RiUWgCvoYUUAtRcGzqvHPbYqZaEo7QYN8pj8LObEKbZndXeUWsRVAu
F77Dawz2rEm9mfA/TmpBYkNJIRmkwsFyl6gr+Mx9k0CuT/H/Hr83Z3fVSTwcfSj2bTBV1fo2K8qv
/j/pU2GE18Y7DyRxB0JUmTS9TKLEolftaoidWIHioMcG11z/RrKXivir3L5XpF1fFlXJRApgwYEU
zxbO3fP0mmED7Ac9lgMa2cwfnKo/mc3TMQrmjAKvUjKp00a6eMWNJ+FUrDWN5O3RDP6oeQ1rJXDo
flwt/QuOwoyCDRFuG28Merb6dE9FuBNcikmCh+BSdNtXi+JvHeWNoslPVV4yRfMphaC25qI4xhla
6d9uLQBBcewkVPAi9v22l8g9WC83+MQKOIBeJ79WSVLA6UgueNuEHXwEs3UbKwvOcVVYhMv5DGaM
dKXVfkeHKyGC4SCfsD0bq1jvjEUjNhPuVVIrXZqUjOYedSMlxhCNn+LzvizW7mgiuqbEUwonesZP
t5RafmrORe2OIxNgviX7g3oEydW7pQ/YfLSbmCOY1Tyob0pzqKz9vCnpOPPlbd1zT1Ot4Yg+7iZs
llD1YlndRKBcFkFktux2tL4cQq+5dRrKhajaiDU64WxpBADNi0hNKYTpYT84ew+MzEsn6+WU4l83
GTgNtHq8SWn1eKJytWSPFsfhH+YljZW1MpALws17RcIZuI2YdLqEHG5Cc9WcF5veTzBK8OQvnZ7Y
cb8ruPS2SgKKK9ZZjiw+vHy+6Hm/HKEMNplcZb4DlqWn1HjjFk/1q3KvT6vZQmELh8eMi3z1FEFp
GvLYybHo0czQ3KU9oRKLjYz5lDpUk/iI10Rjny7KAihm1wExUobLY26EDlFU0tLr9NEi+xcHsY6e
qLbsKsWEZ3BuzIMDjOjmFGwHNeGRTgEmh5Qh4jh61nlcbHLlx1+9k8ut4h2HegFRRKV1Groc0/j0
OMDYvlYDuxr2c5c1q2mclfcANM6RrTRLiAj9UR6o2k/q0nAFb59zZEi6FWr751aR3JArMrWYJpGw
y0JIUiDTWa1xAPpyKbPVxC6K3tyLqOAhZjX3UWYS1z/M4DdD8KoPbgp+GUKniJgbBSqnk7dwqWNl
hC8L8BBAYN07Gfpb8dQvTZauptd7HoPA8lFkrAYnP142KpSTHPKiDK8ocXhGK8vviTiwbzUyI2Iq
Mvm4QS0dk2lxex4F95XJOOt14iP95UE4fIgl8DV7f3h2Snf8XfgPfqW87Qn6bJNT2yP45zZaMa4X
S/vrZvndortVlD0i257dEll35XxpacgQPH3Fp+hW6TllH2/Vs9aREEgIGEDbmOmH4OHSOLd/bZa1
OsciXRXWwdkT/HpTA1dZ4X50TMB2isXkvlj8dWkUdyNfN5DketZngfbavHMY19DZohDcg+ayQxt8
s4lmzfwiih+LdWl9nQHsryWhc9ZvYgeFmafyvO9JAqTuT/+xn0DhLxcUiccrJpcWer+EQ830vCGH
mocxQrtEzxYUWM7TtlKfSzJlU+/Q9XouM+gFH5yXU/V3N1vfRXhKi8OjzVDCdqNcjVO1SOgsriwF
0sdWp4x9qzxGUyCEp+Yzbya5joFCDsJil+0vEKTBeqdmQg8AaBvTRlerV3a9P1FnSzi8U/AZLzS0
ZSJPjs8p2Royh96RrB9absovIprFB3+Dpqbo5ugZTIxA2SUIpGyQqnYA+ZR1WO6VwgmWlaXeY3cU
1UZ2XJVW/2CnAfQ36I8f1vl48O4TVSnH+Kj7SBVfqNjh3/erdmQRA2X3/HbrehhhfyxsBvuF6l0k
9eEvDqzhfZFOQ6YJdXumuJSoDEK832d6Qx4hqnIPgbysWpDOCk1eAgDbIMifAdKaANraYrm6k8P5
D56bMGT/wzPi8/t4uE/ktFd3r9fXSOoz+jD7s3VA2NozbcT+JC+5ya6bj2D8N+X9AYlPiWUmCGPS
pKBaOCX+tJARWLyESBYmZmvxNHwD8RD6J6wpPrJwZDKDjLl9PbjsdKKQeDV09quMVwgHVbAoWc97
JM4JmmD38wcPJ+4fEqG1VJ/gnxjKXLN5c9OhhfkuZRtllDp/mkqmVLYyShxwA2j9af7+rfHoJ4mC
U0axMBpFHgkjI10ww+wevwelTJAWxKV36acYE7rQUaR6IAGVc9dDkxEBbjS6+dTsjgAuyQv93yDT
VFltKxUeFrkMfrlhsrqs8ftbJ/XhrHSGiArvIWsCaf5QnQSOwNG6p3q4uC7HiUWvvGjfq/p9nI36
v0mT6gQ1TQ2x+7OWLu5F2/YHvKy3ZmP/EmzAzeGxXA9j0DoJ/KR9cyK1eCU09Ds9RsFogZ1EHPpv
eM1JSvcMK/CcR5x+sTDkKGu56Tfwhf487PBVfYys1qvK6LN+RDHWe99q2/SgjQq/F0kckaNLcKpU
OA06eRhuRISG5x0WxAExihYqdKLeK814bDf0TIwKwYUfSDgB+3W/89OR/2s9D9YXZ02FBCSz+dYm
84jK4/Ds1Ld1artkd8ubZF/o3lOflEIbdP9qY8z+UxQyU+VQL1wPdAKDwRQ01WAOM9nwx8dw5zB7
V1joJRJv6M/AkZ/gyuyY20ugryW84ufK9VlCg138M2o3QlHx+fXFLLbOLls8PFGLD7NFK8TUasIV
JGDxvVzj5xucuetvgO1Mhz76zehd2L35bc0a+UXCI6elfZaIJYuepHUjxyMdngeYCZvJ64CqRuYb
WZlmFyFWaoKGTBO2u937PX5o3W0x4iGk1nwOve9XJK1N0WgY7AgzY2KrG8oAWMaNhXDFVrvCyz8z
ttA25aeE/sGcZlj3apUfdl90A67NH46sxaw7FxfsjBGKM2dvtw8vLMJwvhAvOCWyC5WSZ93hwR5Q
3qwen0X2CCpKMVOdHUx9iAVnR0hHKjP/aen86eJvJiM3IDfYlCzxjxeN9Gdx9wt2Bsjg0/ciyzKb
jS8rOmmo4LYzr0JZcvMvbm+x/8V+41D+Ht5Sx0/AxNt9OsoJXx2MkDZpKsQKO0fhLndsbCMTAecJ
EU1u8wSyCn8brA9RXHafc15IN6F9onLoXsWfJOP6MXC3Z/N3kXFJadXQj7SPAK39eByApH6AO7sS
yC5bnEWpIdvdgR1i6/oQfh7vt2XUXT8sVfA0lEtdXBKm6FXJ/YA0gpTCktVz+Uw1vj22k62GDECu
BtRRl/23kYM8APZ2dQAb1uzNwTKQK0++2O0jBqw7W+mFOQlkKJnsUQOuYjvSg4xTMPVmQC502sp1
amzxoo1E9/dTTyjsK7SNUfjWpKRRJ+2dxbjYfkgXpte/3QYUvpHpBB0fM14plpNVYLEhMpzJsWzj
J9XwQq3NVoPexc8arP1v7nCR4aG+XMP2nkYRsPbsRlrvvGOvay56gU0BXvFhuQXC+K4moF5wh5rR
WHoAq50rNZfNDxakWGd/3Q4lPAIfwAj+Oyr3HuE5pETcnoPPDwiix+vxaZ0Gs2J2pqUSwD4mKnrK
Uz+OR35ICVUSo053XSf8CMtrnoh0GM7ebY5juSZDNq30jQfaBb0QTlTZShdj/D4amS0aqRaCDtBD
rl6cGy67fTauhfbDgGh+6gsVWEB8cmhaswyy4gtdDvB7PCSQElYXad5KEy7v+Gfcys6jImVhRtxm
aPpK8iWiLCCDPv7eEqv3jhhuwq1epFnUFqO6lxmJYb1IvvCH5tSAV3+zah0KBpxPETOt2jT7WjDi
Lw0NFv14PWW1AwpYURZlBcPjzEY7xNSyHd4qs6VJ8ovbRe1BJmSxn6sAGd2sDAkxPsHv0mtOr+mE
E+OafEHKIZQYDcNBnI7WVmHIjDfTJ1FMwmnlerqmx7nZOaxkcTn5SFDSbTN3MtEIaNEYaAII1u6+
36s/GNOHdU4Kj+8qRkjzdoE16tSMjjtbL5Ii+ZE+QYavU9MMd4mTJg6ARXrW5eaaPt/jJy5wQzIQ
h5V49ABcnO1RbZdm/RGgtTQjIcjoZ3aKoheFWBo8fuQKY0S7Hq+mwKUzECazUZ+L/4dcHxgZVJAD
cECblx+revSZjlKUU8+zdvFhhVJi4sy/nx0skNWAqwf0TjYMU4V7OMUnT6eVH/prtnIehqw7+uIq
kHXapt5g58ULfia7DV19YHyVNLyafnPejdZWGPXI79lmSZALYh/CxQv9QqNiYtUGpOjhy5rK07WU
wa5bmvzBnahgPcH08CWue+GXxQJ8p+f4C+fcTrZJzmOGkTbVy+YbZBh1Bt2d4a/kA5qSK5p0fjtZ
tA8aqdMUFXFVJoLiRZzqBz3pvZMrc4DU5bIPBzpkDldyl4F+SFRZ2Y735HAZnsm0TgymIDzxHRta
LWvHERpHGl0NTJfmJvGDdXSZJidhgSm3feVaeMHv+2oi1I2yJ05fCYi0Gsevh1TDOj0vFFvSXRjh
vlvyh/JcXWZT5hrDzGX3vMlqu2KUyUrdwbPqliVLtyfRcYIia/UKq8J8hCvb7BZMfyCu00KRIwJH
IYnQCHrSqeVsBi7Dir0YGxdr8r+KsMV6TlONkvxhZUxFiNiGmvcjQonajXwnQVgrDdIBdJmY38rV
CwrXzdPId3co69sy7FDNbeTvRKt25zCHMo+qraidSE+50MXr2u8/zOv//P50v+UNyb+lEV1geknI
IcqFteim9EuQduOZx6DpLdZMUi2Rrum6v1Rrxl6vaNA2KzKJKhaM8XWdgSbS4tcm0plS5O/RZXI3
uJ0hQFD2sn/SJIlx//SKwfnPdhetTvtE9R95ZhHLUKjkxvwhoVS4mKziGOwi3q+Y8qc11vC5g2T7
dPUyJI1xWWHkj5UaazJLcDn1g5391VrjRNuMarjV2YqGAf/ZiuzlsP2BwFY5VWOV1ScX12xsccB5
AhNtQBFnJhihCj2Tv/QaYU6+A3hixisitxvT6L6Mpoq3TAfoGccbvUgNa3m3q/R0OFycow0NsvxY
dyAuy87pYJqFq7W/fnFurCFItARyMBQvFZ05M782LV3qoNJn44f/BWO9WwDNJuNK1y3BJLy32Aha
GksN+a068Nq8Lo2gwLkuPheEs2XNB8waLus0B/jg6Tl83/5Om7TJG3nDwjyG+QDao0o5UGDzwnsd
GB1d7mW+mdLUV49mARZmUppCZKf77Iw+s9wKmp65ci/ChLcfxmZ8CPtK5WqvXl27Wj3gmEDwCHLi
k/YD/T+yneaw7e8/vwG7yMme+5rAPcYd0cpaZKENGL9dIhFImYaEp0R7Dj7fMEv/aFVgsZdG2+DW
ta9lPjBRlvAoKrXqm9WuAHdvZjHu7EbCYALEJHVUU5IeQWvUHaWbbWizWwHZutf7jr+H0VWLRi+h
8UI1T2pbOxjiiYxN/xgc2MDi4tTQccPYk18jdPA8bD+3/+JkSX9fqPW++HSCTRZ9qCWGdLXi0bn4
UPJYfkWv9buuGuqkTkaCfMpuXYsRpDyFVDGrZbboc0D7tlJ3dYtWItelFW/ZWSdmPn4oj30pIeqI
U7AHBftaSvIbXodgr6JBB3xP9fcgOTL8rx61OvJO2GOil5YZnxuiYCAU+cAzDYXJtceTQQlv3WQx
EhyO6KbAILQaO0yXORvk7CT/YwthUpt6qxcyt6Dye7wzMgBJcbmZznTLf9MxQoKGGaA9V9JnptKk
GqA924dU57uoMLy4PUhF7KfwLsaxmqLqzQQ0eqipYgQQwxLpLvTibkyJ7LvowDNnZ4+EDV6AW79w
PB2uq6/YlsolXZsb+6q08ieWhtWhJK1wStA+UGz9Ou8n64s03F2QUBQTT0AgsKWtRdT6pWfkruRv
GbzUtumJN+43MNsSbajUD4y5v5LmX7ajOipfj/tKnO5nybeLbJYDWowKoG0sSowgNisEjFtwlx8X
UOscAYYSIXRKGG/j5N3h8W7u6K2C1OQlNz/1EAQVQ1OYT+HOYEtZi4eGPvmeDBsg8CKEdWGRJ8e1
irvvfXLWJCbp4C/5HzSLl5MC2Tn/uLZ2tfTUUktBfSO/hHl5LsnZxCEKvAv0FoFNHG2B6LHXSiCa
nmIjAD4rDwZjLSpUPkCejZDnN1HsUOQYG0FY/3nu1vKDhK1+rT18tqum1X3GdhXasyK9dzndPKtJ
2o6mJf6IpPy3AmLQVYmLU/y8omxf/mNoQ3QdeDOZFVIf3YPbh2qLmOIj/nQFNYRvJqQNMHmXxgjF
Q2WT2CXUJzPYmMPoYYKj0uyD3zTKOrTCEdHqwBwNmAxxMLf/sdgpDNl0e/BrzW/DXZy9G9d8VTi3
d1ov3YL5yeEH0DScMUsCIvtnsP8DguYyehko1pjAhITVoQV6BrCMQTtkYI5jGIMHVM+JTiQdf2+P
YkoATUrcgBICyE6VdR+8plkO6itOYoRyCyzr4AchLiA9KEDvEyzlaqlcQ3rJb2Vgf4NFldQqpqkt
IyW2sWlcS/IEWpt9i8Deeb7GunaIpMIi2m0AY9qR+9AB2BQ0f7AbVdEDFWweC1HYV6kCCp9VQ5Sh
KUwPzA8ZlCD+SRGB9hH1sDYWa4m/mfGN/s1zlpTpYgrDVo7x7vPCRtFuw7wbTrfF2fsUMzYaMszq
b7TfuF6OollAHjdXJ1GBlO6YV/CLi6/JVlW0v35z+erlAK1VxTEJWenB9LThQKFlgmtC1L21/tun
higP8zLOcP6U9TDb4WRZh62gycQwzk9AT3DBeLqp4PQt9XDpllkpFh5mx9/FPGnRqT7QGhucDuL4
V6HZiddSnw3QdoP8mOxzp845IP7kSezatceBd47iHT524p+oqxYVXpubootu/d4n2wFYfEwSO1LJ
LQeQs61RS+tLW7VT47e6iqsAzLb/DFFjgVxRgxOyrzWhIE0UixFhEWkL8zAT9BzUE7lvPcOW7xq+
QbLHM9KE8X9uf+RduWAGB+gxqw1R5rWG5SnGI1MF1X7nvp+NvtXmnhtboyOXjNjcwdHILfYKanCu
318SFwz6OUcrYdevN5OKMSFCM3/2LvNaMCk3i/24MZNjJnGrikM3w8OhzPt+PgopLku5/gHtCr5q
mAauTMSBr1Ttk5QxayWiUJxaWC5Mr8AqrE6FrdhAeeecPdJaZbXeGaERM0AH1/hLnfHNSQdrSxY6
Q5e5tx+76r0sntpzgwpdMwglQG4VVBk8bNqxNlrhrpwcEj7NHHXelIogtFPVCu0MsWc+E2kGtmaz
SJ1+kMLohoVjZizo9SmPa+aiI+pS9TjJ8WzPKFJTvSQSq1p7yWMQwegIEQ1mQm3ipROAklU4yk1t
Fc3fMyO5SHaApFG+HVFImIuTVtbGi5S0G/WMNx+YmKoYDEXW8hMinFXBYUy5pGlNNh6oOKcji70F
1wIIbvv7yE5IcIcqrVnIUMy6jJXOUabQ9qElSv4MA5UrWAljDhZNAfcYJEv8ztID8Jz0ZtWXcPUo
CND9inSAlT7/jRvotW80a25sb6qXd/vqRUGMWfDUYUoyDbbte+78beReHxkdtecq+4RkNaBC5tNt
OdNN9Zi5gjM1W7oSA8gBI3wqGJrb4otG3bhI/y5jO53lCdzKQt57Mx0gbap5XbQGXwM4xbhdB92E
a8Lizo5YrnNFEHsU26Bh2BMtCesTHYIg3qO/l1a6pwQQqFWF0x0zbcRE3CAQ852rOZJTBN77aAZB
38yw5V6LAOjSlkY7MHH5fXjpjhUahKYFbN7MhV9YkerGJwUSUBYX4ghPKF82sW+2Lar/q0u/9hFG
k4Ha040m7RLmeyGanFryRLvOC6doJjfq2GoG5cFUzBQOh4iS4WnOJrDlBIflY/NqgYDjWravEvCm
vByfOT7A4mvkkH4BHKkhS8RJ8W92ttLK4e1LiUv4zZq5N8f38HOgp+b36W+9W9TSItvi6WzxgiZm
hRvnxhTdx7nFFDFV5wl9yKp8gMrEyFjP4xOpSNDK2F3s09bqWIyYx3oPVULx2Gizgx9PI2omjh/U
YGo0tbNnbxa1ed5WJi8YOILdJJdNLqRlEwili899+oMBBR5SBr/B2IP0D4VTzZ9zG9v23Ap03Piy
TyO1d7jcNqDZyNUPR6IeM04r2VQi6I4YTEeLPMYk2xWbJB8Ge0VpEhursYPH5DqAS+c4eTMvQZ/S
BMMjXxv/4sdovg+XtVWNzB9IxLUPDEtUaYXf//TcL5+DDJVRf2aY9b8FNcMwbn08ZKnSrSXF1+c0
BOhOCT6gYOkKJYzYYpKR0PR43Ha6SZCJNEA+7/CIKrUp8aR0XV3L+I54QWShzAZUUwOCzkxaIvnY
/oMsAQq4mXUVzBn/OVR1DCbTQgBrjm3//3wG4E555qr2Xbb5N4EFlnvCQy4URVbgWE1/133BVXAI
fecTMOjQsD4NC5G4IESigxP2whVh00hXPuO0YdOpeBU2wzWYN2XMAs9G25yI1pHtlUfxO+LhXBRM
c7y5r7cExf+AsceOjxWVolT/3jetCrZH0c5J5RhGJyBXQpjxetxKld5gcnH0DsHfNNdOb16Nn1nP
ci/B1vh3cMm3yNqYIQWtk2luyqGCuNQzFradJ5aYfvszh3e+B/rswq3l7Jy3YutShfNMkmIp3RLN
MG0sQrxBNNvRdgIxeLYdagbmENbllU4GXDJxUs4ecMPvI9Ou63ojaIb2+NcXs9wLU2b3FSkSwFqo
VGvNyCyWNVKoVM1+sr2a0K3mPJs7a1oQ0zuG3iHvRX4kP8v4tHYtLc4SauNrLsB8GTVdiLqT6SKT
jKN0rqv66Uxsf7b3sABbAndPb5YhJsdctO27ZXUT+wvfHmN70mmeArt6V8FUDgHvyVmLSj6z9mvE
IFhd+lIacstL3N1m+C11bbILWCGnhx/3fWu6lm/VCpSrvTELHKzH/bKyiRPnZq24aSxlbNkwqQC1
umtzZqhu0JiE051uZzXaBImy3FTi+kjulI6im3lzy3XfbYCdcUBXEtmIHPVW4QUfL/DQ4ptWy62k
GDle2e8Kx+ezZ0opJIuNk38EgoHnWFDnTyiWxHneUKSwd1/8ISclkd0bEVFzPcv5CNG8gZswb9zs
NVGDt+qHfu/nlxAIj3veffwI1Sb8NY0jqDKAOfcgWC8xuGavI0DVZVDiSgQ5xuPAhgkVtO5e49km
qBL7OyVSya0VLokOB+4tUwL6jgzWrGn69v87teSkEgZXXP/b0jJa4Pclv7fvJOMIfILy7GIr1Q6U
KfpM6tBdh4bz5f4f6hoQNLGX+xtu88Qp3rJ6Jhm0sT4DO0gXSIf+P7nYFAeT/vtuGSBnEGrx+DgA
Gj04wa8BsuHNmwYB3Janj3GETTHyxX6DD1oezgmLzDMbpM4cGgswvH8J6TIizSs+GQtFSKMWM6ee
HZ8DoFKrvszruww5+z7KcVbS5IEuKKM24wps84OAOsIKqmc3eOEoiIDmTqx70QRX77UA20Uzlunt
s3lLZ1J+QXxR6oyLBNWR/EFHTvhxzs/2SU7UdV5PWSjy9ZSmr+42yNzBnAO5Ifm+BPVRp9iFFRaR
/2G427wcORCHOMf5cigIddx3ndwZZAwYsKhSmAc4nt0cy67HbfGrpnY45wAK3ll4j1TEUuzOPz6X
G2dNBQzS6wmgZrZ2wWacMcoY9CLVBP7/Z1LDFNPcInCwCENQ/3FXoZJJM73s0dsy+0X1JSGmm8vA
LeOgGKr43x7BTGCJyDaXq8sFhb+fX1e3QyRErSH8qh+o7GWJPvOTC34NIn+tZ4sq7l2GPd7H4W+9
eqIlshlmC0VyUecN6D0QUrVLArUoi7repVypOeOvYgLjG+jGA8Vy5qOFlw0qBp54xtrflGyUiisj
Nt7ABM2/GdQC9m1ZjK2m8SCrYMBnTfRyinZq+87Uq7QC4ts7ES5X22sLaKK3aW0/kSLJN4XV2FOv
rM/VljxKEWrpX/lLqQaWfoITKXU+7qzfXVS9JQ2Y0uHjizj+2pM8bxgi5IEpd4fxLbTt4tBJUqU6
T1yskrir1tDl/6hCMKOpdaNCfuojiLiyr146I+PvtIFNPH/9SmGW2H2gRqGZV2X7SpyKklJamNLz
GTEosRVDIwek0XzMPeaHypJKN7xXvwbxKnc3LDOxpjZDzsRMLTEclPAEKA4W9kTauLhkTKQybnzX
yI24lenHg80AVNLYLn6O/E0VLf65huOXWfsaeCJE+PXacmqcM9XM42BSbVmDnNXdUPUs4iPKSk+R
c5z+eyVXMs+Yp4nf4twGAeixHBRCeMavHWY7RqZptA0VbQHo/e5AuHLBjtYIecxjX8fsWOabf4SO
OLdXeQKW58MC8ne66+DxLKy4+xzLJWVAj57f2/LOhFm16NWCkrZIEJf3VuvwNit1lSamT3tKUD+L
LmbSViBf1iO7UuPOwYPbvpDsTuRwTJkrXLW+Tu7cBb8jzP7pDESS/dJLLJPVsjRZ2kKq2M1bltwU
CKsBVxxrq7MEUxvdSQpA+DPndDM656YyX6RgiKftf3BcXjzl6+NECe3xK9xgmyEwlcegigRiHYQK
je7Kw8O92Htj9Ofh+nEILVfMrEowSQNInuoiT0CePe2YBAOjkoB6RdIyAlW3mx+CaID2QemaHGmL
rqBmagmh0q45d0wEawJeKdY9+EksX+Unrs+roshKb7ad2SzPln1RWrBuNURtpUa4P9CC+DFxy51K
MnT4W0CmjYfGe8qI8KPfgqTNicU5WYwoKQgayifSK2v2bHO8twngpOosjLtRTQV+nqXWC09ULQI4
ZINfwD2eRBlJdHBgm9PJYVinQ9vlEZbY9xcsNEWH/0PANuMuPoqvJ3r/ObFsLsK8P+sGQKith0eN
fDtFeTuj4DRiPViRf0/ohSHu383qzKjYmiYZB85hAdJPONPwq2DPfEHMDT64O5DWgVAMx3T2pR1C
MbNmrCo+MdikZI/4ymdleOTuEhYbiYUyDUpl+8q/tF2+m2zKdh6zHhQoi8NYG81zchRO9rsOPeGo
/lSaJjAp2ODkw3dYO+K6dBVrogOI6oItedGLKsVQmf+6x6u7nwaJFVahVqe7kd8NJo/1SKuRF8Sg
YGs9NXBMi4TIVYYnyovg41hBDjnVumD4bhui08tdcvRpuHtCH8Ija2KtAemmTIUd/xlemTzBdE1M
BdvQudy5+sIJwIWss5x+zDEbSaKi++eati9h0CC6+Doakle8eIKUvJ9ynRo//xbA4zRhsUxk/rgk
5CCXw3jQLWlKOZfJAEsoTWvfS+0dIvznS96EFrZ+yxkPlYIxa7W5z4n+VyWzFKmySJgdg3vOsJR+
CQSdhmt1hojXOOKzcGr/5JX54Z2Szq2Tk7OWSZ5pTKfLAPf2b+d1vJFpUveDgEPfvgmPQ2b9uSBT
mw4gxR+tBUoSk52+bL3O2nAkvDdTchkwBcZN8NgZR3NWhCdcfqgFUOfAyzQxVcBrCaU9+E0aq6mX
dFWqitVYbWj1wOTX2jAeJd136KU5KjFjPmaZdf0aj0qpp7KWOTJuiEtigEQHb6NWX0ALuMYHvDni
aQ5ZY5LFSwRIy+a8t5fOFUgdxDorQ0Yd7KA5ZrZJwNoaZt9u3n9LZX6+Ls12T0bbzNRmkfmcxcqr
XTM+EfkiHdgo0qvQY2ezbDvcOsxCb9v1u/C5r1K/qglbbbbgRnnysDp1Ev7Mad9c4M8WLlrrSY6t
Oz1tJdvUnZ4TbUXnt3Vn0WsiCJWClDMzBLIt1mmnxeolWLW4KfkXYzZbCNfVC/Kr2fqihIQ/scWL
P+oadhz64o9O9q5LiYlfSY0ULUYvXbS0ETr11nNGn5jFfrVfPNsXIOZiJ7R1Uw3XmoIyf9jfd09f
68g8SUqgyvHDZSDnuJhRpd+zzrmHbz1/jenT71Vr8yddy8mVtOqnAaB2/wZWbysa6y0BwwCahYSf
rtfA303aHJTPC236FqCXRxRpD6uebBD8VwP2uAVjSyBUqjr39+oBPGz9n8xLXPi9H4K0vXDH1w0H
I8PYekcy4GevjUfTglT6htp02piapkyIFe4dgMR80ci8xNsd48RWQcMyikpgBNrkobsRU51D//N+
+ECEHyCOlQR6O6tJKCreNSN3UUeZubkqTXqAll8y8EWfqpLxCdoRmMnVoHak8yHwoWkKx4VD0xAC
IFt5GrEOXzvOJ79g74mUU9rWfctMzOzqj5SSte/a4CRC1ZJ13HbFLTmAEWhD90L3bDXgOxg+TX5W
ar/jp5RmQmKsn0t+0C6brT+X7h4fgPzNAlFzAlawYmQKdn6oJqDejf+/jXkM9AAM7mVMNuU/o+NZ
PM6D85YxK37Ks4T3hyIkA1Gs28/wTKN+LBCviCIgO76otF+gaTlqlDymblTguR9ino7FBjohjoTQ
xkw2Y2NAj/GtSHmF+0d7Vfv7AuPtG/ldx0zCIyMi2+W7D6cUi6ZMa+cg1jIKxOjz39LnmFxkqfOv
GmRYGvd3EVYPEJGb+bLtzwJYnSprZFX4yF3ktfNwL7xpmlmN8RlBNMLFd9f48fbft+Fn0+VM4ixs
cYY4IPdLTf8dbe1BYhrIMm3Bs630KQLBAWXv0d9qTtrSXGqco/NsSfxFIol6XHjQn56EB3d7o/E6
q0VLePy35sL/ucB/2QD8YSNE0museiVX/RIk8i8gH0MvhErltVC/0CoImS7mSh/VXhBbhQhuW058
yAD0Xb90GOEGKk3Rxw2jSZJDuDVS10zVxNnibjYohzqzTqVAd1GGwqSUlPHScQodKxRdiptEfTLc
efdaqplVJQBeTQoG+a4Ot25sA2MAsELijpIiwXrh/ELiUkIDc7X3ysrrqAo2QjlzravqlG9rwNnZ
tGZBjTGTUm/qPdHU12vabLpSK4yhbxEP1+AZ1Cp6nrdoOBYPByiknhXy/1j7u4/HX51zfHzJg1Bd
FG5oOIXULY/o1XvhTkRUSERy3+pnpbeXQ7MsB2H5BnNG3m7qhEKABvRDtBFQBbd4alo10t08Ld4W
yyKR7Hn4DAQF7KK+PTZ5yvX8urUPDwwg8ukuq87YnhPWNa8X6ERJAyz/ZVKP2CjXuNzLneu1RznL
gk3aVFMxGVvgOGjzFovf9mPCtIJyzNOqyLZ9K4OwGKIN8xiAKKmgv7R6dah/hgfC9CwUPLg8kOPr
a9f8LQ6sBgkhe50gAThaDSlOUP3dOGmYRJIc4mw3HwUl3oi9GDIr4sCm2Vy2bEiXp3o3SeEQ6i5q
HwGjYuPm34HMp6UKIXWp8h6B2gaAgU+9gRYUn0WD1kEz2URiWvMuv6/JUtJta8HxO82f7qSKrlMT
HOuXH/l7kvTExVa3TnFQqYZFjMMTeU0FFgEbcVIk6FMfvIaIKFLKorlBAFByLv3amfd9gQZbewAo
wwiQTOVn44AUiW8TQcePaX1HfkvMPMKEyCphx5fb+aWMVTjYk4Whr17jCGq4ids6DA6XSa8KJMO9
o0jiSWYXgiTs6YkeJUZ9vxO6LzUBMFdkOGWlOIeMb5SNjfLamCCb951jHeI+YW1Xj1nCazl1iWbD
BZ4CqDbLQ7j8iHELWjIKQOpt9ocX2drFzxG0PFvEN/UuBqBUF/hZf/wMt1hU86TNMrzzjaIGBHce
esZZYrtLuQHnJswzTUpzPED6gSmyq4Y9zxVtAhMVTZDsVu7EuF62iwl+h1SCw2m7U0FuSPg2aamd
dNiq1W6NvL555kr21Igzw556c+mH0Cw9ii8VIbo6S4tpSMmezl/l3kVaHFxxEaspjXwlDc8MSca1
KXusK4/kdU4ZNSryKdfKSuZPdo5vNPwV1jkV35MH6SBKLAcZBXxchTqWs9a0zOlCYFyuhRYQ14m3
au2qqIp8sMZW1wp71YEPLBylhghajhkyfyg2wWwypW268uHTcL9Qkn7jKZT93xgR3MRKAChpuhgQ
JS6XaR28bd7Tyats64fOTc2yNIJsT3xEGlm53QE67fIQGJxtNy/mls0DAA0xVprvE6IRW0Ti47ZX
wr7ItyvDs4kh36QX03kNksZr+3MoUajgvn23Jp5/MMnA76Z86UIFPpE0xupLOhpSeVVLBLudOiOl
J3RaVWW9wm6GF4eXWnoYJPBrA0IMUi4E5g33NzHoAFPHrw5XQTNyGxAn6/EgymY3RlcPVyGv07Kz
s0YDirdB7tBblsCfMvDS0umDt3KyZ+JLxavWCZN12FEXxgxV4rDEbyM32U6zjYbwRbSmPweWsciH
BmaaJgkAMip9RFZJmqPoR0aW0lskTnv11aL11nTTs8j/R6N/dDXEu3dtqJ5Ir8Qzs+k227O1Yw4V
q4Zd3gnQkNGQ4xXfp8FZKXYrL2d/SiFNNcDSM6SxTrw48BbjaejfzOCqj1mtjRflnPjDr6LMKNYg
wOJGoRAj/u6lRxU8+2RK+4nIo66czPIJjYZIH5UkM5goU+c8AW/GPVSFe8pPKSnBOxBTIEXAdC06
fbZNhpxu7HZfZMc4dzySbb7qQfJOn+agV283SfvP6hMEXf+zhQmsXduWAKvSllpFZaKCc/ivSp30
+IOIOrrVv1IcJie5sE2cH74LXsthA+mJbXupikJQegMf4hC4vyIrjUUxbz1N1Pxus78NiBR8PIsI
JZdQ8FQBUr5nub4xqmo4CVkvoaC+ZEtGjS0ODWfRd29fEoIswMddA/5yAKwJOc4KgNv2JYVzLSYt
/wimslEMr6g1JuJ1N68x6mtGPLEPNiRzSuAQvVcS0lp1YiQTh29l38V9fdZajv/ppYaGVAMahO4n
A3GUUe9Xz4zQ0Y8VRiRYe837bkVZkJVU2eoZSk9qgVmBeWiqBRhlIu9iqqpbcdAu2Q1FeH+JS4LL
ObWs9bVNGHlVKATOwOyxamWGVPrzL+swH1pO4JTEA9UGwtq2/VKHAGQH1UmKk25dP63r4wvlD6TP
J6/DjYna6cPc4hm3K+Ll0NhWRdmnRXGRQdUKrh7Wt4qTfAhe3jE1fHl7wDonDFJc0xGxxpJXniYG
OSZvjuMKGBWB7ylu0dDEHDxeUW3tvktdvO5vL++kz6YeSwL9Ggvdhe3BM5UItYOIJG2t41TZoA0M
qv2xQmHcohR95RyVlWxMi7j7GDFrAebGLZbDsAugovLVSxk9H3C2EsBgyvB80N5Zxehw7GkYo4Bo
6AFQO88Gvpw1s0uTe8AFXIUuzqHbC2Lz263mUQb2dRg5d9Nyp5/7Z5XfKRaasAFE6WLedtJHf0Zt
1ohwr4XHF37Z1FvyWpVAs+a9LR2J3mvXSZhEOUO+XLue6s9RkJcSQS2rSjtTU/k9aNHelBBJyiBs
Kromrh8UfC0/w+3ApcTxwUTr9wAsDZ0kIijb55OVaYhetv2X5B7lAMYMFvxBtlOUBNx+UDeBx4+v
PXHi9qo4T8yTP4/14JTz/akTzeoxEdDqJ2XAaV7eOkpZ4fb7aZsvcgkA93sRmJllrqnVgSTFUWnG
kUF6xS/f2X4zD0PrT2nH4A+4NSJxem4qcCqK29KARiAmhVSTqki19XAo58kxhN1X7dCb/Zc6legL
LCarGywz8ksC7yd+vL0wOFGUUXusiAn1vhRo4OnnkbKtWjnt7E+KQKnG4MWU4QN6ZsDMyIUoaPvU
IKMtt9unblOC5DsjvYc8wxrBzKylt47nlCSLlFgnu17TjR37iLKpJ4PaBPRgE3ZdfETJ/xrXSgmc
oruw4GqFPLL0V9sRKtWeybHW3IBsU0csuOjAebhS4SCsyRgrhdo+6FzmaVEujS8H1yHWuknIkPqv
Y3R99A5XcgE2XqKWfEJqcONwRrtuU7iptJm++vakqA+FebTyLa81aMBFNh81fKF0rWDZqLHDDRvz
nNojKst/IOKqXtEzyZx0RbYchEqvZbPuBGOn96itUuXEbKO83Sk4Lf/CtzHVy2kSAePi1fOWL0S6
MtO6zPUNLR0Pd5IAdi6LgTuFxsJbFhOtcOwwRkV46agQiOcfTCCCFTCem5Gi5sLtGP+0A3ePpjLy
HvRjiSYhuqqHE7PbG/U8m8RWxfI1Pwa5Va+p4C/6ZazUEKv5PLyZhd1iZXVBhbwvCJHSPlf33zi1
bX9hAMQtaTS2hHRxEjdodsxzsEEGPOPlt316rFmpswQxmfMlI3oYqSWC/O0vNY44SEj2x5KdknKu
O9N4zm8HzIDXxfHUOpJdyzrACeMTob1dI46Zxl1YatKd5/rVGSPGioOf4/LhMzxyG9brQdla1ri8
dZosA0YuncSPM2QhY0BD2ci2PXru3oXn8J9nb9p9aYi3SOLs70+qvepjmJGqAuF3A9BSxWo/vshg
xiYilEH+EJgC8chyLooHJm712xf+8bWDGjmVSF0UGNGw1EG1ZZUCNiIZ5FXMu3uhdxxt+5KEqTDP
5FYHJRENvCZTTl03fMQefr2crzJ8XuaEEHCmIzsVYwGLVOrLp6ppMy05DTO72H+/1d0lDF/ag1wS
08UqswDKH8Cf8XvEvzaOgvupkNnninC2EmXnKKdKck/73vWp95UXVBJtvKPUdnzEJVNSi4ow1gl2
deztrBCFpPB+gL+QfYgpFQSgcmHMLsQsctU9HB6hKvl22xQHcfEnJa73OstHjnrTrsXSTBuwVGM+
lWsTObTER9mLMZiN8Krep0Hv+Uwok7+CdBWhFdaYWvN3khsyH1ZPqpi1UwWjb41S5kTWMuzEY02Q
erxWn6MFWhriVVaYuLcxJF70igD0qq8HIX+lUpTNCial1KewMj+V1XNitH5VHcxyRrrdohErMYxe
5cFRzb2xKxJbi/JUhGqj8TmgE3bQTxZl9Dnfv+UFw3eeYevPpeUhliYQ8lDYBdC+sEMmWIGuYhTy
yVJiLXGwy+wJxM6LwwQd2ync5jSuV6vUTXQE4aZpHiWNxXVEz4zybIwjolCvtI4G7zDp7XCI2Q6V
HfgnPZlM6f+a47cij975OJQVmMT1uvyf3Dllke4S7RrxCaLH75KLeHium7QFHpE9ilGlJOhVYlEI
jyI5tVRkEacm95OzOfMXo4B99nrJ/PDmP0+kmu1F+D7V1z21/vfxsShuwHkJIyvuSrvP7BZb8Ma9
dqqT1YHPo0gwGReDv5Brp7bMl6jR7ChuQpDTE8z34CuyH9vvYuBQu+NxQgR7rHguxYolgDWwPUhX
5aXccD1soZ0QtOSGQfESQFIdit/qbkj2cMoDHHtO3NbyMcecKRsprgLYU2lFBPqZKNney212pDbS
xfqw9Go0cIUscSKpSMbBbGH31oLC7rPMdAGi/U+pecgOan3vbEzq+x6vVjzGXd+BIaB99TPEaciU
7kvJacDZn+gO3kTcnRb3GGtFp+wlWzN0wMYMJYHuSz6xyL5RfjohH6Zvq5UIdu2bh0YDs6VGr5Oq
pGMf2nhfvWhO4pZ+y+366gcx1oX4GgG6wJPP34T8ejrPmQ0mJ27ZCa60IG4+D3w8FDkb9jjFct1Y
CC0hSCLdGtGHFrXwaOAYR2prI2qsO99vRO0yXoai0nxpLJJLqZE74pe10NP3pfaELvKt3kDYDY0M
UQ8BBB804ycmIWgP3qvZqHumxZfitvwYqQS37iD1uuEqxRlyen9M51D3wbYAhHQQFF69YbFW4Miz
gwKze2i/bnBYwMVs9AyPG25tL4v2/5K2+NLYtD2oP4PGLvVIRjvWmTUvaHWM/RGNMvPh8xrmSXkV
9nHzT8zCnckui3C0aNui+soZbbzNrMwoXNbDqPZ5JanZWH+sxpccp8p7RYag+doOqX3lo/zusdrw
Em65pgW8g5ZIrQCgyAV9L8XUeuFlyuONkb5nZMbNfrrY8cKYZ5MQZb3XnxxWi64atVYaC5QJA/zj
UOzQLfi+hs+IAGYm46TWH7Nw61BCYZsCj88wmYoNeNRIEtHlfgbODqVbZuipl908MCJShLCc4+d7
6BSKpoj5JRLmivIgTWXwWGQryR5LuGSWNfunw09SgjV3iEYgFk/SH61kb07NwSpsP5D69L9NWbM0
NvvZHTQdRPkdur32B8r0uG+PF4F8JGzz0fiWRbn1gYsudq9wdua8w7OQwIHeKxfU7keYJWngbd3Q
IbyhZDyAPPKYzicKB6eMSPqq/+W4PffosfZO7xTdjGJfWY1qO/tski43D1/rNJiA+CeX66B/WV3f
cjzfS9mAlZ6wp8dwSNnpT6YvKTuKcX1+MJR28as9X9vF/vePBtTXV+8egpJbJKhBNhTFmAt4sjyl
NZRFBMk+9xOo1bi3LZLvIpYmZf4B/8QTHJwmrd8d2xddCXfgYeTacelY1WMMHs6BtX1ZV0pjcO15
RYfwBLIwnO4JMwfE1Zu03JkFMuQfRwYrGOvReQA7xocy2eXHc5bybgvXFb3BO0Va8RTTFTAzCxkE
hoaPi0/JPOmtUxrZCCjw82WZmRiZBOxDTwN3dwv9Ntkk2MymkgfeTgPNrWVOM8ohEflPCqvvPuPz
wWAzRtdcXqF2K11TKxNCSG2OvyXxHhuSqm1UAZyudxmCjuPKMfM3rt6TYvziKlUcblt9kKc99GmL
+j4g0nsU3QYUSQHXLNxlBW2QzAtcinEKpsk6UclI+IH0o97OgVXE7wj13VhaxhKZR+DeDGGAsGDv
67wMt0nTPCQxtkOusFZuQSNCc80UKg2+OxGFQM128lhmq6vJ2fExS4KDfZ6snCFegQwIsp2/9VXD
V2QB5QwrQAnYFWC2oPUMNb5ZdjU/a96PugxjRtFfSECZcwf5NXB9q4N44MiezN/CyjnBIKvorq3p
mKhGUVb9mAOlfbkUqRYLbxmHFGZ0O7MqDU/FPyglI2J9BQxIZu9U4xGqtr5f7rymKN7JhM47XiUk
aKqLrKCgOyUgf1NAsFanBibS6Tzc4ibU6qJwql+nKrUJjOOY49NKUxlBdGh4z4ErXrmtUaJ3kEV1
h0acB+Kx92ishiJWwv+zfUzHX9gJ0E0tvsvSqyyW4HZwQGTKjvJ/HEtiCy+taizPGsldGTyiuv1K
k5D1di0FM+F8nNfg67QnzH61J28Xn1WWKXjyn+NMjcl0Jr7zdboW9MfsSpT7mcMOUntAhEzq21lL
iCKCK9zeA39YdWL16sY1PMBvePGlaRYfMigOBLfEhjgB9+ua+rA9UxCKwgIHSfZ+F4fuEflBpctK
nYeEczcoOOmBS944+vMsnYvwbMhhgO1i5MOnV5sXEMubuKLgMGdxMimmqRo+vQfxY+9/PHxFZXwk
H8lVdPAH84yYBbLzBaUUCwpde5RUTf5bJQxjPqm0MIZcv100CLsR8qSpADU4eRU+kAHg5x2+wMRs
dF6+a7OKxTG03Vg9S4zATPwtua1MfJeAreEpjcKxigZmv2Yd0rG7/w5YMs1hdN3JEpvnD5HFbDeA
kJhz5fe8hptgUf1x4wQxBz9b5/k70qgcspXMdFL69JXZb2GEqhZakyep14WKZS+QeUUCNnpcN83v
DeCv4/X8/iBK3jOuMycxUyfzftLIdWqXgaQPv3A23UzgQj3BnJps8xlKL1j7DE0rAr6nSf5i8/Xy
6nUwdi7ZJ4+6P6Uzo7RJ/LYCIM0WrXrxASpJLUvAiW/hZ58J9+WM61jnsMeaP50UfimvKrz2ERI8
1HD5V5iMR9W0UTp0Ys+9ROitcl1xGQS6RVv3xVC6Z8ID7Txe7d4PFYfXfrz8WwXSYsQqqxxOsMZJ
eb0vNbXTC/1s18z5oqdphQFqkj1IC0ha/1EsmlKfz0fcudSqn1K4ES6fGy0xiOgKe5LL54HNkmz7
494h8keTNGwjojpb+SeOsFiZvYDUbol5D4R3ZMTmz3wckHb41RU57Ng5x2nLlM0MNOnT2d+F/6dl
i9N8Wea8E15haGhsbZHb4X4miXXJ12Xqt0FR/VKTy6ENMWB3jIl8cMdMZ4sxSgAS6F1FZ2Tt4kQj
YmbTfhdird9tGhM6h1XtwOU3fehObceQUP30R3osrYdMjiVA3yWSJKpC7h8CNxfMKp0exjuXtYg9
4L3dXSwPHbvTo8QDT4nLJigDq4/udRkmNzsMNLRcjz+dLJTagvZc9tDgyZcYm+jGtpjc/ZmL7+j4
oCpXkyND8wazW4v+7pWi1mtCdxTMpQVsNq8cV3NSbFs94vGP5JO8G74UTXozV+er5iImwmPtEx4e
aORz5ixiCaN/cjTQZ4Lg72RB9cDDUb76TJa3P5S9UVSw3pDA57st2Jxn1kQPCE+rKWAitLEH6YR9
yt9hYjvxf6fg9sLtbEUSg1L4gTEtCnPyGJ58SU+JyCsA1hpjBfyAiSHstvqU5QPXnrvbubH37hDl
DfYQxv3EIS1nrk3/Rz63RMWPJN2PjKAvzkIF+ElDQpnMxiEsv4Xkt33vZy5aqIx3A49FTpinhY5H
g9iI2Rt5fcRJKnq6Egtt9gGRxQ5I/8Lpy5UMEYyvCX/sZlqaLD8YZNF9aIIKbWpUZUasSLlTVWIh
+zfhOJplNrROX1ltin9W3Jolk8Y2tH3Q+K8XC6tyLtWNpOj3tD4NWsSeCqwk9gQcPfPIqp3/FQlL
MRaDDz8YtCtm2wYUiMMY4uWNxAUJZ1aP6oFW3yabiwd6KiaeGPtZl5M95PfBI3t+y9zy5h3xrCPt
4rwWtN6hrXpG9uvLGkKbsXuZkHI5kIdGAGarHIcNrTRJV4eh9mIh99OLX4O2H0mpyCyh5Th3pbhJ
DE1JOtS1iwKq6lxRbpiCpyp5dOBL4fgzJ9LBanOu4iNfSM0L2Vqj9nELTOLhrcoEndVUApqRW55m
6GQxTD2AhlPxflh66nSIqtJMao8BSNBSho3RbMbwwJRBHh+UwyN7yQB1XPfhIDe7FcDY5Rhu2xYV
ccOZU9KAs17dd3R3PNy8WBAbbVkgbLY8BrQDcUw9fC/6HLTGec4JCCdSiUx5ywNh7aL8RFztV7sg
fX5iOzaqovRRpMFHTPxVK6SgwqqCj8VAsbrCmcoMlTVDDkFfaZmKWgRghoCJiuKHUq1K8fOiXoW4
4qM+hAcH90g4CMrMjftCOjbYB2Kw19lfaJra6KN5E/AoeQpJ8KhWOtHt0pBewbe1irvhiLlLkQdR
hnQ0mu0OdDgR0dBA0+/vfNkPc4PzDj3QsXwzBXey9Dr+p5rq02zdURefFOgettuptgIMgRFMala+
EvW8O1BxF8IDpx+/86P93BuK0Z2+GAKlRyxo61WTU8CDWsEKYjKSU+NXiZsVfpElhHL0cjjxC9Uo
sgbmhDh7RtDbf9cZ5AzSVLVGBsojF2O65KVEWQwpqyEYPC9n7OlIFbGl0/qwp7S9xihQeExoqkPy
lTxXBR+K+GRYdkic1xjqt/hhwxo7v/cFLx4igNlIuriQqnHoiY6E2chXxHuAYDXFoHTihcH6Mt68
d0wzXNEezFF+pBeaEk7fQcC5KAR7KzYK+fMSGyo9/wrDBQaPA2sJig70JSmsnQ4V8dlZVimDs9wM
K3ZW6ygskSTHLMeZj8w/p/XroJwLn2BHM8RV0FBakWmo1WZl+I79fuVKpbdLW+7Bl5sHWq5pMBnG
MtQTK0VaEWpJ5jEsH3t3p4oqqBsEeWbOF6Q9FXMkQdOV4ATg0ZSqq7Yw5zli8b4OHpi2x1uK9CDh
dDAGzAkfnhCx5K8LQsPYdu7ZROXEOY3MIA/LUa9Int6ld/mMXR10o5p6mO6viCYWybXXEd881kzp
JRIlqBDNa0UbMwHdI6wVm/2T3WFak9JOlpMmu6AuKM1+CI5R9rjx7NRpXTQl97uBbcGkkrAWFLOm
OgBf63hXa/9QnVGAxIoK0uYu3Ltl7yBWS1JGnGZ9g95++TtltkVyLcisCbssM/UXOyKqHKjUu8GA
D3zUTUfRrLnHvZMtTfBLjyq3ksy0q3V0m4R8Ls15wYuxhF8cB7fzokF62WWItofGcC7uK+6pY0Ms
D/QdMtYua/8b6eJJDAC5iaVKu2/4AJM2zpCI2UspPVXYjswoknE5+2ewyy97HwB/MQIreA8ymPaE
1T02rVk5QCKuxHAmPbCthW8LMwdSJjqIBKL5l49Cz1YQ7bVyuMAdjmoKYwexMRaXbSVen7cTQReS
nSAlAJj2h/c3vK2uOh5eXCXSU2aQZ8I0xZEJhWkke6x7HF8klNTDvz2XIBQEu3mGkdqgDzHTBO9h
cT4Hw4ad1V9eJPpgWWamcHuZUhYhCGMqOKRn3183UM+BT1IIgUq+ud9nPBbdgx6fyrqcP+bknwtk
QsNk4dQGJK5Wsf+oksXtmgDL+eaq8fLzmlaCoSDAp9wRHHVAqYH9XBViu9kV7JNYfQFNRpQfZoMo
MYYoObuhF2RfL752BcwrY23O7M4UwK6eRPMVe+3wRnabq4/H/eb/FUfeoN5yCcEfMpZve2d3p4oc
cgp+J5+1myZOF6uwhDLyuwP0NQogQflD70Im+nbpwduYZgOGaZbl3YZvi1wLvtgC99qMfFVwC/yj
nFgDVL8B55Flakei2jvIPdab5FO9uU17QSGgRstZUTRic3uNjd/+WJVGmA85N5+NDh+554VzRtHo
8AfLbR4NmoMCYjWqJRPOH6LyM9P8OpamjDg7dARM3h0YrCzGr81q4gn8PR4q4WvmSloKoBeEC31a
Y7dp7ZQsxxaOu/ny4pVYWD+7N2WlDb6mVdkk0s3ApXWVroddkNH2b3SPrP7jbgIK9+TLtjKJ6y++
GY2tElUwhW+dPWQcknFY3GVmMhS/xEcw231FmO8agFYGPF9p52rzCKfSmvChnLlWQFngNmdGWcy4
Um/Uur2ImD+wu9qKREbw4zzgrDg0si1r5yNHNwuElDud/5WFX8odc1H5+X/QcmO/wP0L0ybLErkp
vQUO1wtlqivTYj7qb3oX8xaerzLwkMhX/quGL+lcFCa2bFn+94yhTR0xZofI8TcLqo/wtjBwf3Kb
cJ4ovRxQRi5d5+vTbDl7TQFq5jPdumyQ2Lzt7r4QMlVPzm7bH0mzVTu3rfhqupcOQREvTJ3QNJv9
kpCcsNmYnTDSlqPR2NGhupVaX7Vxg4u8UaVJ0/fugGfWumTrjYoTroenpz2Pgd0ZcLXNn3Q9UPIt
AnyaVqkxLkiI7YmMIBa1HSJOmKraCL8Q3GfMTc3lt1Y1NMjnLPxnC7IzEGWxPo6a89NW+DyMbyKp
CFL7XE+S+wenlVug+ymMZpNtCg3KN2iP6MvCOlDmdzb88t35h72yL49Uma/NUePdRAzhHCcy7n3C
DIy36AnvuMO2k8d/iApM5a9xmWnXAKBy7aZFuEYdR+8oTcvp8lcmyxj4Qkp7Esw5g13IqgDtmuJN
nLFj3fIIQOfIn+YfhTU3/s8TVlKlsMfhNGvBSh4OCpcPCwGsWfAQASMCC6G8jFhkzsaOl9Pp6MYG
K/RX1HYcpks5Fe1yOLHklHrc5nepAdImUwt7apvMA4fwWDQVACT8rXbPLJu1O1yDjoW+ufeNkdWn
47QwOr5LeJ16UTYBz4n90DXRnDpLzW65tY31zIDZnFWSz1F9qtdyGzMrvoRyvsmwyH2Uj1apoRUl
o4ja3xZ0nZrpazvpJ4FfTJT+kd4eYjaX4tBcnXfIj9Y7cWjSVEwleh+4vPxkhnWdjD5jlGWxLpk1
5wAKfE1IAcuMiyEk0IC3CX143IQneUk90L/3XCoSzXt9YuUhhuZqRE4UQjS299uu+MN3SxBI/Yst
xacAsSveNhMy+TjBonEifqAnNoF+GjnK05nPGrdGPGf0ApK4mrfkym0J9UnWPBM6RwY8y2E4GiDl
fNUkgZ3tlSLSk8T3Az5+coaKzrRf+SlUeTk25syjrfgHyw0aLrsFD6pSYeRvWZXY4XOlRm0dtGPh
jHr6MWW8sMiBYWSBP+437gnhNVbrwJo5IT2EVndS0CGKL549Cz29SCzQZQBFzt6vAI/+2beaXVak
jSCxyyZ+s+mp1Vx8THxn493WaPl1SVWMy7jkGe0SoCscv5LMJg/1IL/A3+YqBkLsfatAruLJYqJQ
T+V5JDxE0JGIgAv5Md7iVGEdheZKPhicSsMmBry69xqkSKmy61nCXZmPp1n2GG0hJZeOOpbx5VV9
BHD2yoHaac5JhgFfktQqTzTsfOJ6TqxEjQr9MrAzI/ZBfMEly4/iG1YufcXgGMBQEA3nZymg64rp
BFyQW7gfXmORPdUw3AqJlUkWUu/R0KB5SMjb6Z3N6lFKkEjyDLmW9Aw/mKvSBpBN0nVOBYIDhqJM
LSw7uX/ozrHRa7IGnoRZqIJA99dLNDS84Cz1LUQyoBAjUHfLbnfm2IsZgpSTIVFkpbvnPoXy3jIM
NsQ97ehcEV/eIYmz74/ZE+wrOeJHKMcCdbqb24CRsERhp448USZ9idlPAkTjtdXucOXpKauhebFf
Dsz4+I/WIj2OCAigCcab+UofFQzzYCEC987KaBZRmSlfeF91e0tFV4z+dIkqzZPNTPDw6rab6KGB
vHWZcWDUrn+5FVUomw41m4mEcCNmLyk8qvxhLjlIBZdQTN9eOLVTxjJthjONIboJihVqOO2yK2be
KM4fPYZJhbxha+ZpYSCkFt7tYqKDoyBMF7rT9Mk0SQANDv0ICSICbkQSRGQvlSRdzSg0GkokGw/1
n+VOar6RFoPthNPICkZEHIgjrxvkGBhXEvvmQZsJd3wKmsjw2jEyR6WtIzEUv1X0uSig9hKu3X5n
7Tn82Iyj6sseWEMSASu/6TwSEYNxMo91ycw9lBgnRr8wJCHHvDpZtDJGnUt8iwPmv0DFAEkEU1Ra
A8QFFZ2hxU+jFCtkhqogD4RacxGHVaqQRlwKpAd4acDFshEEwafakMlp7sP3r27Z+8mC7S174Tjl
H4SfqJC+qyd+ZHEQb2uqLYbh09TjFx2JSTQ8cnRaMb+VJfH/SlYyyZrQu5eD6IoDzIpoUwu/BZfH
GuIDXHKHfI+t7+20C110wVAr4Vb8v353uwF9urKlVCCF7ixWcsNmwWuIFmUMgHV1wEoPWgXilt5R
abBBdivhafydGy8+uGWlg4/9SmS0mZ5C7GgW2ytFK+bWQAl3bIGqcDEm9y9kopso6uiCZH905+eB
Ef6zaVcSFV7Kl2u6cwxZ4PZtH1jhD4LHinTakx/xqgOey8JiOfMXEvZdMls27BXpb6AepFKnmn+W
FHfrSZA3quKv38C9CSfuuqBTzcNvgH/+7gfDcm2N5UoJT361lXjb2A8tylYW8VPvFj2AkQRIK0h+
rPOT69ao2aYnwmXmdVEQow0PBb8VQGTG9kV63IVpB80U/VpBvkt/dBWmHi3rEio610F6lj7DGyqh
X6+ia4INr0t0bH7VPeIuv9/fKaF2KRXp8ACVO85NeVxGX3B3uPHvFCCoNAWp8RFh8Kx/cHnADplE
sZ20FA/cn0TyxZ7YLrZdYofqRbNKc4EM4dFtX0iii35pDk2rHG79Pxzj4VJ5NDvBQs8CJ5AbiEep
MoXg77G499p4oPOGZ2eMdob56gIPLW0KBunda8qMvFerPLE3DdZVQTkmXasc8LWkSar1j4YsuO+4
reAShbtmNa6P7mTPbK2Rlle+RN0YfMoiBc2zpZwD6Tm8wyVn1QhVx4gGvWd1wiQYXecW+FTVbw+g
Gg/wnoZqlXtX+KD5EJ4X6PtSIqmf9SIz+KGcpHyUzqUKVCTrTKs9j0JzMasi6d+7f6wT8bhDgGi3
r/Sy1MBh1Zrio74bjB+VUF0Q1XzKEi5HnzBxea6ylp6oxFM093r3Qm124IOM2SZJP4AbnelMpiFa
s5UlNRT+h7LgcgFSXzxmxLc6MFYM/LT9TulisrbRi8k3wQiQOH+oRtTqtZ3mZIbZZPYiW60+y2xa
1tMKuXq1RcVNRZ9hIXGa33ZoZwL/2BAU7ek85H5xzD3vtdnB9YyMlNzWGCohvywc08qIfm4ypH00
nRELGcxVXU80qHV7Qv/RJT2oeSAUYd1bZXfHa6Qs/XUohL6OJI/eyEKr64663VAFitm0nnfNe/gz
8Bftq6PZAdDKT/czfbg11k+K8gdd/pt0RKSqeFKhakn+OPshsNDQZpubUgZLTm5qGRGbQ+uFdS3g
Gmz9QJbV7+5Cen8J3X7aN8K5yB6vn93xMBdof2XQCuyOFQG+0RoT+pxa1eUVKjOienBwoAv0h4v/
hzN47vTxlJrgOpU6QKRfUy+NA3V7vSLAbC/awrPgnIIV83aa3nxGaJn4O8LmIwRivWtQcAw2Vq//
nvLrlhvhX5bNe1gUbPy+YTB1ZYSql+xFNoTOinWsxhm4CK4B/3TSgfg5qw/k8dA+jpOQ4nFLWqjF
J5Hg9pa8uHwdtVRhVuKJtzh0CkXgJ2xAcfzzefJ9Cg6dGp15U8Jpj0scoPmdK3Olyd5fSbcSOoLP
fvFl4QLF5701sn+0n6VXyQSzDL/h6FqgNDMS/3o78HeoaR22zf3Tf+DtZAVsQHbjUgQODNBUrlNZ
V0hesq4OhlWdOpWOXcTO8zA8ajFpLto/L22d4vgG1Fgvbkkob6EzoZmQy0e5eCLs9dnpLV8FPYGz
xx0W+o8hv72EMjlUzjlJ1RRnluyD/gqye8DUqV63b672rKyWVeUQEJI5ZwJncMRoSEleTe07J7x+
BnhLbAGvUcnNOwWruzGyZjRDgmP3uLulnZgo1VCTd5n2kp3ZJI/rKkNQ+HAq4BDKZao3En2cTQB0
DqYDruoGx7dF8yOqN+H/bjLGJLXrSpFpC4zZMc0cBSBfeFs+86J//2vR8/PO0HJnVGRqoyqNobAr
kZ20X/Xn4JgyN5lJ1i/86owBt4ksMRCbSwv/8SRrnIYZKl4TvQr/pgZu6o7sw3mupwH4vefM/klp
mrCbUW/RDqA3nASljEKAlCl0KThqRlkFO+qgCeqooOyjDH6S7FlZZ3R3q7biDR3D4sQgx+TntbAh
5fQKYbz7On0t+wcEW4zd6NzYVmv2sCpdhi3O+qX0/41yXTwcvRHwIf0N9RHHiKCbZl1UHYSJ2Kjs
kcgjcLom2pcwf7sGrXZlC/aXo/sBYQ1d8a1LKNZjz1wyO0FCtWBcLN4+JVPudFFhyDEF/iaSpIYC
sprpFg/XGiAPa6QRlA8jqORrscIUqVBDcULGWyv+ykNXqRp0SCdQCuFAu+PcgD1llkM3gSyn4WoH
U1bFYqY6nuU9qkkAKQBSQyWTRNP6ovyA+ZsR9ipGWn5HJX9UgH6PfreMJQekHDgdYzpsdPlGKHVM
t4vPUDQZ+9EgXFtLqjBLnnX5GzVq0ty+sASWhw1lAA8Vc9bot6clks8oMcQifzW4LetroNdpHarn
78dwoyPb6nN96TUT754Wv7tsp0U8xlbXf09RoVlNyvdL5rGaMN0dCDLn6t8wBkjVoDOx8OzLqldt
FjP63sNj7i6VUvuY8eH2byHmo40//CcK89drOVwY5VV1Lc1tGMbxCuLf41O+ipZiGNsaSHFO0Lf1
1ncjX2+sKvljdv2tFVjitiT1UzadcUkWeKibyIW+CX0sm1+8CKfVD1xMk2eI2FtfrnRyJDY5mnon
PUPm+SRUuUEuAmJ6aMxQNjy4iZ7cwY2LY45EakpHmLY5p+lFNpm1eU+/ZyTeLsfIuYuo/SIGq3QW
bGMBmdj75wcq+80SgxXKFI0ujZHDLIjnScq1JFyjM7KQSuD0b3G1pv/pQ8Vp97m3D4Fh2YM3q67n
YuU5fkhTrFFOtMWNldAaRJtmW8BeohSSSnCPRmJFpAXpvfvKU3E46Ij90YwEWDQ2fCp5sU4cQh4j
NEo2x77RhaUdw1k2ihO0kM3xHRyjkemUdXpUyonOsc0XzgSTFpIvFH9L0l1ZAZOwflSkH6cGwVnx
fbvEHt12irHPbfYjYKqq9Zs9rElC+d4496UbphGeVAQFsC48GsxO9me5OHG9v0pZSELIA+GYpjtB
1eCvGCpjlobQVRKbTDqNsgu3+7qiDIPA82w8wToZJRuMaXCISrusmwemjzu8X1xyCE37C0aMhMPM
3X1gqlBu4TMAwCgPAALsKAF8btgXVHkLRx0ZftMP/pB2zsw9sqU2NzsewmUdXb2lLubmjMMhCDx+
vc/LbcpsqLtyd71CwKgrq8wJidVMsvD/+lektvHuM6I4Ax3XEDvRpdN80FRvEUkc7BO54dXWc/bX
SiqzdYjwlaZh+KhsuK3OR04Qa5jaKmKnOfqpTZ5K0e65KvAGTsGVywAORsjugqKSx1VXT/4AMd++
1sgohKXedM8K90MCQ2Lj3GNDBa9DC8iqxnPe8da9Tagzdz5Xli8WuW5kLGYE3dwbuuhG1eyYUpEu
ytE0p3fcqkuIkgVyJNLZcrqPoMitf/iB39VTO7/M15iFMmFXyLPQxuDM7RV1lsR4i+QrxzSNSpSU
nixbIAbcF2UbYWa+gM3Z+I8Qtv635+kIMN2vpZ4P0oiZBwhO1DmG12eM8XNxCKy7LSA584ZduMCZ
cbCJq0C7nw/laSXOnPbd2T35buE7XlYpqJ9oXM7DsQxBnCRUeGPDAK14SWd7Yu6s5AfC4VYfzrbj
Hv/roWS6/LCjPpwk2B0Vc0VaVwd3+g4RmJPXRqpl5iRhr9bXB9qrR5VCV8m7ZNGQvYBmNi6MVV/W
jjf9NZJ1v29jg4jx4Vt2TM/aLEQnddVBM8bw+mNi5HAbHl9FPvE9WwrzRGrnNgaG5n+83ncIOlht
lU0C/4RnNZWR0dEzGW+yPZ4bxRBLLzzdH9NHI6+BsEYqLkXuMoS3QyGdwFHZ4615C7ihWiF0bUSC
GoVX8wtuUCV/ibbcDxq0CjzwNzadCjfxYUnJhNt7xBj9cOG8t2at/g0HL0RR/KD1JroBrcdAY57M
9Mribklzaz6xR6E718ZgR2xT8zQDxVWmU/2NzJUBTjEFKGZ4IfJEeBsuK6TzTK3Q3oBZRk9EYPKV
fpyNrsW/PS/c3KalNl0TXo1131x1HAnZuUF903uH0lXAilJE5yjIiADfqYqGnV+mw1uwsJ2vU/92
SoTUs6LU4VTgfqSx1B7E5Sm52O6OFcYgVjB5kVyERjjeySWy1ZsY/8D7slXAfqbhr+t2AurOf7RW
VQykbMaSHH2UjYgZxK2HB0jQlfiqDIcjSObeVrSuVaAP/HAn2fQAaHWkvj7yU3/1U3MtqAFcGK98
eEgWoTbbVrUscPYP6Hc2KszNUQ7r/hEb1ZR8LNXOsk7RqRYRlMl5+jKJ2irb6di5GA51YqaJ85ff
cbuEFEDBGHLM/V2ErC3hurGrVOGM9Ve7gGkk0SGb2dQKh6uTFehcEcfrF9Q/jW2auD0kZMxIzTPs
Cnq2OFNnITdiqsOdievlZgSE/psPcchb2v4UaFa785/pd8jCuIJaCyC5N8b9vCYfgXX30001XMSW
Alh36+5YUypwrBQR12R6kJIuXaIdZTZY5liqRSXcE894MZRiaXq4IsJTTEuNwJqnQvJ47yIuDugs
B7BsI6mQ8P7nm2s5NpWE4YT9hHEJnedo4B9yMx4CF6K76VdXDsusD0bsClMygeyE3ecbHe7FJIQ2
c+PkM+HHKoFu8gDOHKIUYBWkk3C7VG+laPvOLLHJoKXsGn1NL5Pb0EemeRrBRUdPu2O7sFo8pW2w
rTBaCzgTWlosY+vCduLyWxBvctTmZfawABCylhaveVG7OPbV9ACtpAXxiGmj+In4ryp79rscSKjn
z9irxexrLKhQoueX+QKDNENld51hkscqhyCjZq/DxMPPMVfOC53MKc7mhwfxjoGmjomCC/cEwBIp
Ks9kqXoten9E7Rvbhuz+VZHHkT77gYjIwBoKR2y6oXrsjow1SmxsIHWRri1ewJ5NV+i2nQ2QaiRk
OgYqOI2jQYfhLKfdSRv4qLyzW2KmyRgpEaGsiMrjRKOZb7Ecs6pB5MeeL1n7hkQK5P0z+L7aSHcP
bNOMNPAHA7l2H2y6NnagKZ+wdh0/JeOA/F1UqhpjVEohBwsv0DzWUph7spvzEEbwM7VrFrEFljwY
t8P1muLaj00tdeb29ULHRaEDeW+Ll8jEVbxGwSXcaxSFRirmKH6S5LgAhov0/V5U1ctB9HPvjD6B
hZQmMsJxJpMVUcc2aPIc8vSLyQRM1alZbQ4LxeL94VYvHkhfcW5Kn4xQuzGl6STEfse6qyfF+i6i
iRzTxZWQt5QdXsP4xFnCtXYTy6sRGHsblXSp4rRjXh3eDI8BDrLKs0ZjhGeZLUFjd0+kNPT5EuvE
0iwj8KW4vcHHDPZ51mhaOAiyd7gJnpXr+PrI5l6pUBeRrx07fLcSGjMvGH23XIhmQ3FwsZsXmkf7
g+J/OtOmqVmQ2ESYPgmO5jbfHs93O0/F2EL5qp8Atw3jQNa/iDTZ431AERDvC6zCIbPnUqybRhOf
WCPCoIBOAIOfNcjN42Mv+c8gxtAkcejihSW7s5HxXBcy3EJHCHmZcgKem/9/Hk06314VefWRwdPa
DcvI3edWVkFXTh9W41T4FRuPljkHoyiY3Z2hYCsPzX2AdJsmhfOZFry83voFTd8uB+not10Mkb2J
NS46gq1y4K6sIfj7Aaqc+BNcn8l68WryS1nPdJviAWaWNE8u0h2Npv4zMy/vu8o1W67StfHzlQUP
FqlTDugBRixXsgjIgou+ClUkTC1TH5u0Prw64nX77uiiGWjVffZ1wCpKtHgkPMbhrUItv4uvbh3t
aEub0GMSrzUG9bMtjpwYctbJMuwnlRYsc8Sx2cHLIWaC2f38GJKgEPaWW0Fl18dTPq7jt/FQX+11
AIxPgDxFZAn5TYohkNVEpzTWyZ/JHLZjkvPHzaLX/RhOlB+1Oxs0aK0ptfug5kbH+5i+P1od5C7Y
8pkXkOHVEKOW/pH8oPLQ/SKccNqrrobkRgYlyx6IVqyBCjHshbWtikQDztfkNJGswRks4xrFOlyA
E7QHe/W4T3x5ahEHXr3ptapRQOusROguKi9F35bhhcLNocngqGupqLxvaoLPetjn+f73fZHGm+qv
WiGRcZDgl198+NAcNPhhS1I2DmNnZ9bTP3kgA0AGBAkxo0zyvouA9xKNoNWlg/v2aNFVL4D3Eudb
XOj15qa+nsQ1XH5Txd3CxTb1SSw4e+QqSsIQJc6GOpj06DF7fFFrq5NaeS5OJlOd7rj8IM+b0+Qp
GEeFlP9G78NWtb5yXtfAEB0/NlBBBcA7TRs1UHhOgCvgfL6mo/kv+vYIv8oKO/J2ddT2FzqnZozZ
rMfCduYZHOqLNd/SrXpwQchQRgmPkiMxpdavpGCpqR/I/gxWF8vg8cHzBQ6OptDMy6vZMU7RtBDP
XsbN7rc9UbQoBsN8gAIksPNZV2J3iEhjgG8fU5Bz1/5T3aeG1XyV1aZjkKKGXuXpu7+8ZM94yEtL
eHZUMlYEsdmj4xIhAshXrsKxWWj79NvkskW128D2+nAQvIERt05a/giFPfAHydqv7KSL/KwJwx5c
8jTZi1avOiuIpUEtD8O/KhaKvwMFqb+/14tca/ZhalOeWqNw/otLjDlsSgb9uyuSBOGaF2MpOxJs
HUimIjuHXsSxiYJAZ0lb5fXlbbDHinFUOnHcDFf7Bzljp5YX0ogLxJJ6EAaM4kWsVce438ltNfSQ
2Oh1ZKBjjt2RJVZh6ohdbdnhG5rCJUJcpPwu8ZbIA2xulBNC1fV48SzI6dsTAFN5i9ycFpygLK3t
YFlGw3fqAzBSQTq30meZLTehaCF1jhq64LzzrQnR7fWiiD/zjsbo9wUbtI8xFL4q4P200aHSgRQh
beFE8xhEqZ5hXbHFTYWihVr3ZMkYvIZ5IEpG/b19jLxq4tYKHN2E3sdA0InstcY2gN7+JwOvUVJb
AWL+t/2xu0oATMTkUFUO32ngDmGFNHpVFGE253YziLWp7h7kYqwrPGhLD4/yoaRcCKRE0Sj8S5F3
OUYHp7cOPV7VzvqvRFcI55XIDeRVot8Pb+um6+r4N86G+dByd2Pbh57ZG63b/0zw2F+Fc91lMMWA
l2wMK2fNVJB5GVibKrqI8UVVSPWMPv/avAfqX0qaGIwBD+p4CsddYHtjJnu4zAVS/8Y1qnnwe1vI
ZcpL/wOYpQzfPraxqztcsxlnOxuGMV9qWtKBKHw48VQDwB9Bck2dlPaG3nsUUBEHijC1gnCJ8b7H
DA8B7VWCtyNIsY8WWI+fJeIROl8AW/apxTaMROCabtStY5ke+9gGHSfqPA8x+0iB8dKbIJXRGc+n
wr6GD7HzqeTvsebXVQvjduL3XpIJ8xgQ+5cMGTT5Onr9epx3vol74q5Mq331ZlBhthym6uFvoePE
b8oVt4EwTIUSGRpws8SxfePGjnIJUt4gGqPVTtpn88E+GAUEJwubgNJDV2dFlX2/tuP73zET3K+x
cDv9u4jf+6Au0VafGA4IRj9I9srvqynhGyRuP4zlFUNlCEaEtKWek8rVhLPCLHSpdVV80lu2s9C0
NPafK14PmU88OjPCERuwmOCuwkZGLHTDxE+gpxXc3vR0be33rfVqAQ0F1irZJbGqMbq7ClBU7zcy
VFSTeDD6ytH5zmB9VNDOZkARdSOAeJvHKjonzW8ARdgu7dG+hUz5BEGqLBMpRlarVVMQ5k9lZgtH
qWhrr+bjVm2MzOvEMyczJPqXItfXpfylhOTzTmVnUqtVoe9VhLT3xVd0rXZIrlGALga6T5mfE8r3
mqx1dPT79FxmkFmoVkbBZGuX3qBJ580Twq8fyRHryB7v0XkZA8fG/MrG1q6miYtVP2EH5vtwrVIj
ffQx4/2VaGzywYs7kbM1IYH47nUQLz0V6NBPJwSDxIXH/37f+hoK37GPW7imJKfmwA2DUXxcbx7r
5XHVxPZlIc73P0Svf3Wi0U+y7zEX4xidoKnFGNdofFGtzajWq7ihUCcjGoC0Dkk1DonE26jCqrC+
KZjTXx0ALnydqIl7g0yai2/lUgzFWU0wGMPdAE6KC2S4Ho1nwFJe9Xh9Du56hfCAbL6GLO3u1W2m
qIBSYMUgm9d1Sq9VOj7q/3MqpT3JJHPxF7/Hev1yeXcWol16MaCCwfMAtKhvQz6wOvKvEWVq6UpT
+dxkiK4x7iv5kqlzN8jRYb1b2y7PgaYJ/dWvpKh+PfHrciTyuICUHT+YyQMaSuqWN6O4Y8kakKBa
D/NUX6xQJK+43As64fIBS/Mkc408lfmqJkMmQGkejnovH+j87q/zzQVHInsIMX19ctS/xASnhXmz
L0DhITvpNEPFpltJOv91SK1lvMF1NhWfIgAhaqh2iBKvTo/JEPk8cP/ObI7iIBeMfwyiXkpsctNy
vCx60IvLbsND0X9WMX1a7pt45Oy/BJyJYTH8TW0eW2UIf9RsCWV0kv7cBGFAR7pCXpYZsa/cfu3c
+CyUMeEpS8j9V8qrn4wx1ZtLpwQtJVtMtRd21YvwHc4XzK2r8AIxPR5P98AiZOMmvPFQ2IIkFKlz
SL7D2rZNc4aCeGA+GhlqaidqQwOO6zUsZB6zIO8lS0rk6twh4gQHfptBhHHB+Fzepoiqs/bUw7lN
w/rf9sH0KN8dhAdBiKVRV4KrDrRon//ADLmeVfpU20gzUwJeEXAJyKPn1K3EWUoWn1m+1Ez8AW4O
SaDdItETNPIKucOIFBC0WU7O3eytn59IRQ1aH3zfNr8eJ6919igb8oczsBeDXzi4yu3gWWvj+do+
vDOuOJGM+f5kGyIGKM+G8vYuFrfuIjG1qKUUzMZOh9CIL5KStqaG8PXAjESYNc9Kd5WujXXehEz/
5ZXyJ5ogMIIX8nUtBsSsvfEF/hsLXvoC9F68cKW5NnkRW9AZEPRCSFhqaBGzWBsZDj+OtQMjEDY7
7se1jvYxhwZhXUGfqkcGUJ1BmyVXiomWuN+Nt2rSuQ/t6guJSb7LsHH4ULXZZ63Xgmbns3sUfelL
gbYjq+AW2fjAeog98r/bIm4RahB2FyyJypbgrbGb9teafyBzXJsVaMvotkc95wpapFbukzVaVSep
N1CHMWwmIo0vOn8uEuQJzsLri3nQ8K1eZ0wp3lKYLm9EzDpobJrj1UlNy+9Ibm5CbxVvURNjPr0k
UJaLyItK3ki65D8drl4sKCEdMDoI06+nkvpDkm0DB47UYX9GY88TcXnTCu/CSWFLLe7FVL0uWavG
ZNLTvicdRa/B+HegcBNt8NforlhazI3gGOiBkrzqTWUbK0cpDjTloaI/A0KBwejUJOZ6GGMYV9Cl
bcpe50Bd/tasEagENIUuemE8H6gz2PNNdLQpRleJtCTLAUnA2l/PPrt3ybGzMedgYpXgT9HFX5qz
hT3yMuWX1ME6CBki8rrJfPSP6xZhG7bbjcmWBhJjS3ADir3vUPVsSsW8CYB3ztgoXeHcARIUlEO9
S7lgmR02GQ3N2wntgeQ+hYuCxFYHSLhGyNqdDAp94V+YfQH/OkeaubG4lQ7eAc19pR9OHtHf7K7D
/wrkWvGLkXlOt0WJol2QLEo0fJcDIuP59ayEA7FmVRma4t285Gkdg9BpRWlSAU4IiOe8iK0eXbVW
0hwtDn4L2zBxlzQcy4LwC/8kxwYOxM4st6hUxxApzz56I8X7cSLMV00oRE+pCVSePR6uwUS2qztK
qu6FraqzCd4VpyfXKWtRb603zsmd8rBOO3HRfbZ5vE/Q1Sf0ffIljGRhhd0euMfW4M+YXMsidkMb
+wb/27HvDAAurQMSNJIwVz0u+lEtpmiz3MoX5WZDTat0Os5qOb5uFmY02vE7AROArOVqJ159Q2nK
3ZyS3JcMMPXF8TtK6cb240k8BJw1ztLdzWzxlq0W1aguu7rOy/N4kaN46oLnF/5s//xy8si7jvLg
EsECQtlM14ZZuae7jA5DXLjTMJMhoVcMfyXkzMiM5pE9D3OOZi3XXLXTUY0STvqVbfxCwf6Zs5qd
/oVOZQeXEviC03NWCzabtapsJXG9QDMbznIzirej6WNzLPa41GaBwIq1iEHlz9VUDZ9rYqCJi5XH
2BFNuG0Jo/1PgmMP5UPe1BZPtdh9O1KsWk3b2fLdJCvoqfOc/7N8yCP9SKWC2ksZCXVF4G2XVL6R
j4n082tdqSXYMpblXYtgUrHcogQ80CoahBEHh/F5VpSKgObxuOzOCkHwJ7dedw1hHiBJeMs1A8Cm
voogwOg1SqNQByNo5jove3AVd8tEUx3kCFA7EztIyc4FSde607UqxcNZF79/r8G6F4nYGJmGGzzZ
+5bRe81FUiGNwwUMA4eEFDK4iX8l/AjSsrn9Pa9hpem2mf6wMj4rHIogH973zX9UXzDlyJGfk2R2
m3ejdcX3EqJJNh1TtB/yvLHlSSS+ub1eJGrj6KCa18aYs7ExdFAkMSAmREH3Trm2HXTcFw2cU+do
F7BA8O20STE2rv+jwYsfvKl+ns52mxYYTZdq94OjcD60YKAY+S6wf1DUWGOEiz78MIcZ6rIwQmfP
edj/9s8xrdZw/A+Izrvyw7d3nPrbhwgjCNxGSETaVQrh8ikNDmWOE6217tJfTcW+ini0cYAe/umh
fAhPBdhCJ4S/WmrCXI8BZ/j0TtsZ4KMc3iaimluubtNBeFAq0NOOYKDE51aLltuW967vWgbaSISo
Idmc+ZGgebH33hBmVOvevLMDsSSaLyD3Y3nEDiu7nEAQYHjqErtkPYPnh3BQMEk2zp8cfllY9UcV
U/cs55Kld1PF6knttxlIgM0MbrU3BWSowLKK3A6Nv0HknippPPDscwLCg36/VX4iuK7Z2psyv9da
NtaInRB8uK/YM+SclIrofc4nHoiLKzFZmDxoTmGDKTGA2ttWTKpmwMa95Cl6R2grMmLsxNF6wKwY
YI36Jp6d+5W4AXRpbCmw9b2GzZgeTIgoKFMeRljxRCc7ZcNF04KwWjKqB+b2bag3VZcxxIsNFsFl
4/fno/qwO0TG35N2UGK7o97tzPal7VyxA67HK+ge/OhAvNVoPk2AYX8K/KyeH6CwIKoPVcJ4iakl
RnpEDruRQ22JssrRTolVFo2Qz++S8HKoSB1yGFPTRBY0fms+hPoiACpwvf/l3YtWWWBbkDG4DWqy
64dSAvVGsPlI7QGGf5jYqQqwDUTygpFvsW4JNEvdkcHDqIf2D1c82uSRTvnVVrGnLbEKCkTpxC9X
y4FRY57M5ei7zlSSZf7Rg5l6LKAJ4hl/WcpDV5POAjzbwof3k2i6eQ0QWir41QWedzitnMkgEZ+P
IJ2OIJobUnEIIz+XEi8lsUel7CzpkR1i0u+UhevUGX/ANb6S0ino114jjTzDviazLb+91FLScZOs
vV0paLbJStHTtzJowJT62F0kO2pl8yIge9tSb5Acpue1jJJEKNvgBP5WTnkFHt4VJXYB4ptQnnMI
JNyc3LUDc2Lmnu523lPm4KJa+UYvx+NBxmRZXDsMBQ/QdtzFcd1cy0J5AlTAfaxn6v0zPvPjPxnK
Y6BxFxYleDvJhmw8L5PMoBNsEPmIUnKZnB2IP+BvL3xUDWEB6CUYCmDxIgBMihV7gE3Hv9fkiedV
fTcxXvJ9rOsRFjzt6ZCmWvn2FW2MNYASAEUBiNghn86eyJGL4mIbWsoN7PkrMpkyCD6Y89yMAVtX
wdPRJp1tifOwep3RvDJ87el+IGVy1bE9IXi1X3ifew/jDJkVXpirH1O7ScO2WCe5b2HDdV3LCm3P
ITDiDGHBOXNaWatwnhCXsXYCXTYANkHDfv6wrvSCbntc94yuTwie2Yx28ALCDs+NEIQL1hheiFs1
wtIq8Tc2ty/T5A8zAyXjQqBXH1uCvNPDtJPiTgnEjZa7vZsm9yDWWF+xNreEljp0ik9A735Ls2v3
xymc/UXI8tBrdqaYkdaQsQBf75E+HQifSYqDrsPIYvKoqlPis5ShwyTwj8Q4ZTJmxPTCzo/ZWObJ
vyeExnUea3vxKkMqSK1mj/iW+EpN+MCjQ0S3Vf4xkD0Sq+s1N0o/H2IUWehx8K8oPAjNP8S7Ohyj
8aKE1+tBMQxeNEP2ewTOVp8f7qapbgevb506ZrtNv4ysmvCiWFB/lbITiPGUGmkeVPt/logj0PWm
Ts7/AQHCb/ETqkQUed+fR+bx0jTVKiinarZl7W4TPmrKrez2jWBVt6a7TvVdO043HAFgLZp+7N/0
A8iAYMvw5aC5UtLtfblpNovNqkwCdcgkr3FdwKxxJVXmkuW0OV2geKMbgyhJ/Ly+6LXEmZwdU8Bp
PujxtQLNdUCWbxJZIPJNLmTmfTMRWdnEVsAoua8bq/gbDYVL69FBf7Gl7JH//cMeuMFflXNRJ0mc
V3TkW6MEmT2opL4SSlnk3z10d6g1oC168sPXdlFK+neVRFcaqOrd1sjqTVqNO5ZWyto+zNXHfFTa
o24yyMh03NGiu/FYnJmio7aiivuCpIIPnXZw9U/nbf7qPCpp7Yl/9WksqurOUYr2oqQOaQyypdj7
bW6/xLSH6eUL7Qf8Hy88q0gbdm264/5pwSd0nwo7DmBKhxKojpCdvK4IFw5BE6hXSIvFatxd82k4
7qG4f3vKblXXyEJMIDtwMP/5ByKyxyvNkHu0O9oH6Vu2YOpDFKOUVwSdnCr2Dq1eSEfDh2YgecrN
i6nk0gn5Fja74YwL6oMrJTa04dc7M6PybK7qTDu1gzs9diGoM+fahaVFqPf8ynALJ5yJOXKgL8wA
J5DIIKzf/SyB/OoiwIxoKX6l1V9OOeotTxD4+0r5ezUXgU5rufaDui1Z3yJ9Lc2Yg1UywJXTAHZt
Wewe33N3Fr0OUjNukarro1PGgFuooRLY4NmobhbUyNWNlL7v0jipajhXAMUhk/ba5L+xMY1rEyja
TqSynra4fYT0k4yWXYWJUXtcd2wqrU0BxHqwyxwZlwTAg/6TKHRcpR4SJP7Wq+YgZg/4CVR1uzSM
Ltbql6qOX9sLFp5FuJRy8nFeRvGprk247iaDKVOhVkdgDCnErglmBXajlchkAT50QrYnrFuH7epY
VfZ1Wyd/cby16+z72mwcqZr+x4p0NmCnjLRRytV5L1GjjQS9VZBhM16F4wdfCKBEhB5qVPAjM89a
hT+YulYoZLd4rlFJ8WJSgXxZnNIXFThwhZI3VMOQpmJa3Y0sb+pgfAtVW1PqWH6HTSOcFp7vFV6a
+vI0xhggmit2Y6kTYrYxfvgtWUzyFGibidrDR4N2VE4DS1HVxm0fwB3kRQFMYn2yjW3tG+fMsjfg
Ya6rEmVRHYUms/rswKiGOoLdsu5J/4IRNWs1ibQil4hG7MIxWR8jHQl4xBo+eGPvU1/qQh0AC2zT
UrwAqn0AHLhWbK+hT2hZcDg6OLJkM7z7+bop1KivsdqrMdhvFh2+QBleeduHwfZjKlvdDHZ5wFpG
bDEQwwx0J3m12N/wuzXb1Aj776Qw/cmJObxyJGtXXSr9wBkLS9P1RHNnoFUG4TP+bQeuvY5IPUlL
SWyuZMS51IMGmay7pC4JHvrZiLY+v0VCeKfOz7Fcq6ZR0oFVNdBRGBV+B8CQ7f8CyAlDCpjnNmcs
a8Pqsn9ge63/+qt1ZtODlNBYdmczMrU2E+jCMiIj9TGRJOPs6E7vG9Da5ZpZ99ettHR9a+yHn4Ro
7yqm1DvHvbgpB4BgrOeB4eJorH7VXbxdFp48cwh6sNbXHmZS47iF8sZOSYb6FRMlN6rl2InqefDP
aVNBG+I8rs7M82L50SObc/QBSt2tgnz40k1hA1Lw9P8PAdXJx1tctcOAPCv5EN1U0C06aWkHUVqH
KymxjDNNTdyTbGiU2qNh4nr7hMy9WCItFXpuS6kHQz+FX7DAtXYJoDhHVbSgr04kGT7BBX3Hfm94
VwqpOFOiNCCN/IHslL5YI2gZKjchIaaOWf9G/rRH32GUlaGCnDAt4NnZYB7YSz4d0sgqZ4lgaUHi
FUWClETEkOVrKpdmb2Gct55RQ07CSmNuq8mPKJT2MVoRR0t2PUPEj20crCYSstpZ9EsHBLCCtFWn
Xt1V9fv7XF/Kkl76z5f7meqifQ52hr2S2WsS3hOOOYhBLWhD+pocmexqoY5NMa/4mp1i+jDYFJ6L
00diwrq4+3qcsoqaQw7iIn8NwCs2bJGUwtROMaq7jvj/K2GKQz5GecxNSTWsH8yf1ZJGKV5xmj6A
NZ1yPa5KDZpF8NdMfqlgKyBkrobP6r6wb862RX7gzq3b9x85qYIoCJHSErYwJUIrDf1+hNQUVxND
7q1RMI/109ceHp0+VO7mhJTSOcpthsTprKtO2fE2DecwN6oVBieQajHGT8u1b9TCOh67tI6XgqUE
5FcOk1BffJyk85jYSo8O2yzjTcZI8pVy1NOcl1dmTbqYgMkCZnSYCSV1vJumZyPR2wLbNFZOQLjN
FipwVQ+RXHXYGMd08+atMySPQohMMTcNxPY/eYixtNv9qVmLRk5hn7rDt5NUY+chV40iJQMzeZ+e
dsht0aeG8E3CzKLsmuAb6nXrQNWx4cFodtLgmNo/r/soETjQJAYqLIpwLSKFUav3xu9UDhmmqdiw
9nbq4ZW8Wuaib7txf0lawiA+fSXD6ATLbigf5bboa8cpAFAXLUylC3GNUwmkXCt4moeAEaU5hJOC
CGj+D1/V9ZVVBqErky9cLGyJ8vcAPVeIsVXv31EkNnDtI/IahJuaLgEknLiagj/W/r5e5Q7JZIt9
F8B0oSKxvjsIu9/Oh8iZjF0ScQAFB0Ew4J768BmdRarnoRYnwINszrDUso0GDdqDVM/v8+Uaa6fk
hkN17TOQb6GCOfO5uehmZJvZ2gdTkxWBZAuIgEsWQEPYAdoU0Z/SvwYFxtihEbGSF0h05S/WMBOs
6/t/5ghsHD037wJTIP1dpS9N0moupRwTnlESjUQdMbzEPp/VG1mpTUcI44KvH93mVa032r5t1uiL
sphuLgxBuyTD45J/Un9CsCGM0By0iRpqUJHJPMXh9m4MXhvfb6KaF3Il8NP3NWADxeE+hME+Tn3G
S0EjYUwqOqTjQSnREh830K6qtQfZwpEW3UAnL3RCDp51qSPK6Cg6tW3z7rKM1MohXcB4ViOJ2hum
vW7yTQcmerwN3R6io2vgdy9SX+BqsrcLwOJq6Rjyy7C7COIdgS9gdL0oA/2t9HBJdHKsHmOfrINO
b2DDuIz+SiKzygfqGHG8du+B13L9NqCClYPhINm6eSJf4kezWDWh56r7qX9e88GK1H+sS/zsXjo4
XVnQ13S2F5eD1AtJ/PzdZwupMdBmKO//ll8e3b/PR3QcHzNEa3j8ERy47klNovOfMQet2uPkujc4
VIItBhbZ+6W6+zS9fJZjK2+uhzl5tND9FQVR5KNMSaV3EzlZ0SMji3/YDvWaKsQSPCBjASOSPlaK
MwVdapsv7MhgC6JRRcuyg2YnX0yGagUiKBnXuuBf9hwPKIDu+KDaApGyW5UmFto5UlQEq6sGhFDN
v3uF5G69MmOsYP3dWjEDs9k5jq0KUpp2tcAKLhEbWvEctXbBS2AYgIVIMdzMLx0uutFOYF4PKybB
BhBsRb6BMaCPztRt6kX8WrUDIDlC0H7gBK2QfV/bCWON55RLhwlK5PeT52v4T0k/rtSyRqM/+/fN
HOkDXjul4/TDAxueWo7pZbvBT7aC9Ori7z24YZn0i9IzMvgnpk3IPSzHm2sMOc6Ecwi/uTBfPO6p
pls68pl2E1mMDwFiCJn26F0aDF5VLL/XQZHzYa8OutndxDICQ/yzChwNzen0sofhc5PDtUX111KL
r6av7S83eooqAcPMFx1INA4PLc9o4dnT+D7sf60H2o3nD9c3j+YolbdMeFI0W3ehSGBbuvTSDRvf
vBrFUawcunXWoRV8f3UsGVJTUOToVmyb61SQ59HmKJIUuoGHQJAv5gV9D1HNKiIvoafu0zJFUcAF
jgdXoz17XYNhn8/eGUs+eSoZ6T8AUMkeA4cmlHVvUSwoXEgcIBj7ksuzmBXhEuAxEr0vSp8eZ3Bw
YBGxn1PBZlzekVPzR6rCKFJSnHiV+HwI3Kbz9kaDdFydiaorG6KTnvIk2iV+UCi+naBhVqQGxQ8Q
HDpOSFJLrhTlxGYnbwuDC2zaYNV3NGeF7bDDeWkq6lyRuHmeSqAhj/nffR8fEATLwZJlcuUzoetm
MSFx5Aaw9gUbhnUwWmPsLmd5cQl1C44robOay+BW2abmFqKRSE4fR6utks+dXS8CEEGaztFmqEsS
ozjz/kt541/gVFhh9kfsvpFBbIfDei7Fh3sbtRSTC7YzAaSFFG2dnF7fPurRwXPswHoqFo6xeTxU
E8vvE2Us4FESaHCjAlFnPm6HiaK7RI6L3vY1EMlGnaWQlfFVsNzCHYy+eXlfAiDW0GJc5ssOxe0Z
4l74VYs85jP2CKAL4MSOXFMAvZazwaitx48mGFX5HSivAWysNnjxneiYt0vyKaStqR51AC9Zs1Y9
Bik21wsG/ucXlw52noxw32NeEXHRra/1h5gr6CnlwNMEdzlixnRhtedYJpUNxHc7CiHbKrxb9w+D
q+UaKsDln4C6PDKlowC9pjgyamYZh9HcoZv9fpY/y+EyxOkls/2zz4K/uiUixD/PNgnA2tQRVif6
JwatWCyT+ZDfNtEbyWK3zjJLoyRaqzb+cLJq4B/SEfom1vNhI5iTEL2cSwLXdtBsNgwwYO1O/Y/e
XU99/2GFmGlg+M7a1pqVORR6kTE7hH8CoVEcx8LeRCohE6fb3Tjnhz1ycTdlpQzqU80Wi+Rbc3aw
48WSzOrT2SA6akR19X282746UPPdnG3wr6m7IhVwePI9gen35ARQK8kuKRkORd0jBQb8NLRWKFn8
SYKUwwFD9wgt/rm2AJ6Ignr4mLUHB/dCO1Mdzm7ENHMuxvmSe/zyaG3t+qVQvQUF/zTYDukOdGEG
6VCJTVKZ0NAP9N48Mlpk6xr008tZW/659H2r9Ss7JdTL0tcaHMENRv5buxqDtH2x5WoUXfVnu4j1
6IRRrNQJy7L/QpZMTho6Ab3WWR+HzRU8hNyaj/l3MPcWLVerZK0QPH3nIawwwnDn5bFWKkukQDWd
dzfyuK3YZGGZCswnuGGYUFhb5p91xL7z88BeMzPfSVJZ3pPaiQR9bw7gwTdPMuJwdXmRwEoFKgr3
Hzw2sZ9IKRPnkwV8yIBoBJZSHzjw2IVFKxWNTl68ovP838cL8Z5zReh7YB95gRz6Edd7DM4zQE3R
6Gk5fck/kw9gcGQidTEMnZWudzx82ZuQQ5IXPqoYneLhCsYmzgTT/w0tQUBikCumYPpYIDkfP/hC
L2QjJ/mKJxcJwDvdKwYZ8xvYQaGTT662Il/2rjkJEBEqR7vPknJ/db4CInD9h7y8QQJjWDJy3EGt
1bOciSNzBnDWkTJXMucmgMV3WpWD9LNZq4O6RsUEVoJ6/b3Tc6K2aOAxdt5R/mEdKP8MZe1KfdRC
DtLRaDaeALvdhyLYZUl2DUmlHZMOx+JI8qYBp+e0FnUQiCcAK2L2S6MGlPwO6ULFjDezdw/i/pUH
F6WeOifHsVvydKNEz6ig1PK8UUvbsYDiETLRnbZrTQdshxMygm99xxYUGRigAoO08kR6XMFlJxyq
oGiu/pOhC9s4Qtfb/WvHtOQjNX7pac6eC4byiLqEVPntQH901d0EA1aWQ4FCiZlp0lHIgrhx1YxG
kgLN4S9AT3Z8jiX6V6R4OzYeO6UpUP2uQU+u60/YZ/tw51YCj4ujg4Z/TrSlyba1yzXU1DKVGUrM
nsRNzsNejw/Q1GhKn9gSldcCiyxoDPd8BJVg+ZRqyCFv9vJl+1g2CHdzdJwwZw2fntmNxTP+RD/f
01/u/+OoHbR+fASLF3WgcExF2EB2sbtwIsT13NDFWhBX3ndzZxy8dmejENA6w4tMV6yb7ZucvIo5
5JHopDDGCEiI5ix4mGsET/4JSp/QNdPphkrmPuqR/keRdhrPskqOJNiRItflLWBz7DUNsu00T7fm
+/k5IhxKsIPnr175pwWmm/QqodV2rFpX3nda2aGWPWHoPzLuaatwT5kN3bMcixVfHpCwVzSt/RrX
KOjaNl0zCXH+n28AhYovzYDo2r8/7KOKQNTFyuFbFhmnDAh8q7Mmn+aNTJqwUrcMLjBOfgdXQ/y2
0VtdZSBD+fCktNuWGkWFEQ2ZuEoerQJrfxW99RrGV8x6wp5IotOJICLum/3xwzfl409PbffquB6o
acvxgz5msxmcpvVjaakfqkGaYlgaQEMGjz+c4lJ4oK1YrBw8eLzJVwLiKY9wvoeQdAw3azdgX5C+
UHQrs0QYEjvbS4MRRTzcqnj5++AoEm2g+ueRMSNVx4r1Uk4YEYxFgWWklw9EmLOzFnzvZJsQsQQa
tT7vQo9BdmG9wnzRhwDt7ui3mRLDLH1K4EGWTfZ602lOv+4ko48UjLJhrY/cdrUlHS25M+F5hh81
HkKPX7mMFOtAtfvwrIqwzp3+SWUJ+lb8JTkH8XTldgQiftifo5TxRJjVnUUek4IUGJwRf6+QOx9y
mY3eiCVd7I1FUxnesnTkG9QKi54lh29PnEFju3THvGOJP+aY73MmFQKB/PDFWbAd2lnYlFa4pMlc
YYhuXyliAWH/DQx5dNgiTJvj48ogLLBI/tQsAxxfxoxUuDRXUX6JEEYWlBvGPsFHaQ0O2jfGYnvR
6OECR0noB+vSVZLWlPmVta53+zNkQ0+tyFpyXtB2kxml+zOoNDwM5gWycweWKqpmwLl6dwfI72lK
aa4XnvYrw2P+uJJ+lppnCEi7ZKu1w40SEj4c8sE1lXfJOtcRSHM/MCW98nTb30ZL3B3sc/HENe+s
VAvrVzhDxTjsmOgi/rTpw96fBjEYgx2ejzE2348O7opRPUg4hDc6M8VbyszeErT3uDXta3ZbMCY/
2fq0J2s1DO3SNvtxSPGtFRon90OAKJ7caoDkZwbs0o1dfougYJMNRdX+ai8Xdx4wQyJxIw/59SWP
l3g7jNjuGHWUdB7GD/06WSF68blQC4M1Y+oootrqeiC7L+y9fff4BrGPEQyeFerSBxhtW+0IfthB
LJSWxTx8SF6jYoeLduonTlG6UyyllcJRhO/hKiBGqcqGbYb1vPR+0ZvPhaX/UaC/JobiC55sPmsQ
YqpgJuvfWuB+IWe+kGxZQE57bG9IYhruN7gik17/cFd28Cmpjl1o2snnOMt6p22S53IiMJsb0k8b
61LsNjK7qiIwlEGRfQXbTLJJGqTFJpsbleFz5u7/kD5KTJvWTyg59imgMOSa67s0uLB4OWmNA2Nm
CIz60XJNS6rfhFpx9Sl7EapOxywORQZgzZAxLjCfBVA3+7SO6G6/DNOvvm9BK/qaqRHkGmwHA61F
ElUkcWUJOXrx6PLaORBp0Qui84mcji0vhp/IulwLtJ0EXIPANDnUudULExgTJqj52H3JMz9Pw2du
d4qdD1lRVq3aiwEHbLyTlo2yWVdeOwJ5nD5x62fJJKZ+7P4yfdlm+F0OWgFmM1vjduRHX6qBxYnZ
GnLXwpQUFOK+PdNF4FFkU61u+EI3yQ/Lhc8Zpqx+KzSTI9/2xcmpuyFrIv8hwgpEqY+xV8BzVQv6
fFjNfKw2WpyYrXJy6eKGFaFG7Sb2sZoSSlffN7MFcozYhlr3xEN4BQ1mhMUkDOwOLNct5o7BP5Dp
gnL+jMTv1cC4sArpYaWFB+2trMUsln+5QdTVTW23MNq1knrI/3z0077vpDqmnSumfmPKspSndwVR
nIdB4J0kdSpLw30yHytYo74WFDgYvaIlDUhLHOv/kVWCygoFmg/ABsPFyke/Hohp9XJnhSQIsJCe
FFS2wcf7qo2/hNkbOh7pAihUA6x7X8XbDdZDjJ5nnWzHL4R8I5s/R8Z1nWVmYbGc4gA3YkQacmvC
cQu1I5wAheZ7PtE4M+fOG62pu+raJu/6RMaSpFulNGdLodrFMJTw5IMZKeJd7Lm0gNaQzeEn+DPN
qL/S2TKIO2fIgMIx2KQN7z4VQApZenPCcjh7Ki97m/FNxD6PH2mCwx9KmWlPSoU7+/XEvck2u2yE
L+lgfcru5pLf+eYWGV893m/aMz++HlK+9RBiZHO8E/UspoIV9y/a2q7sgGnlTnKe3Nr6QfOQzSob
0dIrl3oQ00D2l7b3au4rMAoQF0XRYZVFMMihNZQuIur1dpIxo/iUcRtcXMxCMwnAsXkwojSJZ1eX
kwYG4PSw+cYksUsX2Rg756s3uDT+syLRugoqxmQqDtUBE9fEhK4sBpe2U6+LdqBlVN6MZxZ5TetZ
WlRrzZ/q4QwZQFqa3I2KNtE2ZlUVqiXRh0Db3zW2Fk6ygEXyH6d4gDHz8564OIJdT0gszlgTOKck
IoEB3p6/ge2rczca6mpYhXF/WMPjYtZ83yTMW7/NxC4Yeqbdf/6rPdsDXohcC9DSykv9KZPgFPtc
ZzsN9pohUGReksKnSgnHnSk1sZ181vPj6eunoofGZINPNWE1bR64t292EuWbFxHFmIBYRD5kiYW2
CedICnjLkhRpAOYrrWa8rf8Jfqbf+GwxNszvZSKMEDpeOnJGhitZ/FRDo1yadN2b6kjyOOvgMKLG
oT+iT8PNnXLEB87Ykjry8cOpFB/nacanIPhaEqGmP9LftxFe+cfsYGzch7gGhbomX2ynT69ejVuF
UeRm6A0GPWQkK+B2/yA3BY9G7MtEogv/jm1FGXNT+tqxMo2a1OgtIJ5JOuR4JCrUNSXuwuBshEee
WMHYVeGkXgSwuTqxKKyEKZwJwaBqqFQhmcqsHsMhB1PuV1qtFjEH5bO8jYt4g6Wk28MHK0GYnyLB
Ijlwbw3yu3v6nq9X2JDheUHBn30bk/NMBdWQw/ZcTVWr/H1pG4TmwW7EmxStgVsylgvEB9d9zcrR
wLU2AYvrEwtfAMHaI+c7O/iRdApp+Az+YkM031nkpVayqVK4Nfzj4pTZMejFNQToG7vj7fEt/MdZ
4pu+Gzqq0NF09OzidHo66S0LS/elYjgfzgYiVXqbh1OwXYp2L4eavHR41AxFJW9ITu7IJD/UiRRF
KtdR/UbwWTY9P/WZDbO8er9OQ6Alvmlk/7jw+Lg6WhIeNuLPARsZmOiqpUqbkDHsr1J1vaiTocBx
3m/xH9v3+dQ0szrvbdCJB5LiP6NWwPii+Bm9KuSg/zLM9JRLpNxMsp7d8pNKYdLEsFX8c/ivnhPH
qU3AVWTk3Pv8V0KXd3CNXkakkRKLfUYfpZ1DFaCs1P2V8pR+8hcG3JKaYb3jKyIh/Nobh/F+22iI
2w6eDjhS4HfGcD5hS8a/s4GeIjAjW2HwrTAIeN6y3JYOnG4HkRabiCZyGOkiq5Do/6DB6N/0hks4
UVWHAePwS63tpcWFN6h8gpfCRGbldK8B9NFJEr6v1kdCLU11BqF3WkKWmfM+JWLSvx+CyA8Z/WR+
3OQioHPr2cm+yU7qwb4n3ZkwZmjhm0+cnRKE5wORpVVyoUHw4nC67ShSvYeetkUzXKYZCM8KsJdA
RbPm85uMtHU1roRhdOxO4LAVDoUsAiQbUGufnvA2qJrsILeaGffVAdXqUugg8cD4t7feAtjc+41+
RBoJG4B1LsKljDfKk7vYmZcWq3nbD0rHcwhbbGpCHEu0hbYXAyVn0K1BqpAlMHMyK2/7EgdxPzVt
xhx+67TEC9fVKsHvn74awUm05WE3+2xAwVzWnkT60mjbAryVQc9Npm4+K0Ga8sbCrEaQXMN4slZ5
a0iFqRTuev3iVF/Z8Y+NeEmSe1dXKbPdsileHkHAC6GLoVZpCoQhscP7rS9jINjryGQiqz5hHyY4
uftF9HZJyelvH/EnESZVlWZ/4jyvvX4Jm7VhzNJ7NyhRIkPAY84JFtgdr3ucZwO6xsbaNaw8zTs6
46ina8Bg0oHfS2RUbtiB+xV96YE6YOtsta2uiy5+YQeQgFDXIfKZ8wXwvVmmlUncOZVk9UWRXYnW
Enm/rBUjtKk2mVv/+8Lbiky8AayOVfaZGMwGJeA3Xy2QJk8QGutCi8wZlHrB6yIHPSBZowUp86mX
ZjghqjrKPtNoGc3iMflFC4XwswdDAXo1j5v8K0adz1czcMPlUZJbUR4xetgnfzRjGjenmqQA2C7W
3g/KS4VUnAQso4+tn4dkc81gqvRj6iDf6c7guQzJAy/T/sD9lgxg7umXcZFRF02Z7L8LfJS6Lkmr
lONqb/IGKTgZpLgw0XJDXWRP6jCtXi8wc8+g3yTOL4frX+CZk6LNVo6RoA8F1r9hsi8g5Y10TVVY
iA2c1n3VQDJOgOM+ShmkFwHEjXhOo4bgfJEM2JhnJ1FcHisroImuTxQyA+qUhe6l0YgKxMFS+DjX
mf/XmTH/QCn1CadQL3hv9ly4EDcZtHV3VAakGHCSuo5zxBgRoQqixZPz8XeSQhK6OWY9qqZmhXdE
1w5jqghKEzC5UcPJxR9Gad/uOM30B6GmY6RyYjYddpsdOaQtbQDEiVpPJ6n4VAqnXwg9pcNBU/ix
auPGKGikMnT4YJgOhc0R4p28g/RmfaEwTk0jQ8G8n2Q4YbJ9Jia85QeXNAvuzh8TwJ63raKUtMkK
m3geAuGj3se8kS3fx2EH2z3RmJH41ME7suDhX6uBWeMzdMCdqLDJyAi6OIP8PTqpqyKkz7ljtyua
ZiaTs0NvtQCzx6XMYM4it88d2wyBQM3miELWXUFEJhOZJyaHo4vkLoK6uUw5c5UriYvs0XN4c3Ol
BA2cgzfjzCTm/WGjTtUsZv9cRPaxCqzWVH4Tl5+jwn5QTafKqCYfpiYkcUlFkUzqxn3kdXUIFBHw
aiwjNnLFRlEuHxl1kx3zeVCUGUJMjZnLbLkaJxji2u3LiXrZ4+ARE71Tc3Y5cwd88NYNsLkEYFgU
1quagKOf0XH+5aXgSkSJ5FI6+AwHzFwAWAIf8Nr+cSN1Zm8A6pv1FXa/ULOnaBqstqtdKn95z0gp
QgsUoIG5Bqb2Mjc9P8TqI8l17rcnWWu4s+K+vF39Axze0+BP4p/cLeYstjWQxtluX9NNnSb3UeYT
Efiir/g6lwJxqjxeXYZ/EEhuV685d4OS9tMtpdJP8koXTnsIi7Izx/4+2BdBXazxGYqH8af7paJr
cnUarKmyS5hcPLJAbOetR582dbzVc4kRlRoTH6IAb9Zzx4H0++a7nhrk133JonYOsKZiHyaOZ4ic
3pPrnqp/9xWoqIgncjJjOTqCjy8zGOqQDOWk2jyVROWFyei19gi72vReG9d6xNuyN18PjtC+5ZUR
e8fMDgI4UZ989wINXHXJGAEvjSc6KvfY2b7HS5ixFkbnsU2RLEYasYDT45dsecok9F+trJ3Idbhv
KuCnZMCdQ+2U832BDPwqIh7++tii2f2mNBz8c1EzzIZPRIh7FqdNUjSnwIfdyG1iFpcwmfnntRbh
haP8R0uIAbLH4xdfy20D/gU0N2PIrhjV2SomfTF+2rXjYsREnwQu5IsMLH3yz79kO49lVHRlwo+O
43zpNW5Jw8xvQGv2wV4+i3HYzpHCghfj2AU2NqPWBGuUU9zk8WiHeF13FP6zXRDcqf9z/z9DhZRq
b1HW9YLizKIakTdeAE8lRu8YZyZsRh8DwW3VnIag7YKh/IAQzD00IB9a2RwYDXn86KHi9XX0g/d4
4Z9r1U5//DhQCG902kZnB8RTAlTNCHkYcHysinUGyOsr6t6s3CLUgdgKT1otqGHPkZBRkglbzGdv
m/s08ap7ncnAuwSKi2bc9tNypRTDgXqMxWnWTG/ZCGGzFrFj0FiWhFiF+kMiVyvdCkP/wrUIjfeN
jL0SpmWe/P/urnk9gLwg9LCti/7H4+u7uclehJpa31F3K2YvwaTohn61yFzGn3dklbaxf3ge5e0x
YuoG1HEIzcXdZWJ2doTrGV3q9tBg6rqu/dJvWtdI8C9r5P8NTs550TSxMR36FGa8A79vw4rUagEp
3bZ9bguuxdGynOQMvS774bBhXa6/K2jWyhbJ2/nmYjqbsn1WgzkRdgLFr5Kw/v2SmI8uQVSRD/mh
uKFzIh5gY2O6BM6lhZn34F6iZgqcGtaZ770wqSuQI7svut+YYKIOJAsC30SFnc7ZRoesgVOa0utf
8hh/Sx5pcIPqTi7sWuBKHxVwNtjmdAzqRCkHAsuk10N2zKRr8HH/TGFxQ/QHD16MHn5+8ZajU4gj
lO9YlEkPgpA1XQ5uXlD9WBMauv3WilebJBsGdxmBOWuKaLNsVCYFC+Oy0unNZdRP3dAhoFtN4eEZ
I60R3ZTKA/sP9rfD8/r0m/84lW2ToiQggrwOrvhIXXpLMakRbivMeoUT5L2L/OKUPeG5W7KSQ76r
hci702ONduv6FsPxkxmSNE+nVqjbccWH5ddglNgkMb1qfwejfcsBDch9r+ypgsnJgGr4nP46cZy/
Ti3O3bKKuR38QH7P7FZ3i90/llFMmknSdY1FgyCYwINhzFXB4ntH6OKLmSidqRROrXKoei2w+txV
UMP9q9mxKcsix5viRP5K5yd0jbT4yUkKJ6NMBpDB6Fhj1IKnCGp9bV9peQbnzcNL/PRniDyrQ4Fh
+1ncLpwol7UGTDdG4uqgyziy9GYUelb7my5UTTtaXbQd+Def87A8pkLj9DdVjgJWbM7gEYzpdH+y
xolKNGvYWAw/EOeZ3uP6OTQcZLYYzWog4wuRUJHNzfFW/MDuSXqAvhc6vPF9oHjWDSBlHrBT/FWP
jsbQlFvnTlabP9EiLzAv+dX6ko6zfeIbt24e8BoGDngYjtIfrSzOnV+iqho307eLP8cm9MOhDWkk
Xc8aJMaXpRUezDBkVNo68yPEUz4KekF00UKP5pTCr/kJip8l0eODJp6Ned+8qNzmB1zeyEJW4QB1
ge/n+GxX6mnXLwKPW0DzZX45DTMjCvsdenUEre/nCnQObKxUop2BZJneuSIKR0L5hvKZpjJyDdVw
hK8r1p6q4bRxPSk9GcWK1hXKCKHA1UTypP/FizRYsi8oYyiEKV0fQ4gV6XpgjGnf4fV3dtmqZaS0
ECiFxqx2qtuLiohXsx5BB/gGRLyOMIlBetAzobM9GOwJqvgmXU/pVdizd+Q4Z1b06yX+8gx/azNa
/g8sZU+01vPwsJOs07ng45xRWGsAXHrqt7q9MimTJF+p42bL2W5j+HmfNj7lBTb54FIwJDIz6Yfd
fOIQPC9k7QX/jskzTw81nxdddp33LCdnhyxxZQ7mKuJr5iin6IWZz7VKVbozJJz48EVY8NNHEtFX
pmFTcMdHrgNy/zXa7jGpPtMZD3gwGrnyHzpN/p0friqamlzwE/aoC+78ZD+BdkfpvOs/HE1SRwIv
vdjOk/abhBQiN1QjVqOLfnhxbAYvOQMj7qsiGComgHXU1++K1kI3jlf5u/UbVDIRcrsQgWIQv/8P
nX8y9CEgZOSht1KNtVbMTRpPqkDGo4c/KmcPWQMENlTyY8qYSLTH6OAKrUexB8LewnNqEnq7CAfs
RGX6BI+vzxhGygYmWSJWRSmW/zMV1djVzetXEbBvNcrJchs0SpZ/K+h6LNTn6c8B+eV4hx5+lzeZ
J3LSuz7ys5T6SrZX/iAvEGtRG9kEZiwRrFRoTBawMCp59sTde1JJAXAcbNbRGnneJk5dxULgE87k
uiF/96n28y+RbBEQL+qFCBDEB6M2UXvrjEP2dJo+8o2dvzC1z/7d/z/W5lvgSA9s42/hlqNhV57V
tDaPUGDcHLEettZxvks2Rs1dXLIgeEzU2PlxFV2iDs4bQgakH/P7+yaC+ZI/ty4UzR00cPWC2vZu
ot/0kLCt8cT6DnoV+W846rV91NGsrJ86kjvdfbKDBwYiddlFMCxNzYjqAeEmgZEapMYjhmaXETuo
2ai0xifJQ3MsVvG9eTQlViGdZKX3VvvXZVnoSkFrs4rVevqyAtaN5gSbcG7H8Gi6aJMVH5jgNCvq
W0Na/DfkTanPSRX7zIrJmGpjyl19jBz9Hm18xiA5J9QKsF29rHffbempJXvdM2c5Mh0WeTJXHyDd
s6bOSfnf34+e8rsMUtwS2au9CzGMHCSw+xP2A25EqKniTUeKuBB5s7am+LMaiw4M3IeFmBwInWMo
NJ4ehG9hK9s8fVdD3++xhP7rDFObUAfM4ga5B4zN/5GEWP23H2x4OI4CznzYVhFXP/chydl55uOY
CMX0O177bUhN9K4J+fnN5Qkis8vODNvG8GfafMrXswODTrEIKRgiA8AnBOyBxppwyTsXALL4Znpz
4IIMJii55wEHGYXGDBb+WcMjQMqGSwZKP+x/iPVzWE+vV6OK+yx5LDTefevhKz8KbYIN6/HB5lt/
b9sySBb2ncSBGF9nf3uE/7+nnyyzU/imA038GSyYHLmbVcCX5y859ZxnokOnbrLQ/xZg88PQJLbi
Ezlt0VebiIDzmjz4tWjWTBzRS9Huk5qcfKIJQVOMjGyZueGB/j4DnyPpnx4mDWzLB0B12fiWOMf8
t3BByHB+1ZFMiLvKJEoTfrXS1WPfd6bC86lrGE4sYEgLk3tkHKCT+HcWcpqasirkGLp8W3uoEj3A
89l005M8j5FuUs/cxg+wtFHZLxAhqqDGUi9oRLjWZ1j2L0TJVwJrniAjY0sZe8eGt710TYr4OiHp
hMMLndgzCKnJCOip6E1Eex/ADBpnFpKSFG137/XWOqju/v0phNaMl4k4bb/ZnIpsGVDsPvHMMIba
yDvWmPf2wa/FLft9kXw53uMWGI/fAmTG9RzrUTxic579pjQDLw0OjgytBi3PIoOvno/q+xmcrQ5C
13+PyZAU+LTYLyku9Dzp/RVb5x6jjtIqG4uCq4nP9fdOaKBXCN1kzK4B6ZRNk9QPKXqzHjSRcrXr
ClXDJxzRZp/gik9xEmxv1TTVMstHXhWwGUT8Azlit+ofgH8NhtExCq6laOPLx13U0aiYMVJ+V61b
++NIk1x2mR1k1AWWzZ8Me/4sQ8wwngvs1QaJgT3uEj6DDZSadBhXAftlPxzlTwAqrggoqxcQLjnd
Wjh328LUr5h6otuqp/ZryGoABB1O10D6GZmUJ6xtF3AqWpx035mslnct3iqN2ygXsg6egrBW97d6
Ia3TpcE5oF4Ld1PQQohPhzHzZdx0pl8G0LI0eM9YJVaWwTqlq3fjsDfOLiA9tUXHb3Jf+hkP1T7W
RpniFCvMxqxctw3y4gVu/5W5V1wrokpU7hQDUyBn0qNgLZ+hHvfIeGdXf+kuntYGC1wo9Ra3ywch
FVnNPds8+Z3c9vIUq8Z5oVtIx7sDIsw84vvjIY3FywpACoaCVVwqYNsMwlFS+UJgJBUs9ZCIduI4
UTrni4NCTtp5Omgkro1T1LgRjdRRZixVkCnEnXqUTNYQpK2eW0ru92bpfnbjR6J6nxvLvygV9Wjz
3WFujlW1sdRUtS91v8EkrIsCbmW3NWlV5GHlJD/6/NIkdG846dfMP3M0NGu9TbPSfJX7Gq9wtmoo
iiXqGUn+gxSneXueUT0AoLVs1If0ygTfcrNARigIBURfRThQ/afig92N3EnIyOKgXqP2hM5wpbDO
4WFjjD6glujJjF7tnQfJvLD2GDSCCBeV/CpzAJX52F346U14dV8WHDCj8fE68MzU7nqQsc0uyum0
L7FuHSaeNOuScOxkmc2/xyelrRvLzob8b3lNH3mCHC0ojYY/NbeM0rG/gJCNNpTb6jq3C1+wtLVm
DsP7fP9Acc0FcdKhcTd8h87E8YIgJrZQNty//PaomlkGrI4gejKQxuwY7xjJcehXS0pGH9UQUDy9
5roUyMXWc/zSH5IELXPm8Kor5OrwCiKa2NH3RZOXOQp9W2BTIMY1D4Gk5vQhR7/CiTgksMZPb7ci
nVyjUbWv+CU0LRu0Gzh1Tg/2ZJJ21To7ks16kJD2Ge7IR3keYkzLz7BhUJq9IeMR7m2/ZpvNhtYw
zB+Hf0x+nzvDyXBaaWYl71waBB5fUA0VclXqtvXAI/tajW7tPOh8XuThni26xjZdGanHyjifATw7
eaHP+igudD2FRAScKpHhADdtM6TRB8wIxi5leT8tIswbvDKfiji6ohgUd+v0+M9NclwIlVjUinWR
dTowtqIZSeyuqHLNDYrW1TNdrAG5h6jPfMWtK+LYWEhtgVhz/zT6zGxMvRuYAii1GmofKdETvWm9
54nyx5f6q/M+z1LttEMHQbLj0K03V7lIW2P0wcBfSvn9pcr8nvV/GQ/2EzikUDeueE3pKAoDvr4v
EtGRfm+0YAh6cwEaGyhL7Cpn30dxkpqt1bBPqp2iEgfEt7TYm4re7aZQBkszyJeRU713tfxhgYLL
gyDXNqgMFntnXJa3VNjqq1N291HeQeDWbqxi8enQ8ZRmXEHwr1qfhADd6Sq++bf/R3Lj475NzmbF
yhJ9PV/Xsfa9XdtQPrjrborsOQM6oiPxPM5WXQTUuxjCxmHv7em9CMUhh/WFW+0bNmA6hrp7t4jU
q3LIMgLjQz4vI1+8Gu5vHMz8vHR/M70oAVqK724XkZ4YL3SJfRwfaM0frh2EN0JqXBmV6V43CCJ1
sFUkyxTzEEbxD7nwfeu+lOc9xJQd07jhwXiDzZRn6Z+x07Izy3ius4jkVh+PotNpwhh8+GL67QHr
vhCj9c6zZjiGbsxgKl0t9pNoIPP/XJMd/6abq71Yd+jYZFpkpgW27tNsjgKVJIj6nb6tBsQCVdQd
7LrsLxCyyFm6MVRGTW/34SRfIixu226rJFA+Jzb6406Yz+rzhLQ7QPBWXdRvWVtkrGl0SSGfeDJz
rNnY1+xX6qkQirrZ/kGtUor7hgOalnF5IRpzS7eM+wy4TQL/eHcvc3VEIUTgLo79QzBiqOrQLXKb
sXh6h9VHxUNzB8DqRGdR6QznJqrEd0oZIhdjtM+9nVhMzXeJX/1INy59rbxzCXGIuH4MAJxJYqAi
9EBeq87XNCRymBVd3X7KBNkMIFw6hiGPH1a9C6I9uZfvYXJdjwKqnqxgdGcpVtZRGulUDFg8hLX0
ydA4oFB9cc8xVdOayqbOju2DLg+PixymYsqCeXbJic55kNUru2YQ8j8nmTmJfFhX/bhpqaT5akvB
o2BwUR4kB5n1m3U+Pwp5QyvYlkJp+EKMytHC+rbCHLuo+R14+RxzI2iqccQAIDSBD+Uama3YYgv/
X2zhVvCuFYYn6gneB9SLiwVUTGISHzYr0obBg6Pn4w11AMqcuTNwhfyD/QY6hmcRc+4Ov1HdTwnd
/LmB7tO/a9K7HpTJXvUcwn7TCFhmM89hUR1iYK5tfpyGObPXNmsupdelihYCCqVqGmlETJSYy8Ub
oSuj+3xtSmzHBr2k4cPzxNnNrp1SibhTQyUEbUbH05WctO2FRDQFOF//GgtWOIfb+j0/uJ5LcUOf
aq6XY1IReGF+qq+exf+qH1HPD1t+G3awJ3gOBKa38Vu/VZVS69fJ1WpEUfHQW6zPE5BovK6UGYuK
FE/UXcIcmbJ82eg/DNz4PU1z3yj/fSlZCJydfm74ltMxHUuMYLKc6NMlHSGf7mh/7cjK3b4dlOvJ
qpaUdhEMXKtNw/WAfQvfcdZNX7CDfIMQxVy+J+eqglBqa2dO0bAEx/cJ6raujn34I9KiLijwHZXS
asqrycuKEXPdlHrAJcpAxYqmY3ZpzzjWqA89Xa3BZ1BEhpjRpSLrED2w9T+uvBkOQWuIl3V4JWDw
j4hdBEGrQRRUAHFk6OZMpN8J/PB7AzSOeOmNAgCiKzGESnFO1hgtK/D/T6hv6uxGZ23UearoCntG
rKo2+KEPwze5ZhRF84Q2bS1acuN1Tjl4LjqxLH1WEnnNfJB/B8zl1vjM36ZXykpzTJ9ZIUKWg0UV
YgnoClImP6yFm2tTNrUzLsIQ7p6eJxbMZXye8L97cSYDJ5eo+GreDTvPGyebHpiidzCFbt9ae8At
xCl+9hWHY+2KgnrSbPEAhAgBxIWoFbDsT+J3cNnf9UnHAHSgE1k+z/05/TBTnQX7CAeqgdp48Zi7
w+Pxrmgu3lX8CutUy0o+LjgYFL25D7Vt6SwmzAW8TsViF0cqrHjmPlk5gOS7x7toOtIxMqBloBOE
8F0Ctc2O/FfsmJ4v4C7W+fORwZL4hCL1lAMTTGyCgH7Uv10TJmq09lN3HHLZ2Nh2xjD4aY68Phum
GYI86HRcZAb5hnoJE216K5eHJHpEHHDciUnT8PcCv5vsKDJ51RPHIW8qaNL7EfzGw5B0iSzsIr5B
xQTY3hAWXk74D26PZhozVIoTZxlnEd0xJiNRYJ0AUdGYE9fDZbmrTxq+070D6NBJLHjCG/BNYv1E
Sums6r8A3vCOm29c0cYq7s+Gu3Ayq8WC9GQhQRnIMc2itqWg1b2zQFK1Hm5dRkWXh7oWADX+54XG
O86OTrmkiM2YeMRdAiW1dPuoYNGTko9Ue7JlnKQ/JrmrmLDNLEHKhimzYwRv2Dtv1OhfA65mBFZs
jNQL2ZCNf8umTxRQzbu4O3qQELaLgV9nA/WKZp8BcmfvKxPaP8oYwhaKbALF7e3zSNSzH16+fhvy
AOr2gYRqPX1yLg69TGGO4K58B0hRDMsQ8vAUFG7x93gOKC9XHIWMyPaRLJ3y2BgbJTdOYM3tT7Va
BgEtuS0HlIrY0RiG2LI5UD71fOiltvM1fX9kkiJ4JT34xWMt95lhIPgNBVLknSbFrjy7EoocDVF5
GDet8XuxtptAu3UMCTU59cp415Kwz5M4XHMAm6R4WPP3Sy/3vWZhluDskTOZDm37mOSkDvazxUsi
p3Doc+lNA6KrUOXkGL3RISVqZpP8AnbKvOgcyQkBNOi2064Xozg5dIp5fwEYsG8ymswHDv7G4tNT
i8+Fd70HkakIWjEYFu8TnjQPLgXeFOF7dQZNt6xS5qpzuALyWIaHQXtLOHxdE2MNSiNRfnk7Lhko
91dI2l12RbZidVT7q+Z++5ujXDVuYRzItmkuMLFcdQ2hvG4NkW3+mqtCRLV2wKZc2iGQ/HNvY7Ta
aWySxfsuHIjV57hBkdylHGkx/ga34bADsRslaLERLucS/YA3oOyNPmNwmVVue6JZ+DjOPJwyDl3I
UYcaVTxnx9hk7UoXqDmvMTKItBaVaiaVFUN7isRLQxvDBxXE608jz5UZbyInvZrtNzW8T9hxiNzN
5GIuGOVtzbNduUV1iIFUrSH2xf+8amK56clD/6i7j5Wq3iwmZFHO54lWjedw4tWbqauXnKmaXNBv
iX378WgLT/IgGxaq3ggHO+qpEh1/QnVbpEYlf8uWPrl3aAzVZkTEEFV2Bt3A0P2ZvuWDgyWDGtox
2aNKgsJATKuOsb8a6dupoT4zaEhBFG/f8KXXQk97vEG42+lQYwDeog7mTjnxUeMMubZ2qoMccpcI
27vy7U0jURK/P9p9GcNPVoo/Felc+HOamHIu70JbHMLy3met7Ey5wdHcgTjfG+9jchws5wkdf3ix
fr99+wENmP+dZi+BQkmNGiK8Q7xSobnx3lQv8m68j9G0WUy+k2jLBu8RQLFkPWaTqKDNT4LE49f/
Dhpb2q8OCycIreE/sdeTbIhQ7SVzkbUD7nnCUCk5nmHyiTRtzjem5qkIeWKYeMA2QpM6P6BJU6vQ
bAS6/pN8AWoWtNgcL1H5ITrZtcOAQpYriAaauOU0O7Sm+uFe3ULzbPznpuEDEp92vkK/324MIjYw
qyp8sKZ+kNiUmf7E9jilldx8Qbx3Hpw2xFjwxiVYr1L9dvU+P2FXuBaQvoRIxI06R/BB8pp9j+aW
Atq3mAYpIeMlwh0cOZ0axv1r/kGUf+C9Hq2CyRHIAIres2eYZptloy3ly2VDArYNGUbmayMDVdXY
uKjjPovAmAp5x8nstOXliKbnlWRNuYKNeCNELk99D5wiYVjSRa7gYYYZ5PXIywrnuCU204ycTdQ0
G3OFrW4m38FLJgbIIQ5bFO4ePl0fqlgmUxOnyMPUOwyOqslTxuo40W0kfii215cb2xzhAHsb595V
tq3R6hZI9xUp93wqO40GdRTDt2s+8L+QrqCgp+ioi7vFlk30+W6WXP478bYD/2fcy2pC7DKNOJw4
AjloYvf4AXpqWdv1+3QtZ8sptCfmHUi3e87dlFd5vcF4C/XZASLBFhQG5z0tzdza6kHa8R2HnsBo
rZ8Vo9Y9hXKWV0QWY+Kokd0xI3tcdW5jJHC/A5trh+sFsJpgM+G0mRY2CJq5SEfrg6ce9D4HTgrt
HNnNPWsRAH6jdcLo8uoL6OKo6D3Mb53A+KzHKw9lJo21E83oWM981X6PEWzsynjuXon7IS9uWVTJ
eHBqSa1SUnDMBXXpIfdaCk6W/mty7CMXjmSXHKXAQ92zZp1C5SJvKhnn+z8tcRwbrL+n7RRhFaKI
kENzFtEFDLyd7qL5XBq11SKDJvM77rGd0wyQ6Jy7UnhKnXwnzq2xfUjC9/KWMcxPVeq/PO7I0E/U
L7TpmOcX1+gTi6cP+bYD6uZ/RO1Mx6Q6pa5unbD2RPCUtfSPkIsNVPGzPlJ8BmT2hjPVVt1Uh9rp
FaqX8AA5+CMJ031tuoySqTuYPfeF7bPd+TzcZiR438in1K1daC+akkTs+UPXp20dWB9OYO0RP2IA
uBrf0Zs9dhNHvLolhrowUuns5ejKHRIBpWMx/0+5gA/h9kPh1eBKc5g7ik5dMyg3FtOw3hJZIv5k
Ee/ICvvKwW7/iNWhlAqD3AYBjv4ZsG+xJEy5SbpW4lOKekxrcXOoi6bnRaBEEf8C4JdsMreUUdeU
VnPVB334CRMsSL2ye/en5aI96Z9w60rNq7HTiAjn+tqrfGR8gx8lUo0tfRgzm/1eah539urKD13c
sHcANBeNuxDrmnjzySYKjEnKamUikqVh1Di4nYm1xTClsc3LfZhqzI//f9S2dl2qB56lDS2+kDyv
/AmhD8IYSC3yteBga+OuVg2Kbay3RlxzQKNejeRuwRwbkKoIsL2NbrBRcgG/YKjiCv6Y0yIzDFtT
nmkdeWOkbws96w5kQbaceIveXBu34I6FMHjRGcYvv4DRvFGaiNQDFkelln3dq7+ye7HNjmyTq3+W
cmrCo+Y+JcATJkPpPClB6THHK0Pq9mU1Yijn25Uv286+9MPy+GehASrAZCvoBUaZsB5OeAlemIC+
eOaKWbhfowAQ0MigI4roRo7HyEtq9lkwGFXMPhJ/vqKvCmAhSXtkwyRMnMbeNYFAiUEhSsHg3IBc
yl3Q7DnCnxxaioOdCG4bUg7FmT7WWmh4Ff0a8Rh6B8myYTZcZb/pXFgMgsH9ALCEZeonf/VERGTp
YTtXz4KV7S6eKoAaukO9I9mgWlpBUdVF7DM/g7dIbftl/1MkAfCdLLRKmmJAHScG6frpvHT1ugcj
pTc9V7Z930g94k3V590ZvWAcuaH12oML3X2aTLTKWXSFPoVmz/y8TJ2DV7QySlk1iqXrRy8wDedA
LphOkLWW/RMUSMF4UrI5bzacVVtkCyOK5Q+TbelFWXk6KQH4nNznld/+bpMM1yfp0A/WXhiWQLx4
jVrQOzn26V9pArdePxrSwAEYGUbM4S7sFnRcLPNVIcpjK2pRa6RE1T4J0yzsnNPc+a8Tb925Kh22
GDTs6D0yTn2RRS+CGAdH/hNl97Xzj9/gMzJtUmpXeTPptewzWpLszU8GInz9FL42rx0WFQOShW5e
mTw61/MjmFikvQTd8w38TOlmksz/EQBJxO9kP1jRdOuMbzVcYAw7bVchYlXgElwnFm4K+4A+yuXe
BVEeik6xdjc4PCZsCJ9L4JRSZlYuJjqfo+D0bnikRPisrCdWDeZGXhLaRFpKoHSVnC4/5YGeIZXN
Gch+IY9lGacXn3uZrpElQiUzFpaO5DkGuB6zlUe6y5EI1FP3gG2Pqg9vxDnbHniNDqGvENITF88G
ICQONkH0IZr9R8lrCDakZz8no0cY4kVZi5DU88tXrZCgNjjoRXblp/f6teJds6+l5ekyVW6p1Mwy
4oU17bjoZg2DC21wLjv9HMryHo9EGwxiWOHg4UwV/U4iix8n2m4jBJEaQZyOSX3TKdc6FD68mr+x
q3JQeFc8gH2A3uQiQyCS/RaTAIJSgQlgD8cy9Aw/EvRDtjOOfQC/g8rczHg2LRsX1mj3hDxkvjOI
tf1mfMQdeUqyvcG8UH4nXHjDXCWIz4lQiQB6VQVG4rC+e1j2mjy9ehNxxci5swTaeRKrrouhGxz3
WplaNT+CS/d6OhhghJL/hff8GU02Av2gyCJOqBm24dLZ54TyKJb6Kw58f96/32vgQK8PiJMoiYNT
TcxOksx6E/K6v+cLfHL/Xa14ZN+3Ujx4Xv2WdaHoc7WPuNlLXTQ/sZNA/r39VSqbFT5pk3uktzJv
mPyaLFnoq9/Wt8ribA9rxBMZNobe1yYt9qoLPSuxX5l9fnVnhxHk7Tx86AIMLQ9JR+OSB4/OwlKV
v0I3rq2QQ+m98DuTTaGKbtsHmkzlBwBUHhR7i24Sey4ikokLcGBJvx8f8Zxd/CBV6aaJ/OI2XquK
jjgV8HgkJvoSi9LUPX9nR4x9+Hv9w2pGHBkYLEVrakUyAxTfGWPV1Uy8V4w6k4ykhmowpufEBRJ7
yihD593JI9fxWgVvsBJo+63+BNEZ3weZvtO9a8O+VdzIYSjGQU6juBkp0cqjjFTdeb0Z2q1fmyJ9
nVPSIxRxW5QU3Ls08KVE19W1Olg4CJzx/+PQ+NiT5YnEUQNPZx27hcJh/jk9WrDwqRKXcjutCxYu
neGIPIgSPKQd7cAozYhENat33stII0Gz40ZXgQkGLjstDk8u+/2LwLzoygsLnqyf2iq0w4IL0pUh
7IK29FM7nmpgVSlT6BDdTo6oOHaz5tm3udWPtHha91GQBJTSNgRvgsczKRTrppUx0ADVQgZxl5sc
kq7VqYPZnctieie+3N7JHt5ydTxg2cVGYP8/LFko5gsdVcRLwz8JAHnC0nSZpXEbDKuU2uZFEOw6
oGpHCeI2EJhfRcFxfELCj7muXEAaA3GbeTg7BeSCX5SekdmJQ3cONO04ac0wnTL30GYsi10nayVp
cCJn/WpJ/jZxSbuUAURwarVEv0/QXbTCzMP5I+wxoJgqqjmqyXX33oLgbCCbYr6zjcY9ERYvSio4
tgYuqSIqe47ZVHw6JVG8m46ODB/TBESvqW6gxV2hblvz1vEjVKuhkTFz7rSNw7LTGO5d972hIljU
dV3UA+k+H9BjCAooSDl/PWdFbrqmh3cWQfQ62VXwMJ455iWchpQdRjL/3dwWVKhNXBJKgdLfdKgA
52FSEYSoYjPUsj0q6sTPF+nmLsnx/50bVstFIuKUbI3kuZBw2JICODQvk9f/900FWg+JAXeU7D2S
bGtIofDP6pEZCm1xcv8W4iN+8Barr+foapVUyuc+YiwtXjn4pwwqfRt6eYuegYDSRDHjWOfBIi9v
sHUNGeKMwGttkTPfnlPwF2QAuWYKwNXizjsqLNl59AfoxlLgPyTJ9UgIhXJPR7z33FHqqb0uPqfc
KICK1xbJ+niFV+3zmd3O6uBW8B6DtfnhRE4axLltSDQKcNIJ/BErsqreqIzTBtCncEeJzYi0Tojw
mAgDPMoNbWgtAlNJ8cUiv9jR6LAarm0fCXvNGSJ43I1Qdkt5xSohh5tTKIUPYRFm9lau9x8zkWiY
4/caKBn+6923UA2tHhEiFC6fgnfQMssb45vBwi3rQiLvkXfaov+IblbsD6M6OPttLRgloWtmjJYs
GfW7xdLtdKKtP6V9IcNihoO0bPa/ykP0QvK3vm/OFc0KfrmzvQ7Tx58gspA8XvimmNORoC/Y57Ie
a5POilytBZviufrmHyHj+xiZncUaYF+3NhL1H72mSek4vsYsTAB3xpXMt+NSTBoB3t6l/YGH/2Mp
NsfJZSovYV5AJtsVykUzmaoWg03VeItgynbSabuEKWaJ66aSy9rdzn+6ORxLOd8L3adwewgO9nuQ
3bKU883HLb77wG7OzTAveKsiqKK61ZSqDeEBkyG4yonSaKaxLvnDOvMwUvmOZ42rMrjDAUKGFZAx
NReolywYvKuGkh/MW/keBI+63rFlPnSHIGtT95bxW1360GylmrAnxu2J2VvQKqaVrIm7LhOGsq40
FusaV6xdMlOot1nzeLz6ENsZQck/Rp/LEXx/0MTzCmGJSXRywfsgVieGl684Pb1sIJdLShuI/chc
qyGvRFZ3n/waxOYILU4XcFyITjr+LdqlvcWuTxlWILfYWhufhdZb68ebIri44ZF++798OJM4SlzS
1Jt7plZLdX7RjhO2gGWDMTp5E2MjWG5+fqdfyeU5FkizAVw8gdfc0qB40uv+542B8PKprurQ2A1/
KrBBtoCSykLP4WediRR8kFqYOZ80CcQCNdRdwm5F1NVowSREBoAd79NoK9Tg9EjaLbr71eGCFj1B
oLLNr7bf+1U2mebpEbY+t+BkS/AOBxqmRO/pwCxurFUjOY+5MPJpZ/YBmwykNGNDiwdxstwrBSEd
4eMyA+A77HzughJamsJPHpWlLDQAdM+xkZfOX4vocfPeO8RlAJfDpWKUAWDjpA1DLYpmbQPQ4Wo7
dmzlQwKqh6IaqNJCdTOAtan2WcWEDGGzHBhCDoASZOfMQIkQ7BSeP2T3HoZcIQr7wQ+NJVtuNgp8
mcHD4ipyvjL0QmlHFcUB8gi1P8NavQNOjnyFMqwPBX0AIR9QoRX+w2TraSMXtQhI7Jpv6AngV7TO
CtoCwyt+5oSDwxDbpxNrEZkZ0rVNY4YeXaUWUXn+PZp7Gy+ztEU2SvSqlqMac9JVgw63DlyQ0PMl
umrR+IZR0oXRJVFuwlQynYAPdEGF8b+LLYzYmfgfQk8SL9/MyOwX3U9rAsFgxsgU1Ud9PUFiEYXm
AC9Y8Qjsufsffsh9SIno9/SJNjv6ICHXcahzqfkr1ouLTfABLEY6rpAB3BbOwPAkFo37N4ygJI4z
T0GLtMtOKDJ6+FqfcChCptN99ZoaUrqSs6wkUlU2x3tx1i4q1kgdz0QQtdBQzSAgTEzCvvB3bSr1
stCtgYhOGpU+SSXIzGtr2SfWvXq3ylOq4EdwhmUG1s8gk9x28tKuJATxWZYU3PMGBMT7pwnKeC9s
Xex6/W1UuxoQmdcoZM0tSdPEjqiBnLtIr43dEdoHlhAycr13TqZpDcGB2W25GStx8370+xYPGLg8
uXAPX7mQkQ4gSzL1tZVYbouejh8i+EdJap62aaiDAi/IVRSNZ5450qCpfeGI8LdBvb5tNv5B+zvg
K1yqn14Nsnq7T7RZhICDDzyzGX5fdcwJ6qv0LPjJ0/fgE/N6u6DYmO84qGG+Ragliw76VKO1so3B
1Q7W9+UBDH8pTenNEL240RUUwAkDNfAStJn4muHgcARiKjDZr5VdwskntBS849sJC9wY9HY7iuU6
8cHjyzVVLaf3y+Vs/Jo89VO68rA8NApVWNWWwNKZCJiATSFFjhc2OdPSM3mmoNghX9DbwaPZAW1q
iBkNsg+Kjvz0rMSniHCUbc8v9B7eu6YlWtgXgk/+HZh6hl1GRdvVjT/hGrvUPGu2Z6gDzhMrBuH2
XY0ILBon+/9XIIEsKFM4QT3qutRIGKHhw+3GHlwS8bLrZnfmstLRkq53NRFm9wpCu7mVKj/AK2ql
LTdF3zPyYikxR2+QkaoH4z7iqIPFSkU3plmSWyVuaFf2//WX1DeCfvNhSul7N9wdql1i7gKkFyWX
hCG0A3yAsPpMeHehxwEBY/rB2+EarmKSEs4bDJBFZEk3IIC6z5fxDt/cT5tC8VtWiTJzJF23vGlQ
Zkx28vl+ErOgee9s9uR8U/mSWi9hbkj7k5nSkr+yXmdp+y8XD9b6RLfpLBU8cKdaZpmkS82gMTAG
O7NNvynAcpcWx8ZXiKzI0T3CW9VVlZ2or3oR6M855bvAuiiqR1XIXzVi8mwzINjnICfmCZsDnZEC
FInRSa+B8jbcm7kDKaMZZzA+ES55/xsp1/QHsp2+SW8JUPiDn+VN99zZnTKfqA+JRmcj4Lqh/Znu
X/bnJEo3WAq1OHURu67lH5nSe/X2QpHPuMB38bPmZY+lzrKC5oYfZJ8N/6pOFwfHN3gN27lJApm1
tnGk+VwS59SCndfSbckmYxrXlKuc4IoXIZxqGpVLDWeuBdrvVZCVnteGosL6YZAAkMAvyJOvphg/
BM/HdW63GhnJqNCKO31bWMPmgPO0HzhXlDP1mDP0XUlGI6aEe6GXx5zhpPLoUW1aoieJ3oXskCDt
XrfP8L5aJWcVfT2L+fntnNOo0v+OCm5FS5K0xWFAxZpY1N84CYFjEa8HInBA028R/96EXJ3tuC1U
6+5o2/AZOP6JjB8qNxrHkNyMoFZ0yDiGA0htFPx04O4Mzp/4CrWgY4YQ3nNSgzsDoRxKBqqTcc5u
7SuiPcOSgIOXQhHiLcAKK0IuBF4AlWNQF15KMuI1mtNF/U5votOlqZwEo7MnYOm0SkuuxUiWzjiX
c8sZTnNQAhG0QG2SeCh8JWEyEb1MiuGBCXYA8mDIKMVsh1gQogpo7sKLKfrXxiigoxa2SnJCYsOG
sNGEgxzsADSpK/BkHiMI0ew6eG10VCUt3CW+dpqg+r6dsdPnOUDK1qnF9dR40Ojhycb8g4oke+mN
uATJQrZkGoZWSUWC/QM4RvvAjsdp4zJosFIa1Ga3H31vo8edvpUjDXLPy6t4dWoXVpc2o0/2UsYw
GKruwdycuXsW4ZsOm8zFweha5GmkGXeEA6AJzTSGRTuuDoXxKXJYACELHQz7jfk24mBcJHtIS0eq
xifOGb6Iju4jB1eSf2Im4MrttTOz5EbD/EvO179Hxpbm7x9MmEI7USeV1iJMfcnsfUOCCVAp8Dxc
Deh27GSY0EidNYPbhrfDusGKZeQBNYoPtnAa8ghW78e/ckP8ENQUoTS3mFWkUDHPzLCojIqYhc12
lh7R3bu7yApsvIRB3qa8GfkjhwsTrCFvO4ZCEDJlmGuFw1uL4vj7+CUf+NBC5UIse9UI+IfoTOO8
trBr11b7wjMEXGf89UpBat8Cr0JhxK0htfb5Co8qqzYpLHGSo/waDErasNKOjXGFnXT/Gd8KEcG4
BOSLxQYqNESgIfX9vEMEyXPQXTPbRB9uA9edd6yuUAIwxoQugBYaSdztuXDV/ywmwF2Puqg4GV/S
575/MjdMJOQ9NPfY72aQJLTW5D+rjr5s5Y0N/qmZyAUNTm/5Ugik0j2gPE7xZKzV0Gf/sZC8at0p
R3m0hbdevVBCQMsa8VOQ2us80TfwM731pY3QOKC3nA3EWkaera/ZBvBYE0I2BQm8nAX7s5Jc5aTu
o0NuuY+OdXrfnoF4wKAOvq5IBlyTLYW0XuQxs922nHaj/CEXLS9lg6Ot8r7DkMAQ/D9BS+HMqTuH
lldDf0LEaA/f6HkqkPg4VdVF2itlqoDXqor+D6eGo2t3g6LOuVqtqlA0F23UQfsYO2f/zHNOnXOb
vCQgbhFfB+uXt8P2KggFH3LK1ebbH9HogPTXmVONzHjXr9i+ZRj8zS6Hvzg9Rt0E1aGuX09TFfc2
GjjYWLjHOBWfAEv/aLrgQj60zPiPznOoHBe0W4NMbtpzSqJ7n3MgKxRd13XpaCK2Oles4S+zV8Wc
iJrNsYuBfFMBmiNuXI9c7LTLZb7H0Xi31grKsat7+9/beunpXyJKVH/Hjbuq74RWbFTwk0fuen9h
B/Eihj3N2tIKtHA4b1XrxyDlPp7WdJ0JX4kzN44rR3swn0R29EPQO/VCbJzrJHG2gVcpU0aCPpA1
KXXkJMM+Ye0gV/jabGSTTNAwy+XKxvwYXq9kCJcG6qt3DHNo4w45/Pu8ItZqPc68WOwkTcxu3BB1
8+6+xSD8rd6mK2exowLG7/WyDisU5986urhgBS3vap3bDLixPnJzmFDbqzhmanJv5TH49XMwhYS3
2yfgb3vOwWqLwfOKNaALX9x4Ngyfr1Q7beNG5dImSKqv+bN/2LsBnQ5sTKFLypOl3n1dwzWeR5KV
bqSXS8GU4TifISRYq3zzT+0tgoi1/oKsA770OOOeeQEohsNTd0jd3dGFbhCsf3updlIemWtmxP31
FVZ7aY7CZBJWwTuf/tDTucp3AZvOL08X/R2EkZG+BbxAj65uv+e9P3sdzk+L3IOZ0SQSuGldIQIG
rnv280blno0xBWbMSPHn2FDWpowy8eiYJqlAIbxzb/ru9cGnsuOJgqAVDXHm/zivDKEY7gd2SGI2
VWRCO86RNdAEOQENW7e1/Sq90lfmvk29BbwHBUgP+kAszOeItGYBS5ZWanyx3t5mnuSo9eW5un3G
Ct9AsyO+kvUvdhyGj/3eQ74NzVYGSDhHi01rxhGFmPgg5Lh75uk9bfU5HpekXTQ9BW4oS2A1xzAA
75wDNW7LJBFInWDqeHtxOI6ramrwxaokMp7NmRzlprc8Yy5bII0XTiletnFexxTC45/f26kNoBAX
FYaR2Xnps4zRNjq7QUFA0rfiISA7KQaZQ+bdKpg6Vp6c/FNiZgLvWnjmWpwzprk0srxAt+o8R/YL
SEREDUFELdeZh0zLM7+1ZI/XBmxVjKDCA7Q+un8PF4OpNyNXwOe+ZVvwrUQHqUYqtnxArALQ76s+
EnQyTMfda5XasONRAGF6iUxnMJpt2p00foXluU8jAcGrj27lWdPxAAOn1sGOyIxvZlovaSexi8EN
QckBoaAmAf8kvUWCQF8JL3QS/20JiWWGTsUU+Xw78DHd8JML36czL6zJ18CEt5bRZzbh4pA5bVra
NMU+xGb1H+8M0vcFB8wLYsS5QGHXDTS2/jA/rRszJrrZ0YtWGXTcFPVkVQ2h8H8cWcw0frGO9InV
CxDfucE8apaZdeT5JQ5PhFf4LURODNAzrkqDHrpN3IkZ/tgqkiwoyMhzYnDxiyuyxf1xNyMYaHog
u3wdBrLasxTKkXqBEyAlIEaa3jVBpC1VRtxXwYWkZjeCxt1DJ95SyAqwk46nNU9RhGWi0m4+0DVd
89bCehSWdEXIYY8rVFaRDkTyee8BN+ei2wAPAktld0aUEqheuqiKTIdVWg8/DZh1zUWzqjzwDc+9
D6PLfzpamQV7u7dfcU4e2RqeJwLu/yRcqWiuw1r2pUbdalqi3nxpVLgVgcTQKFmFKAHesyRBLskd
BATzExQxGxxjPHIG/iR9eS2hrMGMviVxsgU4KSWuD+j9UJ0xe2LHcRCD0Ld5G92Eb2TkW/o/pR9i
1T2ueReMuZI/tqd2gKupvJIcEhZNLX89jj5gZVPsPXKKB8PQ79xlVmlpHmsdz8uk/TMjvmyhzTN7
OmXHtQCOCg91+hj+uE7ean4MIX5lEU5K78KjZ3cgxwYjjYyX39wfreVZX8baiC/vKm+mBsdi1eUg
u9MIcMy8LJCakXIBv0+kOt/ISlMT0Z2myY83izrWqtaoyqV6dE00Gb7iU6yTb2TJxKWSgQ3tDMxP
5YoCAQAmhvEHKcQIuOxNsoBQDWRdhiZm52ZdslPlz/3QDbUlSauIaWpMFaTckUccICRnLVWmX1Sx
S5GTVch4TyDJ74kXLebIgoUzfWmNLj/7AuD30BU9LDzJrYmU0jjFOEK7D53HeidjWl2tvJKou47s
LewNS0ZNAIo4/6E3ha/j5PxHe2cc9k1/AMT6Jl5qIEVrxrOiNo4nrrKPoaBQxGtIv25FEiUQ/kQ9
RZLrkVYy+sRTKMHCBtRo5T5g0bn7GjFJWwC793BpCtm12Y/nFAa1QHmX7q7hfGJe/DFcBYmnWMTS
loQyHer/xTs2AIuVyHuCfxHAO3rQ02/68BMu5GOotaXg67/i35fNsM/wYm40i+6FdDzy+FbwJFo1
Y2qBV6X0+EPmEB970/OFhbqDzFWmgPMxYNj4PFrqSU6b5SFd3ae8euuencwBIR5atRYOLBZG5k+M
7s2vW3uiE7AKo63dlxhTZArgTvdT8OnKQFU9fzKeZT7gqk5K8Lk+h46LRQu0Ab+9DadhJirPOAGW
W76C932nUycvKV1RQAoaBdnPVffGhSanTOuCs+sJqyRIoNWxaOFs/FnKGMnUMp4iodZz23wtNzcO
3J0Vk8ZN8PzoH2SDgF+PXi1zqDtsDGDRPE/THx5RvrNS3N07AIMR5I1gHQRYB1R+72cBnh9Tq/Gc
P6gLriqaTBvf/i1kDWKOQqz20b8mi1+uRqsRlWe3+E8IwPWBreNqfMB2zi2WEZ3S6RuPBCnT/wRu
jAfn2xNVLLjCF5sk93y5ipXeaAhT7zRbvh3hQej4J2Ul1OdC8nzN3mAGNydFz9fw5x+lnwWwaF+9
1Kz+cRqm4xvD39r2CC3Q3s74qAm9JF19+YNNFXjoUIpfOfCMsWbQr6uR2UgRhAMwNfQDUJzUpinP
94xSQGSnh2cP14OQPS8cTLSpe7h5vBZZVqfW7IHyNPGZqC8ey6P02q31DljTaQHwXEyGXhap1KE5
VdgtDwacKMGRQoOEuRvKyRN9bsRrwysf9zKg2iZoogfjEFBr9Iry6ybihBlQnJqkf2+c3U+g1YG/
jEZkYAB4LtVEnK0vuTz9bc69njAZgGu2hXeDaZRv4eMsd7i+lIK3urXo1ENZTk/yW0D68e2rkisa
5DyNK6QjU9kOesXpeipmSkAK9SVaiIQtD9/gp9/kgwU3g1RawlGD0jD1dLM3hv0GqIoeMt9Q1Mp9
+rrijSvSa8IYTanq5pYfiJWCuvSTqI4XfrXBlix/kBHzx7heBDMuzUZ6Nbh1RQx+uGFp9Ah4obEq
+n1qDn0fa0pIy6QFFQgenbrFv0X14PLxxuCQxfBdgiDfs4ozgtIYsCRdkkAeWLw0+NeNl4vn5bYt
ubBa9Jor6SfqT+rNT9GsieHYl8YQ47Legk3rLMgAGcuVdzsj4bKzkG/af7c1u+Ce/jOCVW20gADN
ySjwuDucCGxg/XNbnTtPMmyzbnrhcS2oZbmW46BpJq+KLqu8rR76w0xJq2lAevERiJibzUXbBhKI
vOeFrAGiWCL6xdB6fOLspv6VJ9i/AMRtPzuu3Lqzew0qsvDR09MyzRTP9UCUW8f9o0lYKw72Kxlu
eHLkALdILrFFo+RQusAxVMhLrPUn6mwNiZzhDTb/VO7RGsonzlJzrcv9s4cBSWFhxGrRsVoBH8GY
38WxqWCqPewbiOb9roDjTAfPYFufKmwoCAVyB/rwch5tuquzAb97iZo7FDNby+9d3Qdea9xpt1DD
OuLNcd9B6ZnDXnZLoLyPDTnV26R1FsUoBwjJGPsRiPEkSc+F2Cfn3Ig79WvdMgyt93DwMb9lFSeb
5x+y+SWc1TAQFqfbmCSrHAqL8RKN598sgsWMUyTOqhQZsHg6Crk6XnbjpYix4ZaAqZlOnr69U+ap
SWuM9DaJfVkn52ra7rKxPuN220bmq3CFQjzF4oubgh5msFw81z16v/Ug7yKRUdfnL+S4DALhkVi8
4z9r/BWf0YBrnbq4S0R7zTob6y0DtubYxdWXcfa6B14nWPae81SK8ECJCPndIfGTpU9zEkvgYLZ8
DvBNgmX/6c3AFhJQmJf8+ddUqfCuu/ZU48wmNBn5+99O4MXf457xHc/bHc8h9Ckxz+VorQ5RfVMg
iH/zdo9iwniFQuSkBgmROpj+U+YxA3SnTeCPiHgU8Gv349O7v8f/miJRzrPs8I/tGowDCtH5Hsxm
7NpKDJy4CO9xXJsBotXT2W/tDpRBT8nsQsmccTMvIDIZ9WjoVZgd5q0gXF1/wgt7kxUa5OMUJ0lq
2wOQIr8VdNVztpedykUN5utlzDjJXjkkgD4Id6jVgxXYWK58m+z54ERISQI0uNw4fA42qRMWnLhZ
H6bWxMkCdW5V6Z3qI6ezXRIGKkWQiZvP0MJJxNRRYkbIRjbdOsmLLo8MeqAlkEEWOl5XWQqI1KY5
rAOqWB8qEuvBSLcAXBap+lhBz8z81f4CBRHavg3mbUeC7obMDt8R52SkFYyhmvqvxSuc5pXtdMvt
xfCcv7055sATnuD8sBF4NLt/NxefAqjrSd1EHr9cGOoztkaVMTZb52Ebk5dPuF2INbcFvfNPSmpv
qeorK3dJ8h0Y6xKnZoAuFfQFMMAuxcuCq8+qXEEBnYQBK6+aRVmFJJLzjVm5Daj37njZWMdUt+Gu
b8HQQl9qpAHS6jrHuagbN5255ApMlgbt6cuFf+Zrtnp1/dMNNRD3XjsOsB+tycE3xRVg+b4jbf2z
5V1yD64AQZQQY8YWWo3/LPY1DPm3DAPyqz6BrI4LrixlDo/y3KmoPO4N/aPOMHS9XLdqykSs+kCj
9QhTNespW//JT/TpPwWVzAGxzqEmGGThVKe2vPnMSVFmXt3glgVUVF5zGJGtBw3gJPUmbiEZRnCl
3kGLfQnn2fb78nsnnATHuzcFxBpEPK6AL91KyjgDICv6+i/kWgz+nd6DsTnMvEa/iUft2Aj+lBMo
Roz+KdPw8T3fsb4Q6tDB9lVtOJfiPQksHvt42QoD3mnNMlu8WRuwVq7/d8iwm3mLUjZsTUBJTuJG
6WHdol0CmAhfrQcxeMfCnmTH13kIydg+SQtImwZKBlFribVDUX/EfIY1T2PPO3t+gcyZymoVqulG
jcMdl1/bHiiZOsoBf7huMdS5E48rTR9pePyHW/rUann+U3oooDfsV9eCMlaoLsztlp59c5nV9acl
TOhnXg3UiifzJ8Uyo7IDS0c8FADdJvSNff3ThmFi7Rq4mImI+fzzPaZLhEasy0y5RpH45vtBl6Lg
eAVJdYzYn/Khv/zXyF4awWK1CzpV2GrAWEX7HXrXM10GGlDcK7HKbW2a5CNj5t4M6DG5yh1Um4wx
7K4fH5dWw7rNKMQjW9hk3X4DLS85XJmQAtnnmx82FRceQRvlmG8J76cT4C4NwOjafu2C9ZFXRU+p
I4TK5QPv0Tjfo8oN9sAKPmvncmHwp0mxKmOZULJRRXZhdGQM878moifKjrzcAQm72Q3vyC2MPYWu
h+59D2vQXP5lJKw9o8p3tXqgqIqUPRbWJq1ai3NjH6vT2oD/KJZ/FjbPnous7cRya1SW9laiJ0hP
h/M89tBXzsGWII0al62JSI0xVI56kkYQdkhM8OHFIeRwaJHKM2b2vS6QZv1QO0kv+11zoAQzuvCn
u5hAvVZ9/2zGybhi8AsbZiypo2wqsBn5UBRYT48Pi/ARVvoWoJxiJJK9nsuENvG4vv5JyQ53sqto
BQxFO+BBus84pCneMCbalfz6VXl3NgwoSxPHuFdfg7YIzkVwIm+ydmd3RNgL8HtcLbbHEanNFl1s
zEsMbEmMSplZ/8aaUS0SaEjYPVZmY83gpXFkgYtQsKNpc8T+7T4ukSFbibnkPen71McDSwVaAKN5
Czx0o2DY6vmoBb2QSUX2AFwXc6kHh5pi7YrkXIAvBV2UqaC63cWtwtioA0G+igV5JL2Mb5fAgmmT
L2wFo4ruMVZCVqGg6rZHZRTI0QrbzjdMyP1pgr2TeyxYojH/leUXMTaoYHMKhBPPeSbeW7E/u2/j
ZLE0G2L5vopOz53XPDMOb1oyf0JbZSPcxcVSEXTyBbqvi8BFLpxTJ4dyTCCHLQeNaX7J1fK5oa/V
naW9/iWbgEwdmdSffASVkJtiHIeEXXsAtw5Mihp0JnAoKAgCInvSybNuKVfXpfEP8e1xjboHqYDK
bi+UG2fLtcBCSk+q/itokQrD+iqSzwF3Y0usi5UOyizBdbo2dFdAIauOhEGW4GRtAgx89dVZFZD3
2YUiK/lruV7YwaUKK7ZbjoKx65ppJrglRkKzXRjqQpA4tv93kmnRN2wYnFD7cPMrTj2kGUVkGyEQ
0v5rrpn8fhgWGXrmG2Fau13fh0833DSIAHUQt2JNrGz8jr0kK/g7RI1dwPDHa2ekQl8alzXnNV0c
75xbOl7c+jujcDyzBCjo054BXj3hYvc1MJVcKDWSjX4ry3wXRb3fGWqv3O1CT1mpsdWsE0dhE1oo
WsHAuh5R3nYEmLI9bEzWOpX6d0Jz41h3E9UDWKtCiQCzwXmlCVCObR2Xl9kInq0Y+kLWGxuDXg39
Boti+F5N1PYvVW07Vdpcn0g2SaJAq5QB6vLv5md0qZBfffFIgZGddmf6OPEtiZ+LnSFpiyQpS50G
xlZP90qqdl9i3Xuns6X8gQRCFNcrLK3N3KW3BIJuvDWnQTeSypYd5KpbJv8oOFLiE5HRlVtSfPF5
yp7l4pmUBAdQ+RK3wVOzO7JIQ+VoBJJ67Rp41TUyKHX/A0hAw3vsAVfo6HvYyWzjU37nGAuSxr5Z
5R95n/u92WpcF2n+woHOmn4IMCj7pPgj/7/ptfnHj+r75gOnDAJ6I4ADyVGAEMaVGEfTeE3Y2nFC
JklfGQ2VK0eK9MbIOKJ/EL2znMOVirkOPnZHDVl56hKXJIrDe8muQUGzETbCX5T/lA8+QydnGrus
tHS+oV/Tm8NgV9REc5n/jwUHXCup6cv8vtd4OkgK90TJPxeaFhp0We4pB+1Ed2OyDVezphx8yLJO
AT+aHrQygVmTb8BKJPDAxYaba0yOBSWO4mLLLSUp65K3HzCXLTLoTdRer26oSBLd+ObV6mKth9dT
bVxyH2H59hIh8DrX+1qJbHM2qNn0DCFzzeaVJL+tKK2AcyUJydmzTZjJBGlW855o7jvrTSzYntbN
/AUDp/t4LRI67FtSbuny1q1rpP6HAqloKqOkNJXyzeEVviMapNCD3B2KUBq2JngsgsOMSpaFzJGm
yx/FpePzMnLact0+ip9huUAl92MexhZPDZgJw+LDUqN48gmpPiim3MdnebdmwbuqfLWI3smaCgD9
8RdSTVgCRxfjr6pg5vYZZTMh5xqcJy06bViQ05GdRaaVCorub9dMqDpqnJ8Ne0gMBsuVQnYFPO0c
E9ucbxRgOS2uwKs2cZqI0nAhpegJNDkmYtrfZWOqXpJ/LNnJ56vAi9XyzZcBprfJVf9qt5FqIA5X
4VXDk+CWqgjubLJwskjBYfpVg7U4bPu/3Cl/aCja3lx3lrO6Aool7YDYBbKNUzgY2D6QSa7dUPDR
8PebDLdt1z3bz+c9hzTe/2BN74o1rFhLTFUqdMs3rJQ6oDPpQQqXF//PYgNu+0FzA9kXm2+thL8P
anRR4ReW5jZvjrAJCmVdAKsg/I3sbAPbmkZJ4WdyOtpUteVyb/CKQptIk/ZiUw3bhVkNZHPKePb9
Bks4YITcRbwATHxgWxghMzIhwdr/N97p6B1y3dRJ9ZdOdXyEWjrOWHH5ZMZa/3rhtf7n6XKhNIoj
WJRSK53MeijLWQzDliwVyWHI19EkakSak8UeJVcJFZiywcD82RgEnvlss1Ex0WbWCb37OohRELKe
dO6j1Jjzs2kTzWal2yFQFwy3n3wyXu2xWE+n7DIOYulamcMak0JjUVeSNEd78aSH0X5CKD+4cp35
m8ST2QBYjxHSq2LRqNBjnY0EWIhkNr9Zx65KzWaDqFLBoy2vMcBZMT+SBr3ElQ5wCWwVTyVQRvTS
awlBn8RLWYNx08wrc+/mvj1PvK0FJvlyJKpY6jXBr65EBtt9MrUoD6q2PBMXW1fLXh0jUV1BxxSY
zZaBy6+2swB0UBUHy5GSc+FfypW1sjMl/hMyh793d/7xFu/D7MOHCbTIfDws5GsoqzGylYgWA7al
xul45t/nb1nQF805fyyCRZgzi44JxyxxINKLW4lz7KvfLKaoROxIz98dMheVsYVqpJEpB5TiLEDQ
G5R+GNM50Cj2qN/DTHinf/0cFfkg1MPv4ZjwMxTzRZUkDE8EfbBldUIUQ5tyf9RuqUG9e080Gqna
sI/v0hUhFh/Tj9Pj3jZwx+fjPTRcd9KFfFnebmrveDMfyFyO04i1oNt+RonAENR3jUi3lXyPE9k9
5xK4t0ViXOLrLK+7nmexu/GeFqZrkeSfjrHlNu2HZe2XgM9hMOy3rMbhuaIpkOWuFBIlnjJNPc7c
3j6J5QVuttGjhuL6NBiFziNy7urUC85AeLlIEqljgTMP7Wo7BlqIWsuXph114d18/C3tGiqU7Nj8
FjxSM49wGEmGdK0qHTVxKl5e4RelK6CQ2pl+q4VEE2P4Xn8S5dGWQHLpo64/LomypjLHTo+F6Gl4
gzAStHrR/uXL5f3iTdSw7fv96rQOQ5rKeJXHRSRQxgGBqZcG5wie0AOBtGVVTfmdAm2xOHmUqVk8
0WR0jJgim+R2xv230BE3979vcUbmW489mXjopdOjpuAprrwrVU1oNY1SPlo3mhk4485AUsMVWF4w
v2ZO6VPz22aZaIS+yMxqgalhCnPEkztCXttIR2qnZzzjZ985uMJXKU9sFtqc1R+VdzCPvBQ8IGxw
BSgMitOrbg6X8zt5ZIeOBJKl8pIo+2X8vkul4MOVpKPP9d5rUmK6afs5wrfHOnAYbg8rQfBMIpMU
+N+5Ua4WX1MRpUyCxGvP8yH87geDsi1z+4jYdT3cn7VKgRcHVvn79669op/FcZy8xzQD/kZQx42z
0OISMmdL71iWCl7XxzL4fOPMv7Y/OyfR1ORoSSEWPMsYlghNgJXX3LLUCuEJQOxVdhNCpbpLTyl1
wx8i+aU8OpemkUaT2tGIM2pn11NU1A8fayx68H9IKQK6VaCanh9jgfdiq5x3lewQbOta+lsKIvRP
KCVvwPSwrp2fj31Ai1tiZjG2HzFDj4DvE2M6zHBlSD1T9HKTlhsUT+2tp4qL4Cw7nCume2ovj1Rd
mN5nbB2tm/bIadQMgu078Z60SNql/jqAgt2dDqERDLlGQHsDIRtAk14sELyreJHTuU+Yjt9VHJCi
sMHwR/EWhc4c22eih7occW437+tZXHU2TmGR4seWUyLzQkFBsk1dtQs4+S5iderarN+mPLqptv2G
MqPayW0TzOJTudDwY0iWLW5wQBNYEWnWfC4nXJOZ/lgIt6pOdRpjajisZvEpa5nuPuW3Zah7307U
oYup5Jlx/3bu7+dlGT5d0TZs2XHT3gWDeMNakzwnnK2J+Yu/5b25EeKuu/KBkrrQl1HM5R1nni51
lnk06i8ol24mHosNUvfUVGwoVcBRK8gsodHBAKt1nWF6Q/NKhlgPyCm2x1rGCjdS27pOPTPYdlwh
NGqQH/tIvZLzEnRcAm2XA2I8ZBn+YJLHaQX0hhx+jHCNAnDnKtBr1PxxIGzkfWvGYO+C5to8BVi/
dWUq+NPgFShNvRlU5BOtD9zq3DL5X7x7pumTwYAO9pvY4++E1ZnMKBE3sTjbu4/hzfSDediRKp5K
8x8ct4fsO5ebx3EKKDml3pZJj9u3XF2z0RgcXCmirtObMbh3JH0g/1Iu4W6EtF0nxvf6jh2bfkHX
N8xxvGk0CQZPy8PQauF1oT93jt6n756gsbXz0T/ggc+AOIdzkbb+CKtVes4VrszMfmgeP88PMfXL
4O8tSw9qjPO0YZueFfFaz//YKtc/n6dJoMSBI0LtvTxCm57dHtbdAtRz6oSWZfBYFcr0X8ioGAUh
tsKQqJguki5wHOTxwHxFMyRatLIvaily+JtqAEsYrhMOqvbjeLauAcaBPnKxDZHrT9G+vCjgVZGi
tabW5+4K1B/L9aRJMgSIn+LOzkposufrdAKWbal1G8CnXL7M8NaxsgW6NyegY9oA2NYjEOQXonhI
tX1+w5iYVyZSeLa15XWqPdjh/gGwMmAhvjbe7zpCym/o87w5dcIpHcLeumY1mgHDD02Inr2Mb4Dp
U3SfkBP6KkTsT18Cl2FPFGEI+UWg/HgIZb7gMJkgiRRp2s3WricjI8GEe3FtRI6dh2Nqtlv0P6oC
rS9P1t/0Ab2BcdHf5D9PJQ6VhZodsMo+T/LO8h+lITSW54wYo8sgy0palmKkKE20DjqiA+FR5oVn
gkKrCYI5aQxqwKT/W+yqUgwV4wfbpzdq4Qntsr2kWjD3k4agpxkUGf96Pyxmga/iWZcCTwDPWczy
kQhSHP0+zlhf2+vFCgKOuIaebhca/0iJDwDQiyvNIIbo2krGQIpEVpZZFCA8+McdLrPmH1yRWiG8
OH1bsufIoiug1Cb+AGQN5z4hN2L1RxlYZ0X5RY2cKqYWPvIyhBrcp2SbJSSIvULkOlgyVX/5Ac+h
K87+Rw/4p+u2fHkDZfUgGZmmhfKBTVFf5yR6uvNWbQo9iz9bqWOMvN4rbFEQ42/JkvaIIjv6q8kr
glp63Q4FkUZi+c2JAdyU7tMxwL1IT7k6gFcPW+BY6bhIm5whB3ZzORoi/tI4NxjrspY6byiUytcj
FyT4GVCTl6MGMBYt/NnkNLtCWOXESpQehwieLfwok4goe+n2UPcfCbllheAMiTACmHrkXcQn6hDP
MLdRMx0+/+ExxOYP0gjQpiw286cgT4O8nxV3Re7KrSblCej8zewlS7A48b0qh3ev6C9FGKqINNVz
B51+AbTEzqKUdcxuw30uCR2dxNyJG3lrl1JjYM9uLPLOuQHGt3OOm56yVtYKDFxlsbjeFP4wG8G+
bEcYUs/AAJEfeq5DVsfy17dJm+gm0xgBdCgANvq9T2RiHNAypEvSdblMak7yjp4Rhpf4gSn/42lT
ymU6fX3CRp/2gyCtXicURK8vPrfkb5fL5gC9ymdNK4SaM90uJmaqwJtJNBNGC25q226YaT8Y9ljR
c+efUKa6s5hQQ4PH7+XOUIE3FdYBJ4uVqjBe/pN9YW0GnCOY7ACd/78LSQnKe9P5jqsA27lh74Uk
Aklo/j6jsAqOu4yy6wY+fBNzwgodHtnc2VNoCHQp3qwfeYc56khmyIj/58yF8BnvC+VIMtElm8RK
+709oXskxJxDaURBatEREE2IUWham63Rc/rsqOZz+y0Ie8ptiqRdJtcGP9sn49Iof17TWu3m7U68
ej6ngKkZYZ1EFWrUJiKmzfsrE2iLjJYx+F152V+nw4qRhEsEKGDltfT3LmUws5Z2RnMZz4DbiKo/
qAVWLEnb1VqQvoPvd1QEg9s3Z66vqY61mO8BTYpmxMurogW0BkY1gL4kGW4Xxa1Ej16MkP/4/7DX
/XpvtNZsN4F1J8ysGJaR9bxplkPDTXGy1yfZLOuzb7RvQ/V+Hxo89FO6ynprUj/RM51BcC7p73+T
/6lR//ql9bUT3lukElgem/MUAf1rQ56YmvEdjwhq4Taql7cRy6zQzScsDpGG+ws9mPTu/RfUPNUc
ak/4L0VrmueNZG5ZoAVvJYrgzJUjFfWYFHwX2Alak6uh4hPLeFM1eAuT//EVDaJLiHiBi8z+D3RC
k0pULMMydqolkRUUOBCqTT1xq5WOoh7RMfY1F0KyAVHNabSagtEUiK/Y+4CVKcQ7xJAotE0k++0m
JdwsdYQpPoO+YvFNXCsvj2+IcZ4KVFSxfknamSZ6bMizQ/NKoCu3fqCry+xQvgtvcB9XoYqvthMl
m7XUeK9fCobg8/4pe+Wig8ykQAscLt9VX0AxVClua/QKCVh9Rxd3McbXly+/xesfVkEF7jsIOuhA
LeJE8BXUVflmd9x0aQpj0DKza3VMtzmxBjKfOz4Z2UucxiLu1t3g4gGlwfUCosyxSuPjxgqk7dAJ
Yep14J1NGzYhY8cwTpk0GbXVjlZxn2thjJA+QVNFpyv9ypAQv74+m54EwO0gG0HPj4907wcjdZXc
7bjT6tDbD1eBPWUb0IIIppkTr2UUPRUr/F8JEtnVn9JDQzTkIqJkuxDFIDnrPGZVFIhXyVuiR1iu
67vRFKnMmsl4k24TmH8uU5cIWKmwMqD6MHa9tlvdhUctvP1GFouaUio4RYprH/MuhFUvBfRNGdfk
H5zdS75k9dmcjhcLURfA82EYkWgYPvHnzyhQCoYfq7Cs7kOmYubQsiClwSj4m7NRyAwgBBuLlWIm
m4a5aOVqknbQU20S/xP82LyxmB4MVAhW0f+MAlUM156qMI7KG6yy+LQao62bTemIZ6eo+z2hyeYa
yHT63r+tu1J4Kn9zynB/eAA+Qs9R912lZrjLNP2S7eq0ejj6bUqx2DpiwCp28q4d1S1g4TfVkcYQ
e5VRqMTxCwaDwJXzw+ys0U9bzY7Ld3jnSvdYdV+lduvUfxQs3PlJZ72FvmXjJEgXW4aZTp3u12GU
Dy4gbDsxlsfH3Qv4TZpVsPaqnFGh0vRjfh39EVnFYqg+VZ+kcwaTHE6KCVF6sXKl2Ppel3ZFfX2H
Y+E1nIS+n0Mi/A5bKgonP2myp9Knf4CkkNDQjrQjH1BShh1jBpowlYI0jtYPZpv+jyGnGjPH3hnL
dTryda8AyV/2F351ja9NOp+kd4akkm98WerUlYwj/tjRvAS7J6SbA6AWhZw5YwDV9jKqb6DITQCC
rD85VTsjvQYR/xExMS1A76uvAcFhEYK2kgJJ4T5LTvWyTkUpKJOzBk6n/ggu55zHxFf1BBcmYh/h
C4mm2/TOtwA4ad5ferHJpeyF8shmAOPAZ1dtLVQDjMItQ9FQhURN3PZT3ZJ0RJKHa3Y859Ijruww
sjhzHhrCAhdG0mz8HSGVihgdM6kJZi3KavhT+4GGwTDbO9YnpCJxSa1beqYuTot3lPpzwCwgAqr5
b6Ptbd7cvhfZDOopK0K/Mi+rlR/H0eIpFLzmdKNhZHmzuBiTtd3O4A61/RSh32G5JSUlndrRSsiM
RAb+B8iRzDcTHmJnhu4Z7SIxipw5LjAWnWQwHeLcGyi5uvTYjDJQTlTQT0fT7ZaE9OIwX/AIcQHi
RpcNQYb31Mcnv5BLXQAauuhEtbJvh15SieyeqdDkIlCqRYBYQZEH3cb+rTojL1BL7tB+ChtnfbWz
DtLmiicpfED/T2hD+T7vmDIwMpJjUe2otieY+AI+/MPTIL4rWdG8eZ/bDZ130refq9Y4eNJ4vtqx
7lyhEHMBrNgmuBZ+SshqvnLAX10j1obVaDGgS2/O5hMxpUasmwEjs4uW1UwhUFGn857gZTirAYQk
axdjrgltWwvnnOtkZI5+4r2YmJewOKWujSmjWP0DNdSfvaQaVvQ+yHr/h97uYSppqE+1kw48Pegn
UgoJ8kMzKNvyCXdGx1Ddvoa7lJithxfpP2ckN06hQK7CGBl8G9kSjFWcgCZ6YRCxkdOQFI6oK61Z
VYZCK0NwrVhZCKEzHaICKbXvsM4JVQ20USBsfeXfqpIMJSMV27W55u8funDa22Y9sI/uqguUPJfD
zu10j52pEG1yUaRULFDY6QomtR0HTCBQtmcyd921DbM5LQzXRf0u77O9580sD0+yDU1Bg30m+bHf
qULNVxrXqszDsXhtoX+w/EVXKaJe1PwE7/RxdSA3vZyY04TC/j50roZlHVPeYmD5uu5Y6PtWMwSy
IK48FlV5gfS699ONzBDP4AuKpHUZtaqesAdKzsMXAnT4onPGZqPHZmgsbEjrUDUltTHrrEnptR5W
rNDfDpat64jlU7HjC3q3AZqYZsGivUs4afLGYFv7K1oMncuOZv7VQhkeHWXJHWzpQlsEyji/UZQi
NgRSP2UVF5RP9g3zxiQw/VH1tZX5h2qtULXwNgf2zIWYLbSg43e5WQW6r8SLYa1FmEnJCC3Qmye6
oxRkiSiJFoB4vNHmdTarr1wlkMw/zC9KDmizS2kVey0igRpZLGhE+t3glzON2OsPEXPN8txRnRt+
+zQWNDsoqcp9JHac4ZnySUWknLcDkFGB0oQdGKhaMpahI9WlQKfX1C4rgk7yjWzShzLVjXnoLP//
EfSCZagBT/2zD/wtOwuKst8VuVdoE/vfWwdkHvMg2FjusuUraAcjBoVqvcRCObJCN6XwcO4xXqiT
1sxy6zE0T/KkkZktFMjB18cqeB4K/zSliUbkBShVY59ZvK/8ZmAc9OFumk1cDM/rpKYPssBhryHj
sGHKlb7oWpc9d5TQmIVTuwAajX4fIxlu1TC61nIEidu5d8itF4QkHbhB6HFD9q87TyIeQI7Tp0r1
6ZlOi3qCENvLHbofwCvnOoJippoTqBHIhi+DS20sOXdcD1Sm0n3TgcjBnD60gywfcbB9lVS4DqXx
2SUX8sI6V18wHx5VQbWTx7OszbLVRgK6CZIWDwG1VPHFJH5O+jcy3QxPqWCIIQzm+kSLt2bdntAP
qn6l+N7ynJI8Zpa2NdTp5i/uJab2ySWXdaD7J0lDcAV7YnSv5Q7arGseRIWYdUwV+tKNLtJ2QnMF
j+wIoPOxvtvwbcbxF5QV5MB3xR/9z8mMB1FdY4M68excHYx252suC2Gi9Wy1xXdcxavYZsrWP7/K
n54lvfJyTTPOzdEC9nDDxo4UXmgl0tnOA1oeV3Kn1iq7403QiEz9AevwnfluOXY8xkoTEqlix5r6
68xFhrh3xn50+a/MB+sUZmG9aHinZfSdEq5HF7E2jaeXwLtxrN7kt1TDb018WyD2LeUSnt3dlHtN
C1HtPati8/HjyrwptBZ/JnyK8KKwMHOyNtd8HX9GcrzPSAthiqi4sIpkkS+P5Qzm2Z8HaLs9Ta6I
0oP2DWfmEr6aY5LRzbsUUAzt32xeh1KGu10PBn/pPmHw73Jco63hYQQytIC1NNsHFb8+oQu2q+VM
y//txVn9ePt0wZTOtOyD7lHqMpEHGXw9z34WPQgPA6ycxHKKDmB0kXJcfjgexCl6+GpdCch3Onjh
Zg1f0zoGRu6aImckYUnP9L5nsqaDXjWO+coswbjX4R6nBMCrBQN5zBR7gh3DjIlcDXF+q1ZrTcRA
HuatUtech+TJnTQqAz9tvmU/A3sxlA9DtsEc0bajcAfu93OePt/4G5Q5EQk/BskV7dTTu2aj+FN+
FXr6sWcImeeI4BpKsRlLKssf4ASV+hr8uN/KgbA4ufjX2rK0X/OS3iac97u6vbuuoh9Yvxi/8IPz
kiyuyGMDf1Jfu/nIQidF7YB3rbJnvgvYjx1mUxUhl3noihtrwDWCeBWvCAVotIDYvtpA25Q2V1ly
nCXi6AnOR9jpbVk74ib3QnSJLuq8lTnvLu3Epzf+WyGFHr6q2acBQeBIs2ttUl2LDq4ojFzVUm/f
KpRdivfcUMSGujJ3Z+Xdj+q4izcOyGq9jZvKNdnNbtvEPkXcAjgmDS3DjDpOP4wfqG5UP37qyaCx
h8t74KoSoGFJU1iOAi2fxrUrXcgLdSvitzl0rmd6UFluyciDy/hyqKvPwyVQuxhLTtZTCCYOMIzp
bmQanb0YlZqSMMDlIUXJTmyZyFcrjuuY7+ztTB/Z3IdmYVNnzxIqaP2Kw28bmjW0425H5CFoF187
6Hi21/Qzpj91PSjgSNgX5kJPq9g1S3qTJomn8S7sL8I1LF5JCmfnTDFNHEWfl+hJRY3fU3OvVyHB
1ujvyNA+HPPqcF6hvt1U++Ey6I7qIcACtU4Ga3lTHWxgFvsH3Ml1sPMJfotp3yKqBnp/VUg8TOVI
esvkM/nxnavbb8sx1lKMskho/WmgvI/3SHBzO13VtdKCIbGzSZH6KO8QXNXqwGd8yg9IHI2GVBjB
0u3RVR99qWi2YruQ0UemnEw647MSnoyXwsQb1unrmWBAVCNo6dN0QDKWku9SvIYcduHaEI6DTSiI
RJR7S8aWx3pnsXAKrNPMYyr1SnGHUdlXgkc7CS4k2v+69OzE4Uk6MGuCK8ZwrGHJMuttPx4rOKV5
LgWe2gPG7okp/Xt8+T83wIm65MnD7fOijDVYJj877oKHuA3bNUD755OdoO8W+sGsRvV/pGt7nBBy
g5kDsXBNSc5QWT7somMGJzpVvKPKe0NmhF2XVVbR5/GfcBtBoKcQELQzSP3Z2zoTTjcJtoF4zjGQ
x6Bzxjgfn0OoqqABlpeo1D8u+RUtR+H2b1GWLGbNvP8H+6wwha1r2DEEGd5h7dI/4WujI4Jaif5h
WhGP+yTCFTjtCp5FcO1dZKZftEPA1Wg/Q3PR2SKmJ3Tn5Ozpg73Q7t5xDF1BcMx4qoFR/jYsHrEB
xeIVuo6YqpPOgI7iY3bmDFX2jMznXzS61NGJpJgiJ7v5MiMWk9U80nsFEd1Wjjz1HRZG4o788mPT
gfAio4Pe8yUdUFGshp5Rd1DE3J4HgDkfkRIBmUTknpjqrB8iIzX+4RBIBlqQaoWDxmdOtaYz2Bs3
nLrGMCLpMh77osOEK2sLPDHKg5XVHjWt2XWqN3/Jj87+54XoJCeUDu6QTeJ3jQGo/tWjPpd+WvE7
E0A5lAnBBJ33j7gr7ksInrScFIcVSvnE05/pRUNjR2MITxKOjzX7KaNhjohNO/kgjHXo9wakzZOz
xzIGeOu6tBg8x6fL7O62be5Z7DPbxV9CSTb/f8dGP40xzZMNIitM3WPGsdBTpWvIXPvd5cSleTr/
pKJmjzON/WpIyD6GTMqGbqGH67qlI20efBKWNijb8mJR6wbFwiohmz+lZ6SNLzVPgFbdoSe4S6L5
XLOwHicHiymFip745/l+cknlJI5NdL2D62Pqm6vX7F8oLqfUvS8BYe2kAhb5+8iPYDeOS95A08Sq
YJSaFGRLSfKZXAg1myC95nARV9p6/fTkV5lJW+etfrKtmdQiWFNZXZ5W6bmEm7P4zqxFKy7NGX8M
dYKrGErodIY5hTn7hI9seSTAz8umeIA5AoULFavpuIPD43AfCSs7YaDDJTJdoFrlP7unU6xWySvq
m9edjyko6wOyFIrkxNjBUhSNROTYh3aSP3lIJSQioGLuJXsByWf+tHldjZc9xiMLnbkT6WDsWSDS
Pccv/HJAekGfBMHFgPMIImqOf3yCroLqDutKjYl7xWTWe3cFmNxP/gZ1tEcOJk9gyF5pKIBj8eEb
1yicuFIt79QqBQST8MzVCrizKk/Z5L3NfIXatVIgyks2ll7Kup9+npTGQfq5OhKUtyGbcsvVWEWU
VxRo/PvQvmXs8veEdVmkwnMBK34H7P/gQ9gdywK2KVdyU2RLmXBCeLD1FV+wsiJ3CTVeDT/QNp7I
nJPuQIFldlfjw6zRp5/kBZUV5TAS4uM8pFsybVEbwV/8q9rg84oSkdfqeI0fi5FC6ha5vHn8fSKl
eJRg+f7tnx1pO00papanGMamdvVV8sQckHVmg1KeaUysddFz/8QQ8tiMNLm1JMoZQWIuqhYXAzvf
FCLvCyElN1aAgmMnxfXh3fBORraXpoNvYTJcVKZ2PJuaoPEZbO8itycCXpA3YIKVicslx7EmGncQ
V8FNoQ+mxB5ioA6REF5iGsUtUieEBWr+x242Ez7qnUYhuUSrHoI1EJxkdMrj2u6k3wi6AgNjpP5p
0JAXPY3i0Sboz/yzFBhvbQXv1QUNsxEQEjqb2sKcIYaZB72vAzjxnEYnakEl0Mk1803hYM1pH7cE
kO5BtAxm0Di7aGcTj5advfQNs6nOTLZc19nW2MJPw5HIQxbQgdasW+vIWg5dj9EMOTVSit5mlbtl
NUE1SP5sPjQurhnR3xdCwcbm38FQyk7ogf8mjW+KDzbn9aOyyHBgSIcSMEP3FpQJkiF/FjDFtyEl
EDaKk+uDPEvf7sJWyJL4hggBHRBKcya4kTWrsL127JRBWMa3iLHoAbvwXtefnewY1ZWaO8QFh/HA
WdMl5xeBsFRxKmHRVgbzGxeOanaKWe3q1WKdC6I8Z8DGXcby1Z59R1iuVdoH07iGM2O7tIErvClU
GvX1wPc9N+U0NmfOlol4KhhiQW2ipQ+K6XAAnDPLkNe4/HSaVPU2Pq1nseDl9PJ71FR4BJEmdtRJ
NSWQEqJqIX6nqCeMaV2qKxCQ3SWcswBqHxCaiG5Qxi87ZIymV62vru3y1LfmJDOZFlGQRbaOptvx
vVFMgx2BdUeBU5Nd+93bZqFrsAENtnKE9jwa/oNafxkRJ8t311rC0Bhfor6dlUkXJ5+fPTZcfi8k
pKV90GbyN2WCP+V/vakPgIbxKszCsEp4qZ7EiQTtRO/LvwWSU/NH19+oI27SPm7cgwfDxGCwLf5Z
NgSZzBkzo0W00ho82DhoYwjfzrmR1ucNBBfxqND2lDnLVZwJDvMH0aXzd7gucAet58EWUZWa1wLf
l/JZmE6E1+AB8zf5jwZ0OZx+FMY0MM/cOnA27u60nXZZTFeax+ZvjvNoERpVUFT4RkJEWOBsb2TH
t5cZVuZycLUlOc2MYS8sT2grk2UQQxvH5Lg+6EQCnYOTwZzwqxUgaiy9RuqqWAWaDt4ElgcFk3vw
bJHn+jrT7+bBnVRK2b1h4XOC1frVN5MM21lWYxuGsu7cqOVoQOHPHoBllqKavrpUcPmi23jvkUzX
TNktX3dMSNXUQTYRf8ltuZncSk+mo77d1PVeK+GywcU55OKz//UwHYeEU0/o1US3PN45u8NVS4hM
KPtBQ5h/f7PiAKumqhXhQORgvl+OxY6/DpBI7NI+QbDYg9iX+GGqhqQKmoUMnw9EGcOr635TlnYF
KdXS/Pc5fBsD2kJiti/AuHeCK2QVu6YfPc7e0AYd6ZgLHi53I90FNn2xTv0YYPys6LsUYuDlWztQ
W6n0AbhwNkexVTEREBHwxnwWhIjac2BO6x5MoMtVDASMZiqOGnQUGc8X1b70s4Chk5U/5BsCSba7
WMtofNJ+KrY0TD8o7nb4C2GQNoLE9sMCyo9p9MnJnqFshOF1vorR3EzCt3TQDNclsLyiXnVmEkZj
sTUWHYVJpxhVOZDxVR+Z8m7GVJmR3CMSEzbZNwngAuxiFsVDzbzHrHPLZUW1rGMQx9wzx0QV4HNb
94Cart70DixJlMWDIActxmbIGF9Q7HJd920XMCQ+VDZG5OqZsZZv41BaEZ0KO2BU0059F23vG4qJ
v+ID+GafvnKvZSSd6AExPkDtmMRm8+qEmP6xy84OOqcnx4W3Oj3W5KpxdYwAKXDWqwNyxCoWaAZ4
sZbTLhS792+QebSuo6pZnR/DpabyHg9Q70v6hEnizhzntASdV5eWf9glenw4AszQABXpA2YzOHyl
GQXmrKqPEnCgv8Zd1wRrWJvye3SYEfzvC9qWo4LEv9vg4FNCfiTCqNyak+4OMPCyAwN+aZc2cBN5
F8TSGJjmA1jRwzQKr8RJXFVKzJbuWMRE3HMJAooCbjZNq7gbBSbvnXEqZqx+tlhs4mMn9X3k0wkW
P/WCwBT7fsJMzjmsVXsvS1eC8Q7TdGn/kMcUHXJB2WAgAEKsKEvO2jXbAPlsyawEj4YEc3fa8tcM
/mY/zHYbZi1ZgTywHbaZhuoEfsuyiK3/PbiN7XSctc6rY9tmi5Ik/H4Dzw+JHMUP2YY8kSwnrIxb
Wdw3WVTZBEGhCKTPOmH5cj8FhDEoQn012dnDfOMSkpTWwk/zjJqSRuFfrF6SHQS/KskeAnbsiRkv
8Z0fS5wmcKI2H5emeMd2+qncLkAR3T7lqzRYi74P2b3c3pmCZiingi2HKxeCmS9RcWB2ZHKavZEH
yhaRLCHeIdGG1wm7eC9y5lpd5zomVoeoNJdnF93239Fs9r5jj+WrDgSi4RTQuFNQ1O7WdwsMUmrQ
FEnfSgOwr8YM/HSgtnd1vJtD1S0IWePM4TEYcMEdaNddDJr5h16RxmOBA1jlRnDxxmlMCpaIyG3O
hDtpg4irHHN31h0MFjpjuDG1Bz5o0fikzDzzXbl8OLY98U3WbNBkqhFYtH2WYiRda40ci6jUBbTO
rpT4c9CTg2e+9XicwsYuINJ/mnDv5ADcF/DZ28BU4UB5moF0/xmREEdti7qJMN1VCz8AFR01t81l
Xy9hvJ9NEv40zbQt4vyxhcc3OjEY+u8nXUs6nZoNGc4G2rJHN/gPRsP9NNyBOsJNQdndOUBNjtzb
lC8u7Q4Cu3PWqijwiZA4h6LoUEqNNvn7XFgs227TNpRj252fGgvYoHuOrkI8BywqOpbKpw4sb1Aq
wyZN9TiVTRhAHunb8v+b//ftOTSFKs2BcFP04n0hFGgupKtH2pubFOw/B9fueICwWfeeK1JjLxlq
CYXgDZEyqKJW3q6X2/+f2IwCyPux5q/Vn+7+J3dNySSE5O+hBgoKlTGn/sRuYnoUOIZ7vd1xMCST
7HEZSgAgbEQm2ulFW0G5DDRSTVfeAzsmnun06hlCv0MXhKqqbLS5b/2mUa2+DVxtry3KUBwSrBrA
WGo9Vd/mV8hFHvHDuA2mK+jmyYHrXd4X4K6fMIJowbRJmjI7SFvOg0OscfApY1tbpVUGy6JWWicv
OLsV9hGEQmaV/hxS6IHiSomR8xdg9rou9wKmF6WQObNAbwMYb6ckcu17f6YzzqZ+0DrdZwWQOO91
ixsFMWDgQS4tcAlkEI0SEZ6HPyJICQuz2zwJdSXKT99vz8gndYtPG7or7x/QV1SHAOgfzDfr10Me
aIVBJrJRAmDkGIQNoNd2l/4wlDl0B/67rYICZHib4uYBSm9zFtREUe42jo6469EHVVobeYoFc4td
6KHtHrR437klnKuAVdKrvb2ug7NZJHxMkQhaK4/dCs7HOKQwrTw6gVDmLbu6sguT8NIsHo92Us4w
bisEslQNHQemjfV3Z0rwlbd3+9ZaQswiNSYs9WBDgnBm2UA6zdrwxQWJNBUkrbfeYDS/gLu3XlIF
cTc8caIbBi97bJLGLF0N2EQVEi6fuaELSSwIWRK1Qeu2JauliIkkTMKSwCA4QPgXUrmjpUC0dFxV
21VUTHHtbcm9qEhOIHu4DDMFortZkz+3EVkYSaa66pEsrUFPs5Y7vQuY3FsiDBWckl5FeSe6pLg7
mJWoK7Xv+NNlEOqb5kZWZCy2zC2hd4ueCOWCXJNueQZlmX0gVnoHB34HR3DNUW6T6FkKY3QNbs7y
HA2QrxoZPHLMcJqbZe2B1KjO7S4Sujq1iOU9fJY75kMNKkc2dqKW09nCBcKVSmDgr2NfNTisnL+H
TV8L0hqbWAPb/0zJ1vMcGTdFQ8UcFftq5I6pHBOBQxAghOPWjT1ibrJ829i6Zvtrt/XiIxroxMAI
xbJUtvwcaDeN6T4oqfz0JYod7RSQCUVwYW9myX3tkV2s80oGwAkNccV+psnXjBAf8sIa/kneOTej
GmUcFUMdmyMfKnE5oSkqqH5p/WBP71sPDPcsis3BhjF+Cz0kr/6lMYAm4A5jGMkhDM7pwznmo33/
VWfr0ze7H+3Q3laIkGNwxS+SxCWANJCEzTmMULCp+WQ/5Um8KYZVhQ1hait5g60xpoJV/NjkEnsk
NmIu2C/KA7AtWz7G/JJmZiwrywEbuC75yvnulOZTYvnf5SVbHoQlCTtv3DdGlTFwlrAJ66nfgtuz
f0P3+BW4kd5xMq7G8b6AGfhF3M77MS4jpkVEA5tlmqTfOTLFLYKQJiPT/3okj+Vt6cq9057VAtB2
t6Pm8/ODVWPZg0cvoWUsnVbG9K300DlZ99iFTpvQlY9FKPDn1808mSBUFYpVlKUNLLyjsbRR3qrB
Pg98x2sY73YwJjdT3Pq8+bi6P2srx/sjJ0xr4QtmjsY0lnJRl/kHhpIrczxZEZbkz2XGzcUFTEcG
0neOj7pyFEfiHQz8jnlusAytaim87N5M4cjGmwwu5zQKBQbXcPA+yr81AeAC7LiGyEX81dM+X99L
m3D00da7ViI8oSltxOovrlsEiDfGa0z/mhtoYkpQ/I2OCvXnQquU65A83gZCNcCRk82jol8Qj2pi
aniPDH5CADI3gczMA0xnO5aSSE/FO737vAtta2HKiv1ZFuQx6bLUT/RoBvwZ1QfBt1Sl+i2KL0UL
iLqOx2mc0zpVc6ys9+EdTJa9e3+nWYKWoBaUy2vJf3rmJrCwsEw2XsLARBqmZPf2r/idvHgKDZ8f
3ySGSr134CLxHdglSqd+PJgjQSI5GjPDcnX+ypRLzOWAjgfpLkJoybDAEBO1SejYDXh3HoyckDl2
TBcgj9mRZpCaYVbH2EeDT3cT2DYegSdSW9QQ+UlQxTpLAM+lDn0bUZ4o1HWlJC5Lt84c1Ja0jTDQ
ilaFs9+1fBLLT9o2xvAajpwQi7UBuvhgO/O6L4/J99p3rYIiDyWNZ3xNo9cZIzyg7iajl+/6dffH
7/jG2Tcu66xv1yI/MlmlPOVKqqsQz47aBN6wEHUezTqaJroYfLNK7mVEZtdC/H4YoAe7N8HGOJDl
K/XWKx10yCXFBh03AY8kB1pQABUvETKiDzLW6DcxWbjxkLHakKWxLt5BsPdD1/bEquluqk8Rm8yg
3enni2VVlIB/gfxe9vMPSqrZJ4c6DkjKkKgOyE9ASIFpEIHq+Ezm0M28Sf0lRzVi14BtNRvWqjhC
oj9pXBEI2I6nU0baaJIcdgoCZ6nYKqq9lFoaQhHk1iovLhVJqdAGBCNdyAQsCN5o35UKArYtO9IY
SqbrXU0q0bWeu+LdHRtw0bttMen0+IQF9ZzEjsopkAo/tPLv/jNTDWmjzMue1FRQwmiObTTF8e8g
vHz3e2/ZteEASQQYcOtrWxZw/oDHbRbIxGy4H5WFYHdkGOmbmv1R66D4boOnjamEmP6XFG0rMeBT
k1bH/pk2+2MMBxufvuFFo6qXU1a49OycY5gEJTlY9zYbZuOx9XbckgnslofsgZlqKWgG7LrCA05R
BE/C1vLLofRtGidbkryGYRRZ/5fG01dwwBwVTy8vlQ3ZSbu0nR2oRX2F3+PYbZeZp0BePfx0JLbf
WfuZIJtIHzmJ/u8YvJAWA02vyjvbKvlJVkyt5LkBYdDTLN+UteqFR30furGDowOUD5x2n6omnw3K
K0gnc8GtKlW/BehSzEm+5cYJHA8AcN1+10up+3DD6wtV9fnH1Gn4RmDCyVKF2SaXN2IBXKwfa7gx
8L9PLM83fQMTfmy3hknhGv86oCyobgRZD7W4HGBypGEBE5nKSnBpptDkNYkVcp2stGu1cNKpVpZY
0ucQORB+bWFI7YhYCEpoukmeI5q/BtY2hryJRMJEgNPcmvRYfmwruQGOe10Fvyi8deHMrVNVOfEa
8nSrSrkitYseQ04TZbrJI7Sq6sSC0jY2gKU+yF6emVuRVqPWhqv9GyXCp1gnRmNm0dxVQUujkzpp
f2X3Qm2DXa78HRYRMO/LLPgd6ntcijdr9lKa4sy4cVWFyd823iV/R9dsRZW/X0lqyJgH+UoFgzQT
zYg8umjzQP89QdCJcZy2JaRp1izkzwhqWkU21Eh71Q6mpc0nETKe4eCoeELd5eh1i42zK0kUfpmc
7LigXVAMH+X9hrewqU4G9z/FOqjMAMvFYj6j0p0d4Tt64KIYMO6LNwf99g4uUeGRrVVFHJ4xkw4w
23GdLJbVlSPpfif3DUqGceZku7/dAVg2dNptTh91UT8tBFtMnRJe1tsD0EEGv74LKwtSGU0eyaQ4
lzXnjxvuFh9VP31WQcYEQIb/tbdEdH/zfFK80OLHwIKfN+Ps6kEUSVYISjZZWX3TXQxx+BfDvptU
wAnA35whpkYhkw/rQJ0co3l/IreamNUCS0pQzYrsxPsAk8tppVwCda8yFsNbjjRteQQD7K6iwSEa
8NpzxV+Cf+94Tq0zyWexhpxnEvdr8JrxrucHSrpfYHyAFueR7kUsjLrvD1D/qPKeuhr6Vx+3CYLT
B0pXBhG39yk/eaZ5092zmxo6LrOCBw7/glPu++9e8B9zuMr1HecTCuN0aocqZJdUrP46MbwgJ6pI
CtXuO94FXKBHYlPJfQVkjmbx+m6bmba6YF0VfVmglKuMno07sXSzjZhVm0SXpiqTCBzkgX+HCq5h
wrPmlQnfa5n9vXduVYkXmHLENDAqQ0bhokiV2CsInI4GcTsRnocwWYTUaZcZ3KQ0bR7YkL9WOVGo
5Tt9BawMLW4QAjIwjaVQ3ZxG+Y/sHVp/tma0m/Vk3YbdayrwZj7Z3AlwxuULX91UixOLda+jdzXO
48MkbpiAO+YBsyx4ZW2dpWEFe3LB4U9H1GRc7bOogMJASRXaOjtLPs/rD5F7MUK8p8b6RRsTYRZc
Wbfi0ChgTuG9fJLqxeH3yKpz5ym0h4N/RgHoHCY999/oSZqo5mmiAvywarwucGmLdqkB08dfQIMI
8+wUpQv6vdXBbmcGixXG5xT+eE0v920xs05gVxoTDoJPMnWx4lQcYK5+xEh0Yu9EN5z6/Gk/BXnc
8OyWSvFHJ34/V40JwYsqugyvBdU4yBXLJEM/puXhUHIcQPbNE73KxANU8CPKQEVhGX1oPSqidNfQ
TU8J79vPP8/Wl0QuOD6gtCK5jHDZx7rPF+i1z7FOoU/Tkktn2GXyng8uw++tUt/759eV+SD2bVl/
4U0Y86Ny5fnT6r9gr5pBxHaQlaEZKwNKHikS9ib0WfzIpbeCh9YW8+xDWsXnZlfyd6R4SMap5BuO
wb6s0yEEqfO/OjYbZRLOvmiy5AnTmmeFAPDj/sttUM/epE2RtAjSP8NBvyKccXrmcKwDZvvwB7fK
87DRG+EhHR2SsG4lBXDJS4TFNER2UDxSYFoybEDJIX4NYykXxTg3MVsS/4z7CVBJPKgwLwOYJ7hd
UB7RVPXNsnHUwzSGAIf/JmT/Ieej9hlIhmCeSDtWN+QRxkequ9n8U/tQVAIn5HPNWwdVxZwHV7m0
8uui/nuwRMR5AV2j0lYIuB11P4Bg1gj8TRZ6DuhEr81rSAjUJvArB3wGO28UoDZnvHQ08a5CVoeZ
OkbOyAQWqWVuy7mO5lKbx0h17xaaTZhIveAou2vLtzpBO8kbKv3zs7oQQY8DHvua3k08Ra7fjvkr
NzXTYg0wvlb6xhvAVzZor+N6g0boVzDY2GkMws44jJietrI4m6dfF0mE0gqs5PIA8LsgSnpBXgTc
UcNbkUigtihhO/S0vkwYBQESLPgB+cephKcCUWtAaDbtNpQBUYDiByEu+315O8vJFbDuHX83Ylhi
yLxzUj530X52bKTguZZyglPYSEix9VrHzhWEo2a0lhVrrTsTqL55AhbPoNlKLU0KVvpeORKQ07jf
nnj+1yjFC19Dosfvop1brNWdM4UL6w/DzBMyBSv/0KcTue9WcVL9z8iuUT5WJKxHZarow+BD1L4r
K0FAhY6aSRaCacd+hUIaM6doPeOYf1YCK6CHnQTlk+hphtC16mZGmWHnBf2KQL9vGnv/4vz8ZB4a
Wt82Fq+YIV3FvBP+c5zzKHE/yL3JQ+QU+YP86Lkn0jPlroKN+MX4tm9u952/joQy90qBe8FtMOYO
2MbdZdXS5HenQDUj2mf+MC7PcDaDVwIFsrasBwF9tUczvdWz1KrI+s3DZofqzd5wlHrwFKkVqrcd
ZWQ7gTY0azzcgI+nxq2HfTlwmNmmGZr0LZjPxOBruZC4U5WFKLeH9bWUz8nlL6fKm6v1VChUNLJm
XnPdF7SmkjuLA5uqkr0nmpjoQ1o1/k8tJwje9aBkeAw0Wh/H6LT/opvpMjQYJqJyy2L/il/hVEEH
r3mQ93Ekb96HAiYfJfTX4WOAvsOQ5VeOdAgKIFt4XBIREXvnT65p9x9EJqBBUzSul8oqFYAo3yo5
K2lx3MNHFg/p/004rsVU8oXdjcZv9jlij209T2geB9lbb4UFEurnbKp0RT+NsJlSyzHeOtnU1hHi
D2a117sIk6EZW1W6EDhsBEdYOSnWnkcYvTxPWHSgKSrDmruBhOA82dIsFY/iNr1o2al96UsyUTt3
gKEZgnqoELtLHXjelUuxcSOSdT0pZs0Vdru7vBDqvTTP7N+8KOoCE2APXay4LWHOd4TgHdcgQ7/S
wYPKsEZuiQWRu3Zt+fPtC3unKqIRtSky27lhoDY3YX/MyXyygB3NSf/iUBQY6OZwHjBMeKH3b6MB
/JmTLcYDPwkonvXvGEz7Wqu55h8QKhTCcL0QMAXSoHxxRz0Wigf5O1dUr19CPj0RcBJogvv8XII1
PVYzf0itqVX6vd3m8IcywAHV988vM/pNe7TgrCPNmWsY478KR9qmENNWgO0iBO+eFSf/MGvy86VN
VupLuhNRUs1k1NsQ0waMJC3gTgdA9lKqXy9Jetv4xeAoILi9O9suy3cBE++NvZqpBpOxybNJLSpm
EYAcV7+MntFS5aazK+BNbdL+PjpN46d096VcS63CbrfIg28pDl6SjDoV0UOAHM/ajStl+UnpMKMJ
Txwp6EWTwEHZbrvjd+Lz3yTkELENq6ntLM7sx+WTZ2ujMAU8A6hm8Gx6Ysg1kaK3HuLXvZFXBrg1
u3SANcTmxbAz6ADddjy4Bfg98B9c/cNJ0od7lAomnaVfV/j8QWRESfcyoB/OKcrIycRFn/AKJ5cU
FNrtsKAEAeQmpZMlEJ1jYNBmWZpekhBYhCS9sp7M9VerA2wrcLSmYvl81CbYN1DPpY0gIgSglNsW
WKZha1X7LxxhNTrDtB489TnUNiGueFBPmNRvGBBhxEMdfsgIpKSnTGwx5W/s4V5IuqVVhZZKmwyl
6Z7oERj7+rqUwQaEZ0Cti5aW2YGInc+OCAj2hVXdkF16J+/TwNdYyUBKknqKHccMbrmPINl3mxhU
xjlvG6rRjV5Tx4IZeYnY+Mk4bknIYPmmdSd+pbGuqNueP5xHy3dUagem9C+rFFt4fvsafe8J8LU5
+OkoIw9i0VVZbKBmRsfPE9eIUskhOplon5PcH7RxeuuC88ldzVYn7eSQ9NU7jc8lOD06onEsRyhi
CE0VC3BiGKqK2ifLlVn0yi5qveCiK8sy+p6xk0Tkgy2lf+o2+oNCzd33A/rQ6qAqq6aJiKZT3LKe
LqAWEqkiPqmD4S76Vabp8+ySWvYVnBLkgYrZ+Ry1jyX4/247A4PPVMBIjmpKGSArv0vrVvNZrEWf
9vNmF27XSnE4AAA6q371aXfhAOvYOphx3u8T4rb4pg6vVWVmIpsT/GehDuNbVJFItr8mefCp/ukc
vqmqKWDbUwcvaazhaGIDE2IPxzoWolOC39YS6+6kC2t8j5k0yKT4xrlgEPryj18EWtI15YAHuu9R
E1df5mtLAz7WVJ2HMkmDOrEqPPPkKG37MBtUMfngXWd1lZxNhr3C/osI0TX5R9CkdPy2w4cFk2HV
hPmB7wtrbEyacXr0f2PuW5j2SmOCd41xLTjylSNfOa6HRlpEM42oEe8D2hniU668EmJdDsGer8Gm
+Ino5+G3M04U71t9cKH37rqJQ+HOJl4zEVZ4pCArJS1JOi+hToi6e/P2ZpjASYXe3ER3Hxec+UoG
2XtqTMWCcOMLGfZMBPumIiq6FT+JubAA6KHJAmrookH8mzPLJrGhJPiH93lXY1nHTG8Ii5QFHfVp
PMJJUuMTxW/x2cZuD+Yx2eEpc6hXJNIljaPCMaOuNKc5NEQBUEVCfUEa9WuZiTSp0ylKfTAxAZpr
syFY/yTZjkTtO7mIkur4DAhQY5YacQ5PVigAlUmM6KWjTR7g1pY3XqYDoGAafSz9Ch6xAG0LhA5a
J7VA6GxotqmJMHXlbBk8GcOEHGTKYSG2TOvJ0iHn4S30bOMOywEcDI5CGIMIbizHOwz6pXHWkDpI
1hgXp2jg7EdXpWTLp3EclBA8M9ROZqf9CL+jBTm0Yz4e1Nzq0J0oKwaZsPi3PET+dMYwNzsTw0v/
i7KS+sCZ475hLsz5+rSkv+EXOHey48CyHV/4/3DlouAVZJTp4BEcvqySdF142BsZgXP0DN3tQcD7
kec0qaFgkcPNicPoos0NZTBGG1X966W3X91fItGyjvQuBbul2kpvlnS93zT/18+r6B9bH6GW9SDI
BTBQZ6Z8yFjpU56cqsMnhxqt4gWt5ZmyLv/vSOxump7z94khUm1gSjN+xY51YGwYPGGaoy5whhm3
pwoZSTYrov733HtlAPyyB3NJOAERcv3RP0FNDPEAfxHwJ94bDnFuYp4Pq4VNvp7eYPeRrtOMBkG5
TG+GD1lQvssam5FdQ5oeEfQlybPXRZhSf+3OWFSJNrZqZVtF4MyjukOX5BUP9C01Et9o7JjOgDi3
vp8zRi4bb5r7qKUpyWmLQrWMK3KJLGvTf8G2TKGQeTl1Zjv3toYvfBThk/BQspmnHszbgBf+2lYT
UODmhzKinubmcGTNOlrAtE7B3RD6e5TFAMt3Ojkx9tjhSm2CZwdopS1AZ1HwnDZ74PoegeLgWpMd
6o0CgcPprJ+I8hdDzo+3M4zUDoCtOU56U1DavyslLmBRM7hMyTOI01YPuzosjbo9xcQ5LIbLkp0F
1qqrVed7tDC8Uj0PalRQQ5IDWds41Zx6CqiHXJ29rhn74ivDOibkuKBTiXLBnnw239RjqeSkQ2h7
O0bpOStty7NFPWO7m7YnZiP7kQYSUitt1O1FxQ/G6L9eDWhxFusEeucnLH4QdMD8h6YisWkLWvBp
mdSK2L4MNCLEmt5ygJyBySMB241u/rTGqa37+61cWP30DCxvrqYx/7BBaQIIrEUsvilvZN0BGQY0
XsmGfek2ynKIh8msOe/9rL2fwR7iI44mDGnxgotgWQRo2ij/hHb9+/1S3aaSmUhwjXZ0eNQIhrpF
7wCpv2GILhFeWNq0nwnQ49AUxoEzVpLYlMJN6VugcMbnSfNLhm5Q3ZXtCAimiVmge22b5iRCY07j
Lu56LzAlY6j2JNovtsOE4CLHKbWwhNqzGL+StP+OA9ez/sYsa8Not9uHb20ygL8kX+ECkenupSh0
ljc790jQBLAXh2/bGqwOIwmYLeEn6x8SnIlTLvSxsjjzX4mQH/Xr12MIx779jHdmAqhGOLLbdd0L
HvrWaiecRtzMErgUR61/RZ4UJGXDROgTTnMLeeO+bViK0IHHFtyjuvoyX9nUitSed3Sv5XmTWg93
W4kc92VvTOIL0x/4eQ2aEEh5Y5pIArk3wdFY9S5q/ngCrM+BcdceIlmZnjJjQqTyk+8Ml6RxwTx7
GBZ56GuOyBHQYK9sjCRmj7swG0bPvnMIIuGHelBl0P+V1UpW85z/LQnPGSWiqAM5o01r6jUFx0u2
pVC1VHOzHAYUyyvUPfq0owDSdU92kSZ31qzEb6E4HA8Ia3V1Ovfb6Fqu9mMSIWEfLMLFtoLueKNm
V508wc9SJst7Tj3RNdRsnoWdjCppz1kvHhhzm2yxSoAVSF1sIs78Dci923OZc2VudLravskzP10n
xGxtPukUlEWMCwSg2IBGKKfJspBeD2rVZIIfw8qurLPvqgnvLojiwXg41OKSKc60PP0HwuxwFo/O
Aj/8SN35s+m9GMh+LN3x8O4H4e6WsSkKa9QJ48NRwf0sm380z48191XMuuDs1IC7N+2tSVpUwJmg
+SFeQ/sX3l/M3d42tDRWM5w8ZBLWp2QYnhM10vFKl43OEjUBaUSytjIQehJi4Ck6oc+8c3VFzja5
m8jCaR5JGTYN2FIKI5hUpbQEMzCbEihHD3YB4SD3toTq6ceDm6f1rrIp/0XO/yek7S7FfMtwaPHG
qG9c1jCD4Wvg8n4dYcTbALvKIn5yPzZLccXQDlWc6o6iwVUHs7Z6Ev1lqBXuwqu+fNPVYcrpVLZq
wH8kmHcspD2tA6pIzR71KxWqJjOkgKqbM6TcWaiSqe36BJ5fhYWMInZgoTibSJrdZXFMzHgIamQz
+1FFUtrv6DsmQPLtN4krdI3PzRRNYz0D974IazdaA0ui6tJCyRL6q9Obgoqg9xVexYDcpQmYSA5H
2diGMp3XBpz4E9wsEhWY52IrtnKEnSEZZLeur2nB6vDqg/PdmOTF2v0Gkjdxl6udOaZeFYg63iwn
VJ1Nk92WKhN2gKGUtmCNOAY+F20pcjfCKvNmySZc3xcU8Dp/2U0ia/esfCzgcLkRjLjw71qcU2Sv
sxplNK9V23mGAOWRRoWDHM9JMxfLVaF1k/hnpTfrIA+BwhjxwWKT11hsaLWFpLrDVV2MyhbmO/nN
ZjXYLG6FuTz45iOfSctaXVTUter+bZB67S40n2SrTRXBrq1v+1gCHTN86Y4JC0KspTmXA046Sdxl
0hbNuYhi3r2GrSZnvjhR5UUxKfAX+cO2akVW53PT3R9O1DUg0PNAD+MapYJbyyJkMak5SEKSWfaw
IRPzs5W1Bn1gH2btgqP7YEzJJegLCTH02KTjUPPJtwv4cI4xY1LKOr1wW2s1pb6WlL/RLp9KCnWR
gvJQkR97AON9RvN9voqZfIJETpAYekB4pQ9Nv/lJ9CEvIovf+fVHJuP91vUbuqPXMAxy3w1Iguqa
ciWS+cYov1B5Uz2svDHy63MHL9TKV/iM9+EC0Q1LlX5Rktyl/ut9wYIWVmv8pVhlRX2MWih3cbkb
FRy5nB9UgF9uWXgHPw+NhVIiGj2ZvoMRY6YH2cQSSx74HV7pDsPGV2Ow4sDrNo6Nwq5IgOXLqGG0
3Rp2EQTxH6sxlCjyFnlY2qxGYaQ268N2tDS4sUeMoo+i1wNh6nFFVQ9YvVH2pSZ1oKm4/QMboZIi
zjJaBFDdQI9HDfn7c/7bzBNYGUqYWxzaZgjJquMqoKsVaFsDPenxEIQyG0HefPZ2z+otkvpUeM6t
UeHD1uqZ1BB5UinUAxCgaDfjshcDZBSTVxwK4ECqVYHm5csoAct1wZK+icTz06HuKYFyJg+DALEp
HbYATrzbiwbdAc5Bzu+eUmFSFZ06WDMN6l3z9ZrWHjdBti5JMqgxAai0PkS/QtpLkyHsrLLvMVzW
1uyUEWK7kN4+7kAkTgXo07vAd6p67kzsonwU25C1hzQEDvB+C0tHC5ckdFxqA7/Y+6IPZDH6jSMX
8YFZI9htPcwy+9aXj1dEL+DAYdxM26M6lKWC08XVZ4f5asr5P3vdLE6JCip4GlVXw7Wa8NjQYmw4
a/MgnOxO0AlPKEITex1nKWB5O321DXQNiW3y3xOMLahZ/MZSgpcGHfL5DSfJOMcQEqf9QOXTrtVO
chVrsfIH+hMjOMKqrb+SVuPtMqIbCIbqGaNcKPfduxrHcRbMkbcuEfYWGCsQamEMRvrAYfNJT8Ko
HxgePlP2Bn4fvVq9qHiPbZjyG1zi4TF2Qz70+lrQOaYhDwzTeN4n9JtnI3sWOIBRx8vwP5lNp11/
ZyYpNmSNTHO/ox7XlInuXHLae4zpcRNL8fPzw7MtEz4Zfo2VcFnnf6Vk49m/1/gmsLnZ7UDqBdtq
O8gsG/bznKIdq17qJHrnxBeJxWMO+pZQRX7PQ7wouT1esqgw3UuXHv/u46+FzDcqipYsCCHyI0j9
QPKyYo81Cheq4jO0lJdpz17L5J+a/8TDoDBERP6tpWV22KZKN+IsxX2Y26+hPlk/EOcMcdKLr3hB
oAspykEBGp2gaD+3hoLIf7lpZ2V3fw7wJ3tA07I3FdoFjikJ5/NZkQBP8GOzvICZO/LOVlol5cJd
eCVinE8IOi6JicsCKVpsOxxEZCpXsMsi/FWwMK5hJGx5pMciImQATUNkcomgPx1ykPuJPp6waXLT
g6KMGssRJ2D7O4Nh5OdZnKYCeEnEcx/Uw7QuN55Y2c0wCA753A2VsYt3KoSJzr0qqE0qnQ6AOiRt
qBE4dBqjnulCTp7EcMqiPqrY/tUe/xvK/iHSCc1MUeOFJ2XqL9nW7NfBmy9whTfF3+D1a97zBHRs
0wLf6xt9cxyDOUKxOvaXHEttYYtWk/9GoMyzrYobYUnbXKDm6oaMuwDqO59oIxFbKu6Oeb3Obyp0
RJNZYdC8FaO1fA1vVg/vgMkDgWdiWdVSiLqDUS2a0t5E/EKfMQXc0EsbYWFfZNkQgxr6SlrSXBCy
8vr+zYmUiT9cvsRNv4yINJQpCB3wd3owS3m8gA+EPCAt0GFg5nCurptfp0PWrl9m+M50/dfarjeL
R2ybBDgt/fRFp24r2iWGeoCCT/XCPdTvUPVScYg1l6hYaBxHE9AM8kpdoiwYKtz4HvfGQ9LTKlWK
aKPd6TCqo2uWrXOynkx2VtVnwfgXFq0lNFFiOS9Qfcy933c5CLzmA8phPu1pieLmrFQXUyIG1UvN
Pw/DMnRNDfNhm7FWYN5xd5+tQS1ylxxo+CdAfk8JC+M4mL9sCDi6Gb2ldzJM+eminCOYP2VA2BiJ
ZLgbXlZqCfyvNoq1vGV5CtP2JvfWKivpQKrisrOV6pU52SYA4KPLmUWKqA7R04zp6ZOQ8eeWufd4
EPFb7QAvQ2M5uhRBq9/NtVqwqSKB01yfqS77HPYdvuwS+lpKvpTYkZOZwZZ2RXOwMMs7K25tTlZ/
XM1Dtsb1NNW5YssDV1dgBAf2VfOm4vRBXMvA2Jj+WmxPUswvJMHbVLpgwGuLPjeCp4jVUML+QRKO
IV9LHgXc/3UzgIpQeBwEqEMt9Qey7mbEGFjipvezTt/iLM+V4CYlOVOdmYBws/jiJP1eV5B3uvkM
NLoXFOmFH9Pp016hETNEP6AOC7TfWtQFNebzr3wFfLClD4Sgk+fbNNQUwYUktA9eSLUtcaxSPmUp
abtX65UzYM3RjbG0EEXkBys4RzoNjSzTPoZk48tE0fiWPKSZlkKP89fFRl4hxDQ1cNDx84W0v4QK
HV6qsOOuUSioTqjO7BxIktneZjD2kRjKbAktkP3/TqbaT3rUGb7G0c/3/L4eXLR7Wz5gqpBvEqGv
TRPIjKWhNmjWkBBYXqplvjV3bDqgLhIwBCnuV8JCa2rMHhsiVJaiS1LPZUePwGdNqJB/zxmO22/u
5LayMFTearhRoJx/P/BcxQ0bVcwbQgemPu0oQ7VuHqtwPEWMp/L5235NpGgZcffvwajKRp4jnJ6W
Ao2CmyO4CxO4p8/caMplHd96YGzl5TNZCZ2snykv9tNVxqq6Lq8LTws27Qdxz8SdrSqjEyqehcCG
Key6Ao8N6HiO32k7XLBjoV4jOfro+/KAL5+FA5KP39Xrd4123+VnSfiG76rlTB3ZmcLLUlGuw9PX
2LegdLzCHizCVODuJR7SOWXHMQEYx27jELO+fe8/aL1PPbFetxoB1g235Ofakzzo682GToMd8H5C
UBAntkep8sGv2BhjkenpVp8gaSnhuT5SpHKUE2Ts9YhZxJF7hJRDYBksjrrf/F+/cWEY1wOLDHyN
LXDe1/NsP6BXcO2kwCEU4+p3Cn5cVvjNGBDkRmAWDL8eawBpxfDpdxkLnJiKJatlGN7PBT+RbvW5
o7FIAHprt3PAaoiXX6EPsw9fcGZpoeHY4ZrRrsOxGbIULNSQjmcbc7WzT3obrCU8W/hfN7I62GQe
1WN1j/59F5WZhZypZPqLGM4+4332MffnjgPJL6pqvioCPEtNuH32g7YDS8XnA2mRuSgedVGTS73D
lMjBRo0tQgEpfZEBVWInBDXbZ3mTJgSK3Q73I0CZF+TNx4VBZlF5Dx/lwUOz4pFT43q5MJP2bh0M
a0LLOxvpdQeXy/OEESrdUf/05HISOuKDhuky2MNTZDX3LZZ4l70Ze+n+5ewdPguE8m6kUjCag2m1
vS0AcNXVyOkaKGPrL8Fxq3Ygm6jitpj5I/oVqz38bmfz6QDNLeNk0wl+c3lJHx2KN49VD9tzy3MI
fbMrKtbOSfxgxWT8k/pLsyasITpZ1eYQoEiJNvO488jnx4Q3jODIQAMoJjzTySVP5sTOk7sUMtO/
0kW/JQp5Lj0CuCq1j6AQz85CEqSfLp7CxFJQ1Br4USyuLE/pJ/lWo3cdfkOAqiDv/7tJwbf3eo/T
7cEzKbhtxxlu0QcOWwIpRsrBSIS+zJRekF7HHRrN4NujUXokwb8PpbRWEUy5C4gYRoSQBh0AnoNR
MiyT+dGppqhvLIafjWGxMa/eIZtK4pEjJG5UnbFy4/bEr+mCpaKhRl4tnxqc/2I4qwktzsLBWW+i
tT+U896z39uOybrpHxjmBBYmFB5gDTueftnhhgB/RwMg4qkLHjq9stuWMEMKh9fPFaNV2849CBFF
7foQr7WDn0tOvS8LH1EJSwHlrVqYsYE6NK+Rqu7pcQ9OQgE//4KXa6zeD8DuAwdZbUBqc4ixPEqE
XeO+3tu7dcSdDNlD0obPqNTIoqz7G0rI9uh3z53QhGFDW39UGMfcL+6QD8edH7njlIy+fa64iO2R
8eoDPxMDXNg8SU155oc/C90I68m/QFHr5hOPjsxvqb+nomYOtb/rMJxWFgNB9HjyfGCKq/dZ3FJw
G8edxcCuslRdGf3eTIWRteAWftGnhPSb1bRfzo4wN8Lw41/QRgok/2kfWwVpXs+SBRS72co+NTh4
3r9eBC/A5KNvLR2FIoiQBs/myOLCkYs1ReeiibKNW/UMgKsYli7n+qxRunM59W1HuB3CLFwIPf+/
lfsPn+rQWyqmR1nLPfZcRhGSPXAS+K3FwYbuc9byHGvTj1559yzOTl1rDIX3MA6pnYKrjVwSKoo2
toA0S0OczGuLTRTtga0QZOHr2O2114Fm3I4aNZc8BPeMGxIB+/jp1kH/hDwkl4EHDyL8FWK/jpDo
Sl6gGT9wAqK7Q1CqOXkHwbrf35uWVgC2QFKQ7q0JLDZb472D25VEBCRReaBfpn6GnK4NYmXOo1/s
Nu3g2wrmQmErr8t3Tn/tn1ElpRNFLa7L2qi5cshsxIDGuE8C2lW4tyutMa+I7/cbk6zd8U5tQQJN
eSVSSR30UAWUp8z3WOOK/0WEjKzePneMz9+fm+N8YL7bHkmFfSC0lCoCxBE3QKmWxqQssyQSpW2O
upNV29kpBydX74g0PQB8GNr1ciZYZrivZxxLgYUiZENIAldtvLamQgDi9mi8B6QHzgsQPy9rhaqJ
VltWisRmWzRBK4oIzfEiDgl1WP1rTLvV1DhVF7TU1tTZwknsXWER35OCPyituD5jd1kXZdDBEx9F
OJgoZhx8lLdJpwrFdOyy0NT4INXq41AtsFGPacL/fShW5AvCiRo/xtnsv2wFNJ3ljOTxCcKMN/+/
dQQDgXhERwDSK2XCNkZLWT4R4QYUj1gmvG2eZStzykdrUXuLNCqWl+JDjnqN6svKlDl0Ub4/pYYl
Hv133JHw7LORez7dCOT55LWBdvry8Ue33J0QA1eL+UNdHDdq4/pgvFZq/zq53CkLYf49ub2OYFpU
5nT2DB+QeXeHWWOisX4F/lheXnCYX/k8q5ETPSzgXa3pFQtI90GFOdPfFIBKpoqY4KLRO2eqZrQO
28LX5XDk1hf0cvHNFmftHzXL74pZT4gngGtQWSV6IsZiG8Fq8R8EKTvz+O0ppLhd4O4Rp9WeJiKL
V2xOlZwtH1XSr5BqeiBkBlk66sAU6cS0ju1nDPFX10i7lr+CdHDRhK/+HdX/oSRhljtCUjAcJWF4
turuqAvB9uZa23GQHzQ7WHnZjlP0L8/sLFU5A03agpVrTG35H2aK+qIqZIS88PKu7v4t+bS1xq3v
t1H+jZwkph4Jq5uGIg+cxFzKAXioZumarQ2DmlHZLHkRucm0Za68yqhD+/ELAtl6b4WOrwPQI5mu
c4KGqNq5IxmZYmIBaXBc+16QIWidhq/2h9k7Kpg2fXbbRt5i/YXmcKM9K15EJnlVTScFXQc/Omlv
wQ0Q3tRRoj9E3C3rPjRzzofhV9yH0MldUcZM9hDiNFQyhmy+wQx46awN/vLqy3S2RWkKOj5oIhws
MtKrK0R/yCSN5TIPArhRHxTCX/5lAOVX+axUVqfklVAGDDEjhnaJKacMkMLXmxkVpIQJXgb80l19
94VEbN3SvzImduoKAlQFUIE3PW4bp4V4qpXeSowbiZ/nNeIJzxHbGPn80Qg9ujVOECC/zsiCk9Db
UJwXMbVLzJiDScqwledaXnmfbvdWVkBaX8Yindk535aD8KtF6FMrHNNuLn2gUZmbdzJMC6ckNXAO
ZwTC+zhfkfHqp/dMd0bkcTt9iSAr+QE+GiJI27PGglee9eUOsEUFm7P4zCnfGGAcuVrEp3xeLqFx
krnuV90O+lr87JH2TYJT4e6DUy5rY5nEVWi9SL5MzJBKbi/ybZsJCREeCiy326QZbNPhDRwmBg2i
xNhckq9Jcs1uCIvswOyGmlLTV3C5J7o8pp6HabF4I7qOVd/Sj2NhSfhTDsWrnF17suW7EOhQ4Fkk
lj2omkcYbpp3Z/FiCJ9W8W9DKzBBu25MuAYrXai2C+LX4El4rkNgRAO8rXy7cnRVRLVMloOjpJ8G
b0r+vJe4L08SdlXHj0fnPIg83fBv1uaLmGfYZXAgEuKIPYlx/r8CGyxKz9elCMWKiW7bXN4Wx7sl
M/yl/P0kkLrEV7c7mS2sMjJnX6opPjnPMvPmEl3/t+JC9vJ6UMOzBT0u3N7Fsj5YPGMA86i9Wvjp
bSvP13pTr0X7B8oFUXFSWr/n9XxneIC4LwYasKoebfmYLwp+HO5lbF21q+P1VQOcwrdq9h13/H1Y
sY/UdPl/5OwrFwjpzZXOfca7I8FiAVY5Xcf6QL81S8kzHt7d4yFALLKuk9J7oxqqW4sy91dliXOy
3XbeRVFD/L1PKjIBl4/mCbWupqeDezOHaL5IXvCLrB+wDmG2jlyaJWAq+W9DNaltLk0wxtJ0v+/O
YT6iNaCYybPZWzezyveacM8Na8Y18TT/8tT1qAmr4R68VPuQ1fIiIrR/pRSVhP3KDehlaBUdDbzs
2t8Pbkol0VLpXEuZRqzRhI3eHISr3q3QyPgFbsbzKlQp04zuC7CnhNSWJ4xm1EVqmxLrOSBc9RrO
4TZQyGqXV7DVBUj+aYxEe1/sSCzi1UncfErc+S12sGZG6VXNp9tnqf0p64/ssdRGHgLBUfMQxtwB
vU7ga+/pFYk1mY9sIMW+ECtGdAp0EbM7ZMzWTQB4ZsljQN3/ZCkmm0+zo+Dgh/4IsDi7JapMefAg
x/qc/G8xevPoQ9bQ4FdggNT1hm8l/OVXvHFtybowZpB6mWNy40Bo+jRQ0gJikI7J4WA7hvpxYXrj
fcxEqVtcl49TPCslTvkf74hDIzYkqX+Mh9sYWzc5sNo4euB/0srd7CVvZYjq8XwHSQNGzKHbkexU
T1e8Tl2Iuir+nxdYLLqX+bDUSmDrg6vNiswjU4QtagSZ5f+FTr3VhfeGl9UEVJc03pzvgwRAONuU
4lTbplNNlN1y75olxjMjkSiy5PRpXACIKBfXiD084RXUwD4r/sNbj7kxOakBPYoAjiC0b/3VU4Vx
txeSZl8CmopMLW1SotgSlJO5v/EaiefL1P0QqMfKL0J7/NW/wSD0u+3eS1zSkTqI5FNSUL2KTPJN
Bscait/JS9knnJFf3SwD0JbSKcBLs+80i20Bg2TEi6VvfsGAwEpVlZlOAo2RbGqCsG3vDoz3KdKe
KO6NtPcIjEJG8EQ7eZxuCHLObyGayDs1Boj0XQCAZlrpG+MOiBXXTpNr1L1NJZY/QsxgZ4daZKWP
jI8cDjHjPkH/YahHKBqCkdyW+ZIjt9oWYB49mYT2pad45nrerArvQCQRLAEviyR6Jsy9MqojV3iE
XGKnkux6QY978z2lQadenmkUrPUKPBVjjmKnMMc4ykTuoQ9ahDqnNG6hi8ovqct/drD02nwZJuPx
ljPI/ll8nuK3yj8ZTWBLXL0RWffQh0rj5dGaPz1BJX0NBf34C1I3W2ikv89UHt+XAnLBV1De2+9y
unnmMPWra+tlH0wJtxxZUs/Gk/Iivef793wwPdRdJAxR0he785131HKWROvuiegxe0b9YfOxb8R4
w3XmF8Z6vmXXQqyuOCfdSDGFHiwT5s1KK9pVgy1lmRCoTM20cJw05f4KfIpqJj6c9JLQCUAoaTXK
8EU2IYis6rgJ4Ya9RAslHD6SU650obhI//siQjTvHVXSX1pso1oNEGa7q3IyBkMXr/Nhhs7JEvgP
qICYOctOKEhVhUzhBbT5WTFVvL3EJrqdNCApDQ3GRfhbiglSrao4I9behgrypHBm1BZVMpqvBqZb
a+G2xZ3+LgBSaWO8DJrkR7SSsygiDpQDaoSN7EvdQeYixKCrMLVQVaoBMUoKqexIWj8ACmwAyMZL
I3kZEfNUkjldopYT6d9CfHBPruUktqhI1n/DPTs998edjb6IlrZgAMBysO0GGsGhDRDhLHacQE5z
wyQgDw8FUOZWDKFsxAtIyeDxw2GtoXTnXXxKA9FUdA91tuqTTmKL3BHakLRCZkAyN/au3gzZmAlG
SbnS8K5+zzYgrFdUC7s2r9bZequ1RGB0bLrxeN9Xkb0b20KsL9iO/efeSxQZ7B95ZsBMK55rch+z
Sigaa017cYV4+UzIzMFjViaGw25EQ9sh60CqFLPRVdfv/BRx023hfme3i5csYPHPfvZzRptPqgOu
zf3IA2BzWIBcyLkqLWBmcRtWrMTh5OcKxISnK8Xq1x0IBxlgimsk6MMH8Dm33yVSQn6CpCzEKPhX
1FBl8e6UHyCNY9UQPEaIk3XwH4rVv4a0PLNN/1yT+Kn5kQl4n1lOXpkWdOCnt61lvWUFXdo8e72s
H1zHRmf6s3Tz0AbXk1qiyztK+QaQjX/ZAoLn1WFadU/fPeE/b4URq6JWjk2sCGRyWvLRLpbL8iys
S0hTCY7q/i8TxbDWCPnviWw9Bgk7KQzE5c3RwKT5dQl7xxYcOypKM8y55uVWYGLCpszpE8rImHhE
/N+5p3TtRH5N6cgiWo+D2TkhZyrWk4y8WrPkYr/Rd0O3f5fvHGtaAxzO196/WLQTi14MZ4fV8SSy
S4MTamFDSERIbClNEP5quDyonsKGZK4AKUXtwjP3eHkawLjdxx/duWDFcvaKFvt7yOWdasPwzt7a
on3sbOwnVc0syTm9FHDDGrJDNHeImfjyiWjbwSP188pbmDXrUqs0QkZoDK5tlRyskL83Ne/Rf+sT
EmnnbERWrIT7AN5rnao+gkWq0YiUxfcnidRE99KFK8EpYgW8z3ihxTIdT4Jgyd3RLtO9oOW+hlsm
vbDb+BEFA5GqZPcvRBhQ08R2bG6sHKcSa07Iy8/fvkzkmBgV9Vs7P0HSvYMtUQ1ybGPcaz1vHvOa
AcO0HaQluVhySSro/Qe/TjxWJmVdwYn17ucjxDwtHP+TLZ22VupekbeDv8liAVQ0mGJI4PdNKoLN
4+51K20hrEWM2M0aLNn4CpNHPjxxcSsjCyOQu55ZkSswaRomSYna3oPJiBtpb2DzPwbTNVYnNyld
K6kdxgp44y/3Msz9ee7EqcQ66pqEjW0lwH3rHvkxdRwEp6bL6Ra6/bORPLdEo3X719AJ3A8JzqUG
YXN9tgnDBkMVTuRmFyqQK1vwW/y6CvtEuzCO3iP6TdJt40N3gtF0ZthBLJpgTN4mDjOMvoez0u80
c9VPPTSE1YnnJnJzdXc6GweCPyfCjHAztM3q4ZOx20k9eeS54ACo4W+OpiAV2lX6IaYRSjQbw0nt
Lz+axNyltKfi0LNo3LvZsdaKB8XzIe7cLV9ttZT0Fc0EfRZP4vaoy0k+Gboeb+J2cy74XuCwWvDB
r7KNLmt8MKKyIv2gbF/cluTgjvyE1Zmf/Y85x+ZCD7snfe2053uSblPnEWj1HSG96xXImQF16cbn
WzR57vjw+fmlPGGpe6DADI6BgsiaFIyzaftZa90wH6mlpk9GgVg4gu7SmHTVf4OyOVWho7hfF6BT
bKCIR9Zp5TcyC1TV1PBTXLoXoM+AomgGBmffmMvc34HnJmcanKZ71O8AhvqIk+b4SUSgEP8yafsH
zCiz7CCauDZqxHu+0QggrDuFzcgrQVpcS08v88FS+uyweWcpNJ1DFgh2811AJCHeuqnSYIpuZG0W
4VLc8DgCAM8KP6hqwBv1rvF/G3BLxmF0k0oztqFjjgslcms9VrUR0GCQLlWX9016mpr8gn2C33xl
IR5MRm9yb2uCA/57lwR519jTeQG/pgMkTpAaalXGxVN2d6+vorW5rBEh4KJpajbTsUEdxKWSyjir
Ja0QFiNLRDNYlv6pehXSLu2B8pAJsW4m+/nSJKhWaMorzrE+2FaJlUsSrFXKgBbVA3AX22xcAH5d
dlmIuPVsobZ3x2Gl07JBRePMpovzhq2eFY43zp9fem67I3sog7YSi3Vz19J5A5YljM52PRtAPRVd
ykeas2IwdXGhk1fIB154H8RvCW4dTDCAq65EoV3B/Yr/LLnwST8nqX3N3tsDpakefq4hoHt0XDMr
DbL6Aq446vVdD/pC6niU2tacK8RFi/mR99srvTfzp0Pa+eUIcPw+WdYSRDpk9RcHYBW7JMfXB33y
FQrGHw0sY1nZx535ZQZJW/xV7dNwEDUQwcysF22BPioTSZNmkFtKWg2MKSlQ5p/ydx2KQryWiW8U
P8zvnoZ+Wo9v7srXxS79ifeaOhlKR3qi54E9uMa5Xg8R14VxdMnG7cmKwpnIVch1yqIsEycdSIlV
cy1Pfcni2Qhicsn7ZEX2vbaBraYbUHpSGr/2QyX/YEUFNKS/TxosW9FEgVx2B22+bJDUVnNHyUYl
BQdMHFHlg/MX52ObZakE6vbBeCSdc6p9VyS1+byVMVhuTUwxGJuH73cESiZkKoiVy+dXtfL3LBg2
qN3pWsqI9FGmw67dxBjFs+NflGhkwZfb5IMxOwbLCZDYfklmN27gDpfltHEkwQnkM8kSrg9m8Xh5
yA9COt2n2YyeTYs8XIA87U021mQzOAqOWQfDn7U3ckC4B/IM8cq57AR7C+lhIlSNx3ySDi3S1uWx
/OZL4Ttt3HFPWTYcKVpZGuG3KibRZhEjQDA3JnXlugKZXJSZKwmWXGeINTsaxZbqMpRnqQaiBdwN
vGbaoA6HVHZ0w5RLRGAYw6Rm2vH5QNu4aETpL1q9p+IxV4mS1Ymx+vnWmp71bUuhm3LMXEiCnVB+
qH/6x4vo2JZpT/b+CjN1TsqXMXH01PWB2OdqyXVtPmG3gl128ZfnsX1nVhXbIUQruF/JAMTKDv+N
a/nAxj+5iGfQ7XQmQDrkcnwrQPSpxpwSGK/eOgj9311QrXDdmXCVQqqaX9hdMVnuxvoRPv+4Izde
9/Xc0DQWL6I6lsDBqmItxkVc8rc2SnTE/+BcxE6vDmX+4FKzq3AbyJK1cEcWfmPNiSaCaLoLbv0l
CyyA2eXleOyLh4hZb0+mAu3dYzxi/fFkvwtG6uIFe6nVvu+5R5iK2yEYqMANSLTzNhGm6OL1uVNh
PHwLrWpkawrd0ObmWO443ti8dhjavHWVItvOxj0y9dFSawDK9tWfe4+s5bak0htv8ewSSHor4Q71
OcBNItco2/Q9WeMCWbu46ZPKLvrkoD3rGU1NI5QwDunLohdvjO+BpcE1dMZVC2ZJ+MQ8F9yHvcXa
DjSxc4djEATzyfR8qapvswHhKDkGHTHztmHHauqmvGqFkA+6NRXZAHyCCHdxkuDMjx1cI+SMrdsO
UVAQxm0FZI0NICP6Zb1LDM/3vjhBvrM/WdfqJrRbHBHWkeU6fMhPj/cYUUdvQZvqc4OMcMzTvhA2
zNALPC+iBaz7R2+ZZ4U6qkRyGxQCOqSBDeKCsIxGlgnm8MBCUqspoEUSuF9cMCUzum+02aVvO/P7
LTou3SGyo5PUXhBFijZ/YGfRL4Qt4dMXSTtLliQm/lze4/rwBMKIWFRFxQF1pMYY7l3ar8UZ2O5R
hWokjljeqI+MMQTu8aETk/5PWv/uXLPEJm8FG7K6euNAu9Z5imXIeTzPmD2M0jb4mOh5zXN1GxMk
AEKRpO5s9+c8omCrYJz6xO/eQw6PXyqy9r1FssK0NeNYPEe2hEQ27UM2c69VLJsugMjPQ5eQN8B1
uEAoEP7/wT4t1FM+gtLbbDBCWT+DmdRe3EZhM5wU2ND3Lni8gCzW3SwR9l+laoWkdPtz74SSaP4d
zAuPkWkfJr8r6t8vXRUJNwFWskjVIPWATmBS/o4dMeXilcLKPQ4fGtm75jYTU+eQ52M/diRuTCDQ
ZHeD+3kaGPKZD0zwSDt5DoCGwnvR+kvqGucYCU1ZccX5Y07Plfulx6GAA6oMIjqH/5rpeueHSB5x
g99MXKjKtzi4L9G4rM/LBq0kP92LsY/IVOYihNXqpwo+pVYTjx9h/7aFgm158iwN3y6ixF5Cz1Tz
RUPqdn70UY0yw0EGFJk2kbn/3nJqYbwE2Uy2LPK8MkxKU213NnU8NCmsH3BNe9U4xi1KeWAPcVJ5
ePoSRwrruUMj28oow8E4TdbBVsvtGKMvi0J39ZFnbajM0CSsf91PwIIjH7oNs9SDEplxdfKOjJtK
evDJslaOkAjXhxR0HqtrA10ODtw989sHTqZkhB6BsvIksmh3jpLE5Hf7Ky/V2qOoF9cL0ilyak3g
G+pJIQ/Riq5KPCdWNDc/6LhPkKZDmGMIV2w7YoEiIEvjrzyFIScSc2GaL7hC/0XsCAY0LyQ1X+VK
qOF8KJiAloBwC6t9yYdEFoYDCqui9QS+n8zjWm2iqbLt6mhRsPumotrFXt4nSGMF/FVz6QZvjt02
HHOzCzGfKcrASlPV8FHy9zBjDTfnJ8KY/8ek+b6YcqsT915jZnj/NtO0XwGwNAfy/eoEorCWkPSa
shypLcY0QTvYDkK49MkRO1rPL99Z6kvV7AzzI5cjQvuC1cgnNVOiJaU40AGtA5YSZdrr5kIuDBgG
D48T7+1el28PBKwsBVQkU6fRfGu9x/7fPvGITIMzYh6DVvnsOvvewr4YgjS4hfdZmyw9dGTqNnNg
/IKcZjeYpJEbY69Yw+otZWnk7YS0X9ghLzjcD5hpBYmzMJYNYXQ8an3VE9OMdafa6lAughWLep0r
EfLg7xNaUy45k8uWlm0xsUW6vRmw9RAA1Ymq5eyu38U4GfUDIHnmdD8ji59vbg4JwANIGmfMuayD
JkFTJCor4q8erUy0v3r0eDEWMvPMTqdmJE8lfOtakQ9BnO6GLDKW6R6zfEYrVAey3g4wPxjKffZ+
cIkJcEl1Pv91jmJPulrvQsyJkXR/lZTyi8ceHhMvJcmGGuofVl3NLRpjBvMYP9dIL82QEuY/XGnS
Jms5iLU+V7YL3xpskCjlrkOdk15XAIXU2rUR+0bwYyC8ttOtVwksKQZOvwZKk7o5mh84AwwbAtQN
TiOgCOACF4oBMiE0PEEf0sPnTYXfn1EGgBUxQOg4bOF01No1OiiP471lalYEpFLUiCh6V7BkMu9I
I8tYVWW4kRHINz3n6Xo7X4d9XKQcv5EACrm0ZA8k0yPtDqY6+oHevM5p35oVEQB1RxTHF1KGuYLo
O99rbH2Xw3xtIHmM94VzR5jXJ6yw5q7bXw2K3iTVyd0+MNAvrLr73AnAN/nMVa9OTmxfnCuqcPq3
SmZdVuS4RazaaJ9gXo1Tinw+MW7vHPpput3FxZW0EQ3JnysngZK/WfRndfHpG9g4P4SfZCl6QWP+
uFmVuibpV8rXyRgEF/1HSSQPKkTWxhExZk9BXbH2oYD3aeubEZtmnj6glKzgtSIDwnMFPsYCJ20L
OpVOLUEmeSgc7oyUprNdntSPwdxW8iRfKkZowiaPacs8oGpblDJC2RTfORlGJlxJ7CiASNzFuSwG
es8jesMIG51JDtxF2crXWuIzDiCv8nI9r7RGcOlL6AtgTfGvYJLhHJiF1ArmWhOuN9w9UsS+i5Ne
vS1unrBqEHLkORcvvA87mXI+7+z+HDE2CqzjjnTuTz7dEvN2Bpc0CyjPoH5PjcR8P6eMwBRLozhH
QQtzjpx/Jn7jvpAi0YSSA83nAqMjMI/8V0jlO/fCqJLJ9hoknXIN/KYcNpDh3g9okCnYXeZ0ukZ8
2OxhKjd2ezGgvpLQ68BVIBLC3MKp6Tm7sHNdYMoXO/H3I01XtL4kSYjIS8VhVXi+E2xJJE0ehohW
Kq/ops7TpZn78TI0wyupFNZa6m0IPP+S55BsausXF4DZnEvaE/ku08+64n5mqwv9EFLRGRK1fxKr
1Yu4nwZIqQMnEqdNsWlxZDkwFNUotVuwHcQ7ea2LZ+5GEUjRSp9CLMXnp197vSL26xV5sFv/NTJd
3Jvhx7KHC8AYvVVOjPhjvT027QVOMyjeK6VpZtLP3B0psQX5CJrEzQQ1XvyaP+ajDCZ8gPtuOF9L
niWgxA5bd48dhIXuXNrJ5Ayb9TNGept9GPtMAnw850WZA1kSLtccX0DsnkNH9d6T3V3KxIFk8VLJ
vfKbmpCfm2XGwrh98m836SEUnLdDxon/uEnHGP9UG9fUH4VLu3ez8hp7Pk8qC5CKjj4Xey1a237D
kfQU4/DW9ZO2BKCe1cwmER7/REMdh1J4si02ypor/z0Wk0+iGHl8dkkGrn85MY+7MJTZw5FrfDdL
wEjFQSAFwvgOOxtPZ+ZnxalfV1FwBlyRtulfA39fNcmF6AaMaVLgDchW918xI6O++5YBHNW3l1Gy
wu/7m1F7T0eVucNwfjdntP74PlsDiqRgvCUQMpBNoZK1qFDcUARR+63p+K2woBpVkNvnSH9kpiPm
d4Jg1eOTXkYyf51ppfIqoda1BO8oEcsRvNKV21FS/BbiNW6FNB66K2+zPR8SaCF+r9vxfOx3KApR
d43qHPtedLHJSDYHf+NqfBEk4o2rqhRIUh0H2khlz4Fya0Sf9JHRaEx8MOG0AosUb2qbacHbx5YL
BmeCSYXSQ2THNibwxlxHbr4W9mxr5yCdt8BDW20fdYNc+WmoPw+5/B9qCCRtLDJ/bM6+m7/MzRUV
vDjLtgvz//vdC3+cmFnrV6UpRZgWdYt1kRHB3BWVyb/f52SxSNmZy2Y/8U6vDrsYMAD5CBrwPomt
7CqkkHIqaLab8DmyWCwnmkR2oDaaTRJZdGMbVzc1gCJeXBwSwkdxIrPrs/+8GfSnmC7gggLxW7Vx
qpgwHRkhxLKrYWPkl3A32nQLT+Cuh+m/Leup29GpPlQ35Ihho8FxF9zEp9GPZrJYc6vGK5n/oNQT
y3DkOAsxuSSICpr9qLM3BSPWGCLpx9u9/QCs5BciIydj1j7v1X3HZ7hUJknEZ1txYocfi/nPV78h
r/FBJvPV6F5I8kWvyg6M90WAUU0Tlpl0C6nKevCxtXRz6p+7IZQrWGS0ay2yBP0mlQtoUBd7I2qW
v9IaT/845DG3LPmcaTwNDlr4cwfqLYOwb/nrbH9sD0UrMrEwaFSGWyXmUjhI5FA/Xu8qWAG1PjdO
Tp7SpYJoRkEjaO8GWoJNdxC3fnTDGou2VT3P8ZhOnJtsyfz2dvNqNRYFSJStTOKGUMlzrekIxR+Q
dAN/L2UZB/1gR5Knb4sXSXuACsJn7dde4kFa9VNFPO2tYinVvFSIIjjCcP1TgeKnOM2fX4lPvbaQ
gHOVKnextCW604RGhZt1oso8NxMNKnnnwvj556ggDwPjJS4ydwWDYRX0mf7FISUZjiIhT157xJo1
zCh3ugNMbCMlNAO7Xb1t0NaqpzOmEfahtahBU6Cj5pfqfoKTGngoLVwWrqMYAaNXQM0D9M/4dRD+
LClx9UZXmUN1cuZ6xlqBi5cLoKDIuggdrv6xG94Ey3kRqm4jmTJ56d6K76B6FwgL4ffxN36PDASF
myfco4JZ4mFTViGkY5g8FnsfoZeCWdSiaGpS2ic0OCaUJBf65dXRg1CM/Y5xwkEp/sCFTNfU2tfW
fi4XyEByVY2LFBcaesstQqVOVN/9NPm/xbsjsg8YNIu+Ss9xJWoow7I/NjIBUv08A+4U+8r8vPl8
Ly4sV+umT8dDZMgxr4ivXafQ21HNRp7GsVkdby1CDXOSOsqhTgi18KRy3FPQtodfC9lQAlfO1aWd
OVGWFIrI2OApEum+fgJaQqR0lr+NqdhuqIWXZmOzPSSof9IXIrFjz1csWZe9JlFe1HdFGqHDG+Gv
o1gD/BzzgLMICDKGATxHRHewmlsyMWNIQJ9B3g2dh2wSoRyAJaONob2TyiPE5U4x3OmfJBOTjlXU
MDV12vfv2OV5LNrEHw1UiXXEPRHzI0ZqC0oFrDs1sX1Zg6+XHfkT94eZpgjVRh8vvVCP9uba7Xgm
5lPeu3gxrPtxLKLqAxvanj5OeSBHO1kKWwcm32dl6PlLquho4rfWsa54BB1SS3iBXtgfSf/2WKj1
saZsgf51BiXeuBhzZDreRAy55fM7SHMYCbGVls+hCTsGD7Ryo35e5dlJB4XqhsaZUCQ/05Zrx3y8
H3bixmiezYPcG2jkKJF0woll0MykXZMcNGJyioWzTlzsCxHKCgPWWZCDv08tnf/trOftqAE7iRAe
IsszM4jSD5wfMSXRVixTonuEfI7O2G5lrI0Cr9hdIW6jpn3jSxqFd6ph+UEKr7Va+g/48WJw7LUN
J9zzfiDr0KMAlfIhHapfbyzJtF4e9S8HlqM41PU76863dms69HSGeaOdXSg4eKX9mw0b+qExTJcc
pZQKPXvKaD19EosQD/79JCMAJqnhllkn0VZOgypGusLL7J0SP7mJIGwz7aPqAlFVotVotFTTvj4d
QAwuoPFa+60O9Zc5a7peDEo2XyGqMNuqUx50CXHir9aKkBwSruKC9DHAC+F4WkMyZM4BtwxQ3jDX
u2EppY3HSVFVJ9kWMmFsgexOreO53LJ6cL+dweKWbOQ6PaLDP0x2xexDbC8xRiTnZIC3bkozb+sG
X20dEXO4JMx82u4sYiA9f7PqkVag6rGQdSPXrArZL4q+9zXXYpGWBYTAU9txXV1UPG9FXEmYoGqQ
XXU/n5N/vccczk65XOXG8nMhBRq1Vv9Xj39lNIFBzs/+CULQ0o490g/xC8zpMyEnv6cS1OJ6i/WW
i9ZBOVfNv3sVHnIN9x4ZGrDnGg2yyArf7GcVDaoIFGDlDO0ATYn7/8Y9lGwzt0kW4s7xfeDVXfH9
dDfJPIjtMn/ps6voKpAa1finklcanlxFEWF+jKBYmLEqH8UGNQfwgiGjDN4KL4HCWMUhWPlxSoQI
/T3mJtilJmgheiEhd0xfFTF8xgFs4zHw+ZdJGOJlDefW6LXQPP7ymeMY7gwfCSRDZgmP08FRtdlk
uQwx7tnoyQPYyfShFCj660hPnotcH6qOxzMgFGBtTcaGwiC/ziMpZ9SYBoa61BJUenJz4JH3YaYv
EfTNkRXatlJAX5bJmL1YAEb6UWBFyluS0YHywp2cJJe8o6Sq85eJrYdCojeelXYDJN6EZ2IvFdPR
8EUQK6rXN6Cj96snvKLS8EAkj2cAnj0VbyAw+fjJnmBZw8XvKOvy2UqYT1Q4/5miQ6IZkhpDCmdz
jbz6W+rOay2hH8z9AVKGsDrI/leoritYz87ZK1n60cBV3Kg6/bD8BVqp7k/JVbscRajFxFm2zVAU
4B+J850mcE5T+ZXlmeAtoVLL+ZjyeJc3oeizlkIas/NFE9k9unCUkO6qvRwZV2iZakHX5UZLFTVf
fpnpxddw1T+getB+Y34qr6MpK9rLHdmM7/yVmrlY5pHJtC6U3xmabhHgrZPAHHj5y0LluNrlzR3+
u1UKeWIdy9IVSB0/YXewBhMqkDtR0x8hN3GJDeYQSOu6q+eiRAk//BrFo7A0tUBnl5HtF137SSTN
sCe0TLbJKQ2CWtzdA0iDaNMRMv8MgVaYAZ7yft5dPQ1xg93VbN6cxdPVm8DJ73DuSAM2je8EarIG
xiVt5Ei7HhHghmrgLCweogpw5yNECzy1KG1Oc5G7BK/y6OBi8cJdt6Aib7iMkSk31sGD4gbiCSxc
jskerG4YWpKfcetJDNk999Zy81u2M3SxBptutBKccEfFGxfvKsCRHGGI+C+zIfyp4CAVjmQepzdK
lNvSY1JOgfqHxUOaa+HT82i24R2gdxWKclhN1Debq4XbH5vOgf2+wWeR9K2gVvvJn3N+9DhVc0In
VIAHfr3AyZVcleBUTbJxnsjvJfdiA3EhLA323Ch5oDJEMCeQF8+iOFGFC+nJ+53MB2FfKcEZakyM
pSFcebtl0MxCEa3wrtQ28SNpmmHuXAqC+lDBh9g6hO3bF78wSgmpts2Q/Y6hN0bDfOOx3xMXsO5i
3I7YbWO+toDQ4wEpCmF2IEaVb8HhiWUkRh5elO8aTIblGBlsjxIEfjSYfq+d7XaZ/lROdND5vOkx
nf7cbDCIs67UDc6Ah17nmA/XY/ukY3//wMwSfCNe2l9zgMAvat2W2vBLRHNrsqiEG61StOjpt9c7
3QzEmHLt29rAVJ1Tbb62+7sO0zRN8ZfU88Dx3dHWkvdIhM+UE2vc22Fa6Mr0gGoYXWRdL+DUFVGU
sNGZ44fkmNpRorxzbSaR+Q2HHJxUkyTaSVHdEKjMrVWNJuwaLk3Z9vcZdczOAG6h1DgTg6iYzLCg
z49EnI6Sa2K1jDWZprz9ah141ZlKX8nMC+5c21a09rCXGDRL2bDs1tse94H+qm8vkajb8TBBmd6n
pR7EeOiHVy+5sXsLuLxr/b/87wmgrhzBM1HYvHSQjTaqbQBaTdRURjaTvdxoDLWA/YZqWsBhMgPS
JhG4u3dbS403eccnlChDQ/p9EO3uzH4ZbmCRRrtgtxNAncmwpM5J5mQcr14lNMrJ8gjaFGqCWt6L
anFdG1wb3PDbTi6AGGV/sSwZMwfG+IKSytGqjRu6FSXBQMK7mZ6Q6lsy+/uCeETh4ibTbN+03qRw
nklQpcbk1dDsRw9nT2nTRwM48mcbW6/mkD4pwz4+8d57qfZX8nnS2ZjwrTRZLhyI2UQHX0Th5Sze
M7PXaxwS631ZDCX7aW9ofvTNVcc2n4TBSKieuknOaaZiF8OJiKPaXAoEZGNe+OrzWxl3+JZDBuuO
yAl3kfrQrC4NH3SIfJJtgOIn54E1u435jbCitZKD5ZW6rc9orjPJlfJr6lKrMjqSQQ3IdNptAcE9
LHx4S3vV6XVFaRYveLWQ8LKATI3XVoUYkYVQWMsWGJP+YYeyDx1lG+2Mh6+3ZpgEOTcIw5AiDYlF
82U/3ISBQUXGyULvPdSQkOqsBQS6+xAG+4KQJtV+K72ncmii17OvyMMl3TQRazQwZG9Qmcu+o6Ek
Vb/l8bk+LKc+PR3g1WpeAP0IBq0RKlQ//aYbVXm0ypJACI+BwNsoSoaOuBxy0TjVq8C2vTnp5WD9
OMuzT3k3BJCmWMm/FGxgmEy4dD8LXWyqdALm6O5o/T4FifoSbIajpRdwOwby2dcQ15Ifmjezh0zg
QvZfR2ZAVBA0CEX6rOAxf1GFEmY+JDD0sxb4YDGtkFUTKlpCFPf+8rpehASODPSJdAavM6NzkF/Z
RClyBvIjfvLsHU6F+CQcHOUWAyhVxJ5WAfyhjoYvVFQLaMwcRoF4Prhhu3lMQWcqAMs8EIbOAHba
Eyv6UwPgfP2M+1ULC1XCsOhPs/0SY20Nd9Kzgwy7QBO+PBnNEpsBasm4SpBack9VqoYYlRl99UdF
5/KS3jLeElQNhAOu0k5hVvey6P8/esImyLlCBCGSUY3tyBhkXO3ZWs6Dhpy4AE03zeFmqV1kh5NC
q+O6h+CkxD+ty3Z2WchPNFYkpC50JSeCrl72daQNxSNFdQYki24OFhjn+CQTuwQPE8x7E9WJdu+9
3YaEr7S5jHW7kj/dTzRBVjbYIbsaZ3ZDEdquWCb3P1EWV4+mO6TMgPTdhaHIkgCixMx23E5pFgHs
oe5T5xQ/K/Q4LFZTRLItHRgHHtACvas05Vz4R23YXAfvrZmPxncVh/uAY79Ex7eMac68Id44lagm
x6M6RA7qjXH60EdLDAo/mOoQG4qxzBUEX4z8mS9o4l0DaNuKisTmjomnd0/9IlFkbommU7k+7NS+
pGaHZzgF8QVSCbopyuRN6mq+RPCgSyq4PTFiwz5gHeGI9TbfUjLlzJWDr8p8tJPC+pdHou5EStgo
tvCs32tZiLNOTntkmktxgsJ8WsSmohuEzSObaFPNFSzvtcWXVs9ivjyZv/0Ox+T0F6QfubeZZAAA
t5Hzv9vMvGgjJIfLOiFlA9rUaPOvGtFwg5uzvNMCvrsRqwyzAuu8Ar0yax59rd8LbretQtDYf5tk
hNWT88XlowgughOSO863BOKlpdYNZwO7J52Gwl9uEFeJI3P0ctp6wjRVbGZBsiKLBo3pjlezI5//
f0Q7YOdVIdt2yoqmlgFFrqVEf3jyL302LWKU657yjRyzcuchP9LMac21JS8rynccWuXa46u102+v
kJGQ40lYcuwEm8mWQGod9CCgteeckFrM88HZLSiOCyFjX3Srz95Sey7jWF5HIuLvcDTP+r3klZov
xZGwyFFxA2uiFAVSgA3JgkXlJb0MrxkQTTbyVL424/iU/1CAZVaVlOs78NhWw+DVe+hBoG46TbhH
QgGB0Z7F8b65nVBtEv0WAwU9voV4ZBqZJTv9rs0mFQ3TTm+wJ5RHYDhieXVKgVht+FIFFZRndmPM
ZVFZU7rh2GbM5uKojhEmL9YWqaRl80owguB1En/jK+yjY1APyOK+ai8vb8RQMvPGzCNyECLzljNZ
UiEBmWdLiz/AlvdwprUOSw1DBGpONh9h7cNGYimboTpyc4Cc8avl8TQkSZPA7LLYA/isOmfbj5Fo
R8oPqwmPwfoXkecIZagSXJQYsj0R/n6J8uttKYqDoCJHXzQCEmMQ2VOJpTXBVwyDLzz5Wy6QWFGt
2vVn6ahdfqVACwMJ+wSjQ5nEx1ZWzrTBtZERZhEkDGsNAS6q4BPS7YGHoBmQyYddOrzYSnnI+t2e
baTl/5AteezAaHKBmDFamN1+OPEGqxahBmM9W1C7+W2tje+gvdfsEVhrU/EiFf6w91a9r+mVK37W
JB2Vp39jjODz/RL9fm93pH8p+ovyYAdqPvXRMNM13gAx/gxRBl6JdSjxmisfXvFfGkAFgYF9wC3G
MjiS4jB7CWNQsWVp74J7v7ug+ll26GcpWuhVgacLmgnfZWQM3orODywUnwZiuBWdcz+i/GHg8fvv
eGiOHU2wXkBt45+dbsk5ArFZv5wWhIuk2PHM8QUjV/NiwOdNzNoNgMHA5IQVg419QHx7ZAp3faOa
2Fu1pfm0VX74V0vwQ5hpxJNZ2WhcthMdTwKIjQxc6wGiVwtwitwSSkbhSfpPhxNyQga1IHbh481t
q5HxlMY8KwJDfb6Tvj4khN9u6pozYDlC6hYToG3035iwpWeiZssQSVtZZiIjEi/BeSzdhCEo8U4s
q4sdCKQVNM+RP28L2kpTduM761erysKEHAVhw4aZbiIPVStNmcwmZvvRCTn8jIgaPSqF/V7hVALO
leWD2wJSNZJAFLaRArJu47Xr622+u2+DztdcFLNh3Hm2dNRqInjKiY/UZhP7uPKKVGagLqay+JVx
AHUK3cAhfxjwKzlsQKOjbO3PCLH2Tvke95AjFkcmggTDcXTHON9ILIS6cWp5sbFxbQocQqBvTL3O
KPP+PutUqOzuPOCqf3i9mGXTBB2IZ2+LdU9GM2RPsETeTf1oeSkVUvNs97PsiajpcjZLiw0IOK5b
8k+iYVqY9oRm4wBSP+YnixrQ0TFEER7KnDidOApeaGweZ7tkuopkvNrLrjsX8VJUTsV/wf0g9F6h
v54THTUalHwPp/K+hYQHdjtDpFOuugC02vKGrREQm0Nj7XzA7B/USGbyoQtm1QzDjDntQRBapnhy
1Jrnb/V1oJRzIA6o6E4NF7Q+mdCXUPFMNaxys11KpaBfbcBjc1PzphzdT1q1VoB+533M+cDIi6bL
9he1NTdid0luo08fdy1OOw8agk2+77XPjdhurPZhjNIs1H7/A/NbjPDQFWg2ZFFEdoBlJAKQXZ+W
fuLnrCiep82odGZ+2QAaQL0rhy/Rv/Lv3pQiq9N7OSDodObbE3paFNTHKaIaXk0a963cwJwXaN7f
zAYY1aKFjcNu/8JDyVCrXWvcCUQFN7si9wzGW1OpPyL/GA0hhDY+d7JX7rTtvzAdWqsBmEeQSPdM
RRKm4scbYtzY1vAfSLoftlNzsYvOpORfCP63SKMHs/0v0vI1xe5glblQNvJ2pM0t4YH+CFRCDQl4
wNO9rXW8L3YOyCK5oP3q3gc3/uvhGkbqCt54YlqXOwzkwtKGD/3QYs4nvtyWRtX4D5UgViGeh0Bk
gQiTyvcAhIm/T221Qg0ONWgm8KAvWo5Ao9PCiLDegXwl5BACaOknVVQnE7xDKHYMXmokr1L+Dn7c
JkzURaO7cxX7hlIbVML8Kq+YIQVAcnnM5B42LLtw2DzjfbD5k1KR+tFxx7iFAzVieMrQqFx2FmaY
HFS/mLdRuJhK5U/AcvOV7mGDoBiw82YfH+LJYhdCwp4vKEb6J6OcGmqKL82jDdH9s2nlXk3bPvjn
7btDxRK1OSISe1eR6WVXJqq4I4s9z70M8rW7gculpwsq8EQBJD9hrHPUJ+UT/fBaWUm83VxakCGF
FUY5NHDVeEQ1eB89Can+RRG+mJN5B7UEOVQMdvnwJ6Xg1uLo4bG2TKzLbk92FlYQ7LbVq8F0Kp/E
NNnp+cI1O/r6NZmAwd97fnVP09pOv2dQGEvli4PEyG++dpP01P1kKcxzRCvAIlcoFxqDvLf1KgAz
ssH+5idXXzVrvQejml36XChq0S4dAotJMfHgjdEVuDNVfdXMBq8TtunERlhrdrCjlGt0GPGmW/mU
eR2BeE4qyDepywMPJ5F8P5xkUGFLOjgrQDX6Qe0bLJjybUcVCqBP6XhuYGS30luMWySNG3+iv5Ps
bkxgu0xYPMrULNc5VVO2hzp5u0rgBXEg792AfkbeJjZQliYsQ33WS+e2pYRuaOhOZWVvK0lsN5CT
KqBAU9FRoHVzSmU46pU6VBGq0fMhFFzzUSSRBlEDPZcLJz/nnCd1LKxpvdsRnq95H1BWO18ItBmz
goWLDmgWfOFB+mW32O45vKrOD6eWclXCEKQlpeUbdzWU8c3aiauqrtRN+yGLkt1URYqPRuNYQ53h
o3aJV8KQGxAQ6n+iWDWUuls8iYBSA9F4OFUS1A8qKWKdw7dx+RvxwR5lc+dAyu+ZSYWtfU+9yZE3
48c099TXbr6boxjDrGjt/hF9gj5xaeFSDgYaA/H9swMcdefgcPK2jbefhNMmBi8LISeh9RTo57s7
GApfnmK5cLekFLLOSGw83BGbbayVdx8t4lFR7KC33+wlim5takrwo3OnUieDu5HTW3enbTOLofDd
vxt0XrvYx7WZ4jtVKlvlnhdfvhil03lHnq8Z6Pp6j96berM4v+1nGJBRtaLpxiaNQm7++sstgiOa
tY7D35Ef/vHsCo/tRqSKBbDOREEzXXCVs0Pr4N0BVX3o/Nb7fRvsHXNf0lyQM6EWJijq3YAuzJs0
GVBLwI00oW+5BA7zEyHEa2GPvKieQGPE4EoTa46uoaTwW7CzvNL74741A0TljehFKPzIa/bH7VYl
ECmyWXeh6eRtCMoFQUqqZEfBeAmny8QSPVFKdv5Yp4FA0YwoVaihsP7eGmAH7oKGQbgtUOgTsOno
Sb6Ps3ymSnjtIahicPQGZd/nMS+4YrrgAaNBQyTdl0nqfx6yFBQwUvyqWay5gWQz0pRQAiJV7Jql
Ud/u9Y9ZF81j9Ffp4uAA6Q6KmVTrJuNjEDr0uR6S6+5UL7M7/sEIh+cVnwzobEopg/QGE1POkQ3c
TVGJSf3MRzyJJbPXOwjtGHCEd9NdUWLItQvxqO+j+oBE2xjW48DOGxKfMiJFoVd84stt+I/WAr2u
0K/XxgrESMZ3GjCc0UBwbjBTAbXqmRpR2bGgVFfIaVa+EZxL+60QdrvdsJdtGNE//1pBHDLUJ5Fl
Fb2Z+dxwiEBjYa14UTHy+9BC1j4zzQqlwkVydcaqEPIh6cnfcBbbfF+Ss9IMgTIBEWh6gFIv8xeZ
JHW2MfewUueZo8i/tFkJnpQs4aYpasJHHf/b12K81aQy54bKx46qFAvYpegzVAUN09fLbccDWIgM
4n4TmTUZFXKMihEfHdAv3EyMvttkP+nYC3fb0Lt3/4KIZGW2RnaofuXTww4Vbi+J6y7G5zxtrUS7
DGQELd8/C1bWPBVd5pEDn/YTyGBUVOXTGmMvkDO0MHG7H+hJVkWtOnLzX5TLFXbtEc8YQaZDc6ly
dsKZzHN86Qq8xhaNnDW1iCQsyj7MhywxFVVXYXx6cC5duLfvZu2GZOhN1HgNgxeZPXsr5kWAn1Cl
l+RnvBYEn4Bam4RsCw5fza4DkmuqAcdbToyzvKHpv5LIjobWxXFfKlNpFD+iSvcpp10SIGIU6idO
WMFIE7izQsN3YmDtrq/seqzE8lGERPPGMWbOm8BYTVKyHcl0Bky96xiCibaVJ3Oo+05hRC2QCW6s
jQI0sLoFCMhf+RehcYHY1mPnI2QwDjsuse3/AXODZv0JIf9BEGM3OuH+g9krhxZ7URrSaKoZEtoh
aRjEiCWjVFdNkW1yJxMZNWdUKqjQdfrQLVBYwba0pHIBZ1pgrxgxx4i4AVsnz6zzirqms1q2e4VQ
UHJ02yo/bMiQyXxMGocf3tyVolmWNrvwd6ZrnBi5ktW0RLsgaVVoQxOj2PE+Tmij99KaePlYd3Zg
NzYm5IqA7/p0F79++i12h8b+H0SoEhNvHouETzJmYk2eK9e2PCiv2C/rE/uqstmwNkS3RjKzIYqc
v3nYq1ZsJolxMPx1E+ouJANmhPnifWghox88Fo2/gKl9b2KvaZQ3lAsL3cTqR68SdoZmY+xClyk2
xP21+JGdfhrAJbb4VRxuEMV4/pA6Kvd7FGFss2aJ95IedN3xtVuUcGCEJamqZA5GgIecfEHA3FBe
dKHKneYj/+bX/uPp5n1HGZwY5Vlm78Va0uEeM2TmzS1bxvfGusP0e3WtqhlZ51BXrVBPl3tqpAVQ
smBqOjknCyCcoou56qCFLUGO7BnNtMGX7OQ4wMJ7BHRok6iSupKCiTXdCcP+UN6bw66wdi5QMAYa
tjfADBtLOk2KBlukkgzUO0jo8XXyOD5OGwVP50O1FIm9yjC/Abif8sPxVHumExItXrsu1n0iHq8G
p/HnkVSiby7jyOoZ7ICzziHQvw9hE4vXv++mSh8fI8epysO7kTEHW1aARVfPiUwwnbESkJWTbVDe
gUU7dOlgU+9FRFhPSFBrviRQHxsCptUGrw6pUtfSFDCpG3V4tN9VqL2+4eyQvT/rvuT+RRomSvmV
rRV8sUi0Ny/kmwtgKcELOLld3Kca9/Awpcpfu7DPn2zbzRW+MNl8U8M3rEv+xpyXfhsXT258S/EG
rcXHfppDVUJd0Bqs6rW+Y4N5JOgsPSQJvnQjvFTyPGKnW6ejv+OuYNWdyYY/r1d0LpwEm/5d4Tzq
geeBCcOQzjBVc5nAv4PbjaOna2077dgUN9picJXnPITedzvZX/PDH8XjIlz6Vckuso8/v9kOUh8F
GWcA1ywnxdxJmp7YPTiCSOHVdbqGx61Vgsy2QH4xGfbH8b24S4MPtM5PT6a+ZU3ciyIbjAtRq9u7
FKSnagHG9kK47Jk3TRwBBF2FCHdtUYqXf4Auc3gKLFIUz7HEmFtdIL1kIv/Nak691hcl2rB+D163
GJP6h5wObGV/pWh6oPIsUDTs0B+77bSRfvoZwv/pXnwtrY1Sj5o+29nEt2XSrOETazBcj6klU0tt
Dqwn5zy5xeEIcFXEWmHuqdPqWaFBCXsbKx4HNp7JzLPQn3E3W8pJpmyw9MzvCfVG+kuXOVpGfFxU
OGzZ4W55i5Eb1vu7YthQkKI+sKzuiHeTSS2/FidIsfXjP5gsqp0m1p1pFZFA57rQOsouvu4ormUA
rKDkBuYNFu2Hzzbze/Zlq+nxDc4Sh5qgZWK5n9V169rF5Qzb98eFBtfXjwiOP3h4QFfsR7SyB7X2
wE9IKiyflvtt6HHzilroRyqAWNxMluImKQgT3oARm5oxFaHcz8ccKLFcKUwwcytUrXWc9LkIC0Hi
fQjvEyOk15zIAT+w/4JCv8IxBwLCnryeHCp1wWOteHv/ckU6p8jF9nSjQLn1WI8/3N9VP1xvM5ll
iFrFnoYAwU7faoERQIyJKDvpZdf2kXf666j0op6VjpVuepaXPuqMkEgHJCghz/nSCdr9aX3KWUep
G4ICb5GCPqnPATV3x2/n9Jr+KaLGqzGE90P7zqahFa1bBzPb7mtW2zS5RmVebG3t70pHwvevNMBB
t079zcJYjWDz+3tUDqj26SOv2c85qvJwwOQBycCV3vrhjwuSXbeGwUHz+SmS/Qoh1gJwlFf6IaNf
oe71vDUwYEpQcFvFRNErZg3AadZBPhtS3G7Oh7og975NQkABkoPQNuXdFM8879p1wO/R8Tlf0FQf
UzD7Khy7jx51NqZr7FMM3RRFNWO4OjesLpLzubUDdNf9yhdLsEwEikJ3vsYfMsRBIjJR4894LVwj
XuFsXbvFxeOUQp69TV2DG15i3STEZb2R5CnQb2o5JhgzUNfF0axdtfIQuUG4QYGlO6ejzqeQMFbs
JgWKs7gYhAdxq83rhK1UILh3JujwufXCF5vpQFU+XMIWyEOH8Iawpnak83cz14oUW5zG/QsaMivH
3B1q0qHcyoLwt3fP2p+dzmGHmlL097bk9fWIxV2kLH9e8xoe+nemWOkFn1PbTLLaBrLy/j+c6f9A
adWbspN9vLV5/lGjyHxQ7mdYWuInWLuEJCXSzH9TwTyzWGBWyKLSSEC7JpUTz36lf9RWQxKx22OO
JYSEpNFqAapXeAZOJGq2KIgCUyNUYOd1ihdxBDmneMHIO60/jDrpDJ3V9JKLxaffoE9TnP+eSeIj
IUAU6PzdWElGlcR+ERSQX1ufPLNCUU4hlOsW1HD6z4bdH7XGc4a+BhgGC/CR5HKMQZ+rwdq83HlA
duDiN9jCUAvoXUDC1bLgiwqNtZ4KgktyMixvgQMP+yL7rq3nIFgOsITMulixw+G+NSSdhYh21xwS
9vaXqoUnjTf6fC/6lxnNPLsjDkWleqR9UKf/jVP8VlFGh2ymDV71xnjAQZrUBcsWJMaz1Db2zI6u
f0yrnJepAh4dT0fyLEwRypCzixN8Xnb7L/poKOqn45KlgeShobe9QzRh+DAQKoHPTbwSwEsekV53
Xs6XwkRh/hcEO4i2+zOMSWmtss9Kyo8ex3UQgQm5lrQhzf9l1cIhm0/0NPniqfe9oV/SwE0mwHxh
uxtKJMQ98gV7r7WbH3KBsdjvywf8No8zZQ6KAekh1oYclRhEiOeXi+tZ/VTbW8uKV1TR0wfTd324
Lgj3olCVw+BXAROWk4LPte6u89faILFGJXGUw8fJOKJO6Q+I70eOQtKe9UQ0Qo5LQF7nPCFnxU6m
rSHCgxUpsq1G0cd0CDC+g3/yhaWgZMjDci0duaYTZvtUYZnKyJOinPWZWdEb5acNu7Ay4r7t/p1K
QUvWVP9dlPgAJfUZGUuK8adZZFQtvfZAHIF+N7o1hH36Wr0jhAbW4wVfDnej7MQWzQmXKgHrtHeq
mVTTynLDjUmQi8eSLicj0MMbmQe/Y5TPuhvLG6Q+6i9wy/32hCmS6GRkvJbEwqGNW5ZjZxYc2XsX
CQYWj7QE//OUvIaWeFl777mI+EosZf4FvKN+wmpUjY6f4gmm2mNNIxTlGR9EdiRDL6F7ivXOqc4d
l4BGRR1ci80wT5mqSBXd7NuExi0RYVcS69/wqiE7p6x3aKkcgTdarrA0nh+IgXZz8zGJE2ZALR9K
aUd20OgLrXyNBu6Osj56eo0GppS+K81kQFqqtxuui304X6dWHiItBeKPvekw9QFyqY9pmQ/rOznB
t7KXJBm9S/8POg1RZMoEk5oBe9Dzoz80QMokF7igrBAij/lG6d6voIjM5vBsWVcX3FYnZ7YGlhQV
Zu1ol64hRRf+H8cZP7hVabAEf4kjhCV5f6jk1zPxa6noANRzmwfbndmggd6P8IXQV8nskYzT6hkJ
EpSElXHcVHzvujgMlu9fSFJu+rOXWCeYCRZWzCh8OuF1cHAP8aqjN3r1mXIX6TgkQpFLeKfrD83g
2kVrsetssj7SiBnaKnTjlP3wNKxLaIjHIqJBaWtOWS4LdqMV2e4U/SVTbJVWJoYO2OrZ1ixXpUuW
2q7nw7U9fwEHk615IKFN1B/EWMNFG8bGUvHpr9iIjBkpU3h2Mjv2o3A3w9fmPm3+BAzkTCnOrUVs
CMosyEwdMTmIxUN/rBymo/KfXYoEgN1Yajy1V4o6A9OjHYdkCCnN8+bUwB1TCn0+mkupFzRSeJ6W
kxo0DWCeYxv3oLjOXUT1aLhwOC8J3hGlwDwgFIaIFf8rvyY+8i7A970Jny6bu2qvjXo4idIn4nGy
Y14+fgrFXYViiE/2YsdfEekKpSPZsuhfk5BlAT1GnPfcsQ5qzIxz2GC4EynYO4z2vRbRYy/bGitB
CzZSY68u/6bPYr2foPWBHzVZ5W/6FJESWxwb5OTnUxq47G5NpNDLy8lZGwTVn5ej64bhUmxxgsjy
AM9xkNOGL+baxPJq8VhaDDtUUJL1avfMBur3MXElKaGXUTz3EndvASxDz0lazG7b5JzSaHxIKF7x
VMb678NQF0v9OXzsZc/XO30ewjAg1I99/sPrXNA+CxREVwstGKZ5eHvSqoFWiAtXSMxOR1AEHteq
kxZcN2YEMmr9o11aQNmRJ82XyoelzExsgJCCho1q9jWt61qGr1JtR5zo2mPsDVByTfWPfSKgO/PS
ylcxLbTGmRPpCn0JIwGECa2VmeU9MrHnjoH3dHUQvgBvd/ll82rfk8EeyI4lmh2yEgAlzDzuORO2
pmsko2+ShzUTFaOi83EuuqjETJnbyaFzYCT4RJhDCtKys7Ip3pRdJiIv9LR1HKwc6TJGcL17pE53
vhddN1a9KNISGtiMfVgz3qgfeOyJgzFmoEvAg4Jf6Kt7NOg1PmjuE/IVyvyP28L8grqPX+plo16j
NUjD+Rbv+Vh9NWxkr76siG+gZnF27LJ23FaZ8L83oQlTQ82s94OFZWsboPR6gg/j0M/hwMOd9Txr
jUNiWjNbmZxAedKZ3+tQ2jupzrsbds5jvQZMsps2ZHV7M7Ch+IFY5qc+4mlIkOeyFsmZzqPb8qWU
s99ml3RoSnNRmKTV8EvY5tKIvKzP+cLTmN1l6L254WEp8337r55uaowodMP3YsMWS2f1om8FepIj
B76Nh0DBjvvg3GGBJ0OC20fsEy0GIji4p15L5msrpgQyO9zKrwMfCIYZEfcY0H5PHbgpTrAAcq7A
bfxgGIrNgrKmwxFh+tpzMtaWcjnO6x7PKYns13g5y/o7xjYxwkM+fIHrN70dfu0zTq1gaXrmK/6D
87XpJjEqCsqdmbIMNLNiMeVD/0jj8jYtVZeoMyWWbrbL8dkMDrJlC49fYR76gNktiJ33LiEHMemT
tpJmyEvtAi+RwYW9uev6HlXtM2V7XkM/yZBTHZ30icnvs7aVQRSRM4w5VJchEw61CoQBAzPdTIm+
rIIgkZ/tuEJbpeTpQBBVoyumicwOPF4oBEUNNxkNviOnTnvnuhhxhfa9pemkF/dDwMsKtW3/2cZP
GcxKGnekiGuUZZhuNvYcyTd+xMjlHP9ll2ZQ5HPzfIIH+RadIroDQdbWRUnsA4r2m0OVxsT08K0D
CZ6NvVmnz/aTu8jaJ5yafGTJC8eL0JjG9lebj2D1s0nJsj62IPoHwH6pmLvEfENke8AkhZZgzo87
jKf1M3WzuMql/hTpyhgkuR6W0Y9kB6w3rUR9CvouRH8VYyGCjbf5xTQ3rS2qACxVIfvjLxqAFgOv
DSP0aRGVGsmY6+jIA5+SOv8IETXr2s+Q93ySdmA/p/SPHYCap79SXr86MSLXF2Fzvh9wj9YWgLnK
7qkkhREjRQlQrJvn+iZ4arv9fPp5kfFVyv8IM+3Vl75KCNvqeh5PEvRWzlswYycvew/lXpxAHNzZ
QRn1p/WbfRuTJWT5uw3Q/eoE3KJyP5yM6iACKPtIoMya/b7Qr5v5EHB5UOrHAoTUJnP/NNj0sN/V
oZizIbwt1uVcULelABfhhHcug0zcuGJtFRObDDVwalObX4hIleELlCrJHiEypf60MZochYXLrMv1
QAqJWCIk1R3GZXbjos9ss612EWZYrraPjMa1MM6EIUcDqSMftnwJtisk+eTpHuXuKDSDX+EoGIgC
6YHKQv1umFkeHXsgRk5/l4ZaethFhMco82gcEhjE6EPftA2cFqD/A7lc1p6ElreH2wROylTpvqbT
DShE5PTBabOzDnol5g1nI8pcrbDKnwktTxm7c36aXaOKbWonIt/clX1MfIg5CmUJ8uM3AGGDE2YO
xRONSLiAfCKbPfm8bWSsts3jZzau667O7fvWdaOqzm0YA4ZURXUUETSwnc4OJm1OebOVV/K1fi2f
85HITcUJH0HBcldiryS504tzMwf550i4pIBxfSIWR9YBCWMMNdhgJom2oWUh7UZztCWCcFkhFGrW
cwPyHR1lH70zrZJPW2CA4dRpwTb65gLaBJfCuSG2FzXBCXXbC/1yeBU6uimcPxwXMIoBrJOdFHoh
WXQsiNphVXNxXhMNtWdV/xPZwWG3qmDXAEjPK3flTvpJ6kRzwGL92Qqy41wfg1HcaduK/1//bAC2
ooq/qFK3iEy3QOnmN85V5UkPoRNCkb2DHRQ4/W0emxV3Ayf04chfeWvXWoeicrnQKeMQE58UmzEJ
XkL1v4dcmf+Jjz9VRj+LjyS3S/LNWQvfZsZ9zaSrQG3fkgXaumgN91p2KqsBME4ZASI9xDD4yA5J
El/0kljR2bH1j0zefgBNbnDRNn35JNxz/Ww2Qx+L1IESD8EolDcQQhRj0wrLfrBfqUYf4snLAEAU
u5aXIQDknNCSL9dBwWdiPKKgBgnVDg4UPtkFJVpCsGt8iLG8eV93yTjpbaWUi/hvBqcTD706Y7Fz
iytcE+6BCsytchCS6imIm9j0b6tH8z3M2QzAyj8lYYGkXCa8tc6RM+0c+cOuey8qJxS25TdLV8ik
E9s9Waj6qQ2zMfQIHzCMiyfFHpnTLrvhxXZgZkutLABqeJawd/qwUGfkHCCDaHlIVtAVLvwoJSpP
HPqCmBih6UzYiOm+IO5uzCFLWbua8SDOVV3V9aVidw7AQsp5TX4WjF1Phaof/mzisyP0VHEeKPuH
uek7XnXdM3Jv3QyqEg4VC7zv4YAM/X0YP3+v6fHFawTl1K1OsVzNOwJXgKVtvRdrxffdFKQP/hV8
tjbYN918/BobMFc9/8iQcn10h3zbQfg5Vgj2UXgI+BpTknWkUvHL9M4J8UIKtZgdDB2Rpu/l4V0e
N8kMRgo/YhxalcK9Rhik5TiVlFiQ7dkHhDCwPYh5CNiGTjOUpqkOCXNj+zscvDDrVcHT8d7Tjr8M
OKVlo39qV4ZAanTwD7wgUuAOo1HZKExrjsw7+yGJao0i0b+duuvTzvXnFW+UVRYTT5RoL0VoTehr
jl2RW54rn5E1iXKRCjwlFgXqRJ8LL+aVUFxvPHlOaILCiq/b6oyAcbOSi8cMHgVcj1haJ9ZvwpKM
B58IyFTp58L/7qFxQoVwSpzW65FxTgQTKCDuMauBrfLHQuspkY1LlzejhyLMa9TEzgZepXbFdJ8V
llupmAWZZ+YzTMt3wkvh0MRnHmHu7aK2MXpk8sxdNFaQoYV+YlXKzbnOzYL623lxtNWRf4ZqcNwh
cKH4srykrPPLkYMO+duoOrzLcVr+Yygk3kizvmIjaxmueVpj76VZcHKXz0LgmErfp6m1fkfdFxny
I7iE2YCyZE0ZbbmdmigFddsf6/xqwgwZXmaWiR3Ca4Otsglv/jWW1eTMjntzU8ThAeTppirwtOrG
ExFZUuHaQc5D0HcLOdCJyDgeVqeyYanQYUEdy/BpT1Jg69aa0oxYDVS24jhxSYAJm4Qmt+MmcY00
Kz914Oqb78PGpcbm1pZOMGaOCDVDWBBLVNFghqXbvnC2SCwFeCEZZYvPxELzS+HevlFIg4+o0CUf
zwmaDCR99cJAG+lbpEcgYKfcpqudIkDjPuxCdsVdDFBzd3bsbipUQtwwUG/yNd0Geh7dvKljARCU
KlIedu1ZdpSkNh8ts8h8VGQghXiGjpxzpGioBpKlbbvX74WKQSYDV1/Y82JrMDi042wmAQgD5YqL
7MR68lex2OqhI6T1N8LioeG05zGa0jzXrGpFAJxACe39bhOZmDPKSdKghrdr1438AG7vQ07Kmxo9
N49GlmrH7xJZyuhqwZIYovYL/de6+MVy7uGdHRJawsAtGLpqkrpugCyU3T5sQserVstQbYQ3Uby6
ohdINHh+ZUvVvqvbXmw17VZmGEXYWgSr9LF2EyvPh4hnbkyY4jFLqr2Tu5yKgXzfcmFSXjgCwBb9
bUccxHineHnU5UBQYa2s66VmN9k5jlOuFBzc1lWWNt5W3H0fGiDW50VOYX7OxoSTQ1aLecGYncXO
okrQ/RZPt1RM5pYxySQi1goPxgE92mNjB1zOXeZ+n7Nr55AloSYRfW4R/ZX4l7SLZ8PkYEQjecZE
MtI9ZiDvKcWBkku8ntGtDmFm9Fxon84H9TjsORVcCC8QiWYiZwjpcJG0uP6qNRiHnZSiXBaUHMa9
cGbTEvblgZEpkjJIolrJxPKDCt70ZjS1gBtAINfxj3gCjcL+pbS8sZnfPL1sY+aOSK9RruK5zdeJ
aHPhEoHgQ7P6iFSdtLcmiCJL2Zd6AxlgIyuhIR3YBgzqg8+LWwZi6Bf1XhTk62l7Eyogi0nj/Ex9
KKJXBPllWfSqLmdH4VxwtiA820EYpD4e10GzARq55E8AigkrNJoiHc83KolQMhCkZU/STF//AdKi
hGjPg+uEyG21Lel2nGEWZEB+GHV6KwBNJOeln3RIGr4imvCVomKDm36tvOuVP4/Q2Ljh0B7MyzBr
8pgOOIBBMYZDcqNVnLGDWDJTrXu8O1L9PUeYBXak6pq6gNRKWeq3JxEuwDVAqWUY0SbfPFhar+7/
qjN8YKF1O/xv+5CCzfLYOPnsEH2MRqxhjWSRIJe+FsKDEidoIDxqGV1vjpB6AEpy/ocK5uQ2KEI4
U2R7crEryPlniRDHj39oqybNVjB8Y/0wOyuPIyk0O7+q3LKCFu/ylmCIm7Ph0iaQL2uFGatbPJht
4/9mA/TROVd/4OZ9Oa4SOy1esWKaN8GY/hO6fJTk9qC8tkwURFoRHopTu9fNvQTXEJ/C3ESr2KZ/
q93nf5X4Cs68pYqRkZ7v6O1l1ZBmIAd/iSVoEMXSamLTBkO3Em+vTwJ3HjHnVjaZLl0Gl3Oh3G6m
CMBfgjVf7t/bKeA9aWGqPuXJ23MN40YnGzOSwIXgrpt2r4/rJAiybDs4VsbtUIB+tu+B+O0RM6q9
Iss3VjZNn1lpq3f/Xs5qTQtZidiBlHXVvpzBHUHdkjAzVNpYb8wEyfIoSrvEYMYSfCijl29D1acT
U7z9M2mg35cM9tQHxg7U1xhJr3IOcGZRR2y89H6zHUf1K3ubxjnr1sjrVDEC1RuyO6D1/fqaJN3s
MKUQKyNJ0t7YdR7agDf/3kek8gHI7XdFYtcz6YIY6Sa4WnABPNwk5qOr3wzveu4z3H1UIhvDMQy2
MLMmhLhIjZ3hXmIiSncYBra0jXGlz0y9myfuR+OwbBFeiDzEEw67N6rHOUVN6Ft0Th9s9YpHnQOn
qB3166QTqE4s+w7m4fdZL+7zXoCtvY9sVQwYdtmzHIuYQHBXPcf8TcUtDGUGbY7mSlo7xj1u4NF6
9wreBnxNyswcuwPjcVyJkOBD0bSuznGBdTDexUq9Zg2VBU4LtDmIt6qVhWxBXiHB6GsfpfKp60ub
+UsdDRBeS8W/y66sZLZqwfY3byevvGozftZ1TRHXqXEtquF07U/yEXQjNuAdTMQca7AarggNPlCc
fDICDGxc6hPmY7WCgxVve8S86jL9D5IvLCzpAcjAH0z25d/87MHCQcQ82fKduUFpixhGpbzW6Aod
kpoUn129qFfEEecTUdjjDXnrfwUNAsyPmtM3HQYTYBNIV8RJdjpmKyT5YmUyxGPZSsI+y9IJiNgc
hzDANhiZyVbgMSTN8ThRk1hyS3IHXEMBdHrYJjwALMz1pSnh95TctX8MJwc0A8r3xXqeHoNYtjlx
qeoPjmJHkrJCOwatBMAx6WluswflNUld56Y5/FkO8O1jCy55S/gsHZM/BKmYe4ujYHNtYUJq/n53
rIOhoCQtXOFK9w644STZ18TrQdZPKwHeUjpStVdaOQ6c5RgKf64oYRiw/PYg7Zn2udwzaqeHC1yw
DFnu+9x4Nday4kb2uijkJdIvKb2pmlINcYdf/NShp7GcPazyT4XK13u+GYMRvx5ZtWHx1MpReobg
yJ+jBULW1Li6HjKuClUMKJnfQAgzUHSXBNvkXkd3T9esXm3lpyatOcOVPVus+MwxtU5gYLILblfj
8V2ljdzXLWHR053l9wxMYv7wWMZsOrz9MnYM1B5ZrJ5Oi/WRrPGr4+tjSmSnvaxF4Clg1Bo4JJ7i
eLnJogA9ykv7O8Pd8WoQqyfRqnM0elh9USRVWyuwLDuI2XFRmqL0ahLXce4JLhcRxoutXiNr9RRL
A0d5MX+K7AtP06gsl8vIA0A0dMs9/UFNQa9PYb+DEEmIzk6ROdKM3moszf0juUBfb65hFuKoBAZn
z1Ns36VHuTn4GqJ4mHlPZx+cSmSmH+l6zSk+zby5XnenyNKvx5BEYml+UGGAXU/GIuHuceEF6hQ3
6TC2SVUzPk03XliN9xZROAUyNBAqu7SuIY1YkXu344Y2LvUEHAV/cBeqiiEB+tunEyjyRJWV6vEz
pBUHLXhH9DXrURfVN2mvhy/E6eR7btMjnb3Sharlnyv5XCURSvrUZrE252IcNuHESTRchGsa+ax/
gH+3lLFcns1caGX5VX7kvPUGZ8+M2MmFDJf5l76EFlpR09VXkoftQKf9dHCoQB74fJGz5oaW1qyI
FmTLc/wVuCDJwemy0y4u3z6rw6unbPRTUkqkvL0qrcKgYoX+9IIw1hd0gSjsgyiGzbJTtywG3sW4
xifjvmwgGR6Jw1LH7DyuzxgkXUaiL1BQuhxYum98nQBryKVPiPsecrrGkaqMotxx07hdWdtPU9Tx
pTB0efBO+YTXfK/fNnqVOiFxP/S2eNGFXPMo6RSAlMrtVdIRWz2KhXbgFJeJsBveyXFR8EXqJEFb
4QlP1xqHe5/aWtp5JuJH2UiV0B7INRgBD+K2UDO+HN/d3VQxovRfO9O51ixRudnrGk7U6iPz7FO3
t6/1va8ARbWMIKikFWQ6x+4UnlU/lMRdoknfgx0FMeCb3txcOr2xk44mIGSKhOCMWhFEKYjJ5XJX
0JuYBnDLPld7ol4K28drlFlEZUzCBR9OXpSY3unyxaYackviKZEKPrMMm1tSeWCN7ECfCAaMaLrn
rtZsYbQLNbK+koRyei+4CoUWhvuWiAjjc12vkOqoJhqcM9QAYJjsCPeXURU8VfpSizGn2fRP/B1h
/fDqbLeqGCWi4sUbG+7lROkXvXInabwPBg4sPdx+mlxXhMHGNI+3zoSln1v9iZn3biB/Uf0HgKom
zpibIwgun0kCbllycv49bbIkytx7Sf1NLiz5AdLQmohCj67+QaIsJBbMTBO/8/2ynFEjvrJ2DzTu
AgX2AAumA8ZAmQvbjCvFFYB/W9J7D/+Q1vl/4l4XZytIizCXmtApQAHF1RqMT4XgOIwotrJjvNYI
2AVsumrwPJjYiI1jW2akcLmqBkcR2qrNBRdvTXui4UVfaHHqUuW1vmfTxbf9xYDI57KEDEPHvs6k
/I6Gmx/ZKjz8kQVsP0C3tNaJY+6r8R8cXmwIDILniwye9c+Dr01bGjm2WIkYkd8PMJcVoFeZRBBe
lTRoqnyycBRVQ5owZamPjnuviGkh7Ww4S4RV83dlWc0/hY2iPIiSPy9L+Ey8MF1QObmGaVlyR1M0
gNkGE1yjwTrD+5fVRc01KSXR4hKX+34eDTlW61U7aAhqjwC43V1sHcK0wu/dlSKyC9HOnOxNH2et
TTVvjQ6+UFJ0xcoRmKpSYQ82PHn4aiae2Yg1dcw//hV3FAurIlY7C2GIOqjbdqhHyLwsdS8Uetvc
UdSpW1NHsd4wfkWy34ffmSP8L1ejskmzsge0uWoy5J64LttTCyFT9TCcR26R5vNsq7Et4Pc4ptby
t3cwycAciRtO2JbN2Gqlju8cfg5SL9sREAzVoE2If+3Oh8RVZsH97S9ebhx2GFppXffIsH/2yjWI
HbJzMf/0Uj8F+19a9R+eFWeK6u8eQjJXkJNK2fXXPx1g6dQMFwt2sDcREiMB8K7Wj4QeaQ+MMKoF
SzHdbFkFP2GB56mw2pVP8NcUhGpvc+xL9PdLyGDUZnCyWHNMFnWB3Nsc0BSSzKn/xTO1vOlW8t9W
shrmnzksp53PpF7uNqD6cMU6cpoQIAicvxtHlE6PyfMv34rX5iu56moPpKHulp4Kv/f0MLwQTxWc
WcGd62bpj/QA9k/ryD19AurXyclHn2t/P2LHRoADfbyA6Y5lfRlwIuhyv3F0sZQnjBPV2Wfd4dp5
JtaFHqTRVc50uC+qv7wjszkRNxE3kE+Jy6HN9+tjjnEVxOy5k47+rr5E1g3mLq1pwjFPQJaNxR9i
nZTQsBqMPE7YGPzKz9gMv9vCw8zZmVcjs8pswU9AxOB5vJMMsK1om35Eg1HNQz7uHx2damG7jaO3
w8nlB5PdSS+5v2UzCx8M82ummPTGZTIerxJTw5KiPD44m3NC6CCUvv3MSg5WAC62+1dYF9ehvJjI
9scYUmqrlKjPYyEmX7swh1SN5xNtM4HIOXssp4PqwK8mqJgK6TYafvCg31dvh4FqM+TBPcvkIBio
G4JqQpGkhGkvaBFGe1PnHF8VxOS2Bdb4z3zKz7H2nsF4FREso68D7FWRW1YBwahgYSK9ovIZDjQA
Wqgz4jS3IQkgqiKyKS/dvklDTlBodL0qE8SP5OOP5boZ3nVvR8efZF9yHQn7OspRQOzRhfMm7O38
i568kyB/YTS+0Hu2ytSVOezBp7eOep3daw4KO63ENbSEnp7AuHSoBBSSp7D9KqrFUadY7HAB22wP
91e9cptltalPQee6qecs6/1SI6fyW8vLe6MLCC1xg5yi4fTVCrT4el8HiGvCDhmD9Y3EBFXcOfX7
LHn9C7c4sBJOvGwS8KyrO2sYPmZK5mOPQIkyYFNGrvnyedUYpOL9byk3LG7HWn/9JkHx72oVQvxE
LglK3QpM2mhvktWloYub6KFpQmbQ+nw7R1YgBGq4N/eKBSnHSxPXAKQ9tudWc2YR7FF88RcoRRqu
x0gxF1yQ2newTXbVpuylFMszeITvLTFZEvvZ8us86qM+8OC512wGqz325n1H2kHw8v2P7tEuesF4
DsodwUz4jMlaq/9nJPdoyGZAc42CCYhiKp9T7if+TjoTQsWAJsaLGTuMeE2maJUjQ1Yx6JnORuCK
LFVbsZQb04aEV0QST/4r1nOl/dFwKVCscu2+8pCqQr0R1SnXo9FeHOocGmHi4JRxl1Xtx+G7Kji4
h2b/8Ac1Mn8MR7zehTIpzW7uTUDjsjPJnJRZ5eKZ+lTGhCDyQrZhH33ywAPy3kxQ206Exsi95vFz
4k8mDjrXpv4/pxxI5yn91w595fS+bK2NO5x0FWNtDDACtQh+qXEKAjt+AnotRl2i7xw1pbMsSrHt
X/O5OLaPm5J8CnAhPngbzAsusPuCBvwvUP5fU9EmAQktImrG0ojc/ZI9dmC2MC2TnxvrbnpFDIU4
8yqzPayQ1ASPLyKkNfgyfJzKCbqO3x4+kzdZwNAdVoBtk3/fQ0K7QvpKeNqezePBs73NMhZoQz4t
rleC4T6o2EAIPkaUrpi7CVWuPjJbispiZ9JxR1CLVzKQS/8SUeuFHQmn93Lbe2wPD+DGuP2DJPSL
XKHtc41mhX0tGbdhwoh5OkuVFwg+to1OZP66q4EdrYze9rb8x8rL1BM9W2Mss3uR9+qNY5rWYPNn
eLM2jZS5DtMXUyCnyxu6snMkp4BSgR93iEZWtnAHSUhdeiVxpbEKMHQmwuXKMZbFxwedcUCXbx8T
CmsI6GMUg34PdYyGg/khAPBKNRyh5eR0almerCI5iG9b/d0bXMYvy25vmHvJVMZg6f0xSZ03oRtk
XqVLIGUINjpo3sLMaFWwV92lSofNqxGdreGWpdWppIfTOIrZMq1yADlUQwEfIAtQM8SptYJ2EkRR
dC8iKISgu9pVZIqI+MCXDWsIEDT+Xjib72JcqzxyxPjc2/7FFyH3RsdLhYJn1CrXwWd5S6BYLB3c
3Rj+9z4nfRkIKU7EiyE1KQwvZLnGhsKjraNtr5KHAG0BEocAETeU0Pl9Fja7eZLTsrdhomE0PtwK
UwRU+4peqK7tsKKGhz6PXXNC+Qf/XmfpQKC3Bzbxp5McGcShjTMDCuhx4qvK6/cIrWv5fndp80pm
YsnbQjSBlx3gJdjSqmkqXD7RIBqE2IqfCTmisuxNlkqBtdmwoXAIUNzQeEGK5/qBae64yxB6LGz5
nxB+lkMSVkUEv5tFcrOWdXzv/RaYhi/UNL5kMXsdyDWMqsXIjHeUDxyEdHnYM0UNZk+RwvnaLj/w
huQPEUUAag12+tNWFdgMXK7a/K4ibu0617IdgVQCHRgT14YLxwxcOVKnhx/ZNbDm/PnW4keVti0D
3VR170aatimvLY9HsyfNXBxzfkHW+43HTlLu9lkAZwRYZommyM2+o+hhcUucToiOj2Kv1ASQiOxU
HyUIRJ5fcvopV4dIqaFwkcgjkRbTw6cSqsz5TD+OMkVAj1o3KeR8zp1JzN008bt3kA4xAsMb7pEp
wtpD17GSkc75Mw0YiUAfgtEoehKDixYTwUDqssusO8vam9kEtmeKEB0n68EKmE++dJVNk+J2g4ro
W7lo5TgAwnjXX78H4EiPESfSCdkfXWHYMVg3SU7cSOkDEZMvrGKQepVY4De/r2agYVgW0/0FZeqH
ty6uW4PMyF7Oel4phps9nNdnH06gXYH1Q3whFXLe0QJcjfaDqJ1W0/cbqcU8rUKqAyTTyd60DSRl
N1pnNrAHOarngPqYm5hWXRc3NppTxzmIwFda0GnLZpq/rE4d6S5c4KMtmrgB3eyIRt8plBlxgLzo
qhHBuvjXQFL1Lr6Qerq5RTTymcgDK2CTbmIkGZqDIFHgWpmHxVuLH7dKNSPJKSvF3OnWj3q1hGn7
CE2askar6FPTY9L+dardxqmeyVSgsb5tZaILOUJwTDbdoNZ9xuky+pJkNNFhonmuaWkZ4ypmpOQY
yVPbcSLrTO2tRjkqpERkHFTMOMbERT/EarBSmqGbb6aOyNgIa61z8lPH0Kl2nSfI7Fcc2ddwEkYt
2xyrwNJonFoqI2BLMDX86Otor8fJO/E7vMGTk5/8/w8i40Y8UzCp5jBtAOqUEN8VkOofyB60m+2l
giRWxgkSX0Eebf5TM5LTi9ikoMH3sjNwYzGAIRjFOxjnE4d1FQ5kJvGQw/tckO8XR2CzD9NsXB93
47vVBz79tKyzDvncdwQI2C53DSr7xj/BTxZsSz02O+w+C2UsQ0mS1kgwxYOgTI5EcOXhygU8z+jX
0hlsTnM+EDIItnTLFaRCC0Vnts8Jm5COOjES4DMFilh7u7I0J77qWgbRDWqP9ak4oV7X0C3IoLS9
QD1mS2C93Ys1Ofb7rTnuSIZnlMAuYUZoMCtk/NLWxa5E5kuF9p1o8PX8sZOxbMxlDwmUQOJBmTSD
R7nn+jOcoVn5zIOd788TVeeUw8/55D3UlK13ADlaQXbTW3aW5RzlnblWqTY5375AoIAw5TDR2ZpL
1JsLyJg3hhR5Y42acYRU08kB+SJTlu9NohDNhCJXSpp8o66t76oOo5BuvJMWA7ZqkhJe/owEloEp
X0+0YqpM5OXMipdS8V/ekdv3D9R7ReASgJrWIdTfBPYLF/CcEF/26qwmSfpsEZjz5jE5vypdd5WV
IEdwBCpwcQoMDTybSQeH6ncoYfL2pBBlGu/xkEZ/onq+yyhJhNOuG3Cyhor9ddji7Vv8pVxJIyMS
xi6a7KDnFi1Oj7dl+ZKV46ykhkljv5VQSQhqpLC48iSO2fpLuqOp5APWQ/YseWr4FFWf9bLTbebN
ib/Bg9NU3ngiG8R/0xl7+X4pN5REBDNk7p5oCSnF415auA+n9hb2svnFFGadgUwsQ9ycDrgFHqEJ
bSj4AEx3FBgS3Y4/v1C/UN9qckwVtMJufjp0LWBrw+m277TGlmOGuX99z2re6f8yRJRF3D5Eyag6
mF6bbR7+Antjl1e5uCpOXXgTe5ZHXjpU1oy25ofxXIDYN8wKj4j+PKHsBJy9zfGVtfyUpumyIadY
ZopSYD5PefV8qFFjtYpxeRReT23GJGIf7q0hL/34DMqEIjQnxp2Qw6oYQlbMx3dr8n2webYlj4hR
Iqars4TCpBf4irDHVbhPeb+r5EWXs5RpYNKtMt5z2qkCe+o7Cg4jdBSMr+JFr8T6Ls4kCIrUIlVL
Rjv8+UaMk/OFZ1imAu9YzMuam3o8pVAKXZfT3D90BQpC1WIQia7S6K3b613N3wPX6WKOyEYbaLr3
cQ1VtezJXOL6T3qeGt682WiDvCrY2W9XFIU0g/KhHW8hSl47cqaA+Xkro/hrV4kPwK8Sq89xFKak
zswYybjE5NJg2DKKB5ucrkwhabzeb3B4sVOMbDHutGcTuUV+Bxzb19g2dR1FJKz/5XGJdCFQ2AWO
/gGMWMSX3sWcE30+eM8elyuT2/0ZbUtj5gV7yvUm8vCpLDt4WkgYX98v3sFT9I46z+T0LLTIlQPK
j5yCtqGoImg7RSRt4W9zmHclgrgMQmz4PRH1rHP20/PGrx9ySGHsmymT7E7mLuYqb+Dl4qCbNyyI
ErZGkDgaqPoq2nofBj1QdEYRe2PDVS7ny50zcTosbpYBSMB4e80xP5zs+dYC1gLDh2dDS/EM1YVu
9gU4qw75wr7bIl+x4hz6agGEuE9ya4uieDHO3O40uutjm9iZu97CHBjpIHGrlytCBz8L56gKJx+t
VKqxJEwKdkKr9o/0AE7BNg8SPZl0bAgm9fv9bBhcn5P3bEdXdDDdMPp5XaiJaNxhysGgqNcTREdL
3QLd9olUJBW0WCRn7JzowI6gQDprlGHEPO3PMfZEtPCQmOopowGaIkmFHipBxD0gm/YHjdhc9Zja
UD4l0b7oOe1BxuMetJnbw5I4qAMLNkAdSK1AOzZTHQa8b9Q7oyet4fRMattIlyShOoiqoFun15cv
tWMSEEpD3DHBNbeCo0qWefLPRy5GerRNUvh4zIcWl12gLlTpd44T5HlFJ18RfY3XmdiDCMZ+OtUF
e5VH1ausHLVwTcRotcLFU2mC0NKv/tACyiCXqlf6ldBVIS6rsVjvKoLHjfRzo9VJ8N2dDBl9aK9S
zDaw8dPI0ekIq/rqmi6P8dRfEzx8S6Pe75id9YZqLZS/hItMp6wQtaS8bBwVKSIIiWISeq8iK7XA
XjAgdXVFN1xljxLcyaUxYp7qruTsu60gBE9EJHY5QGRB+3n/lfYIGyswsYDcls/AKTkFO+eTdVy8
1IV7Q9atCssEUz/NQba+t7AUO/RVKHzSEbYsv8jxTRspetk/uK4rp4PdDPxMAgJlSay48/HtvOOA
9r+dtiejZSXKVEFJ9ZRBBiENr+ATxYU2A88KZPC4TsoNZ5KaW63DUIsa365KkJ3KVqEpoc8zUs4s
gXv5vkHnuzagtUetyS0l2NmHdGUxFtAqt39dpd7gaHVFmY0H1LjXFUYa45xOlAGnPpMCAKVGURtt
Dpo1PjKVMLLHoahMQ3PEYevkhDdubyMfz1OwLFHRdm1YDgMc3dWIwSgxOWkHVPledJz8yyOmE3/X
P9wuyoUVi53PX2AP1qabyYpCF3drQwyc5fG3m2TMqrFHWOQ0mJggwCye8yb90FETsOSxc7Wbmyab
xGLl3Ixr1VUcO+qSJ/KPY0Pjn2zEn4jA9dG0cBJTgzwc8b3IhRTbUypKhOBvb2U9Qm/0VjuKqQX4
8GRubwK1aFH3f+RHtQpkQKVbnHHIpZ6T2Epkc2xaGN/5ZfPuGhLnoqQ0dVBuDxyxW618hMLxYoOe
Jd71tmUOrKOB86t/cQtovwotXbxN+MrMFYzf4ehbyNtfKDtbIOntFlum8QOrXiBb89XbRjBe4i0k
5mxaw8mHWHDInb1FA/JquOmZI+eH5GjWu30eZdV4Rsq52lXFfDbPVhqjZZfVJZfTYhnTuUJvULTw
zC+7WCDWEb4UvbLy7wrRtbrw1vOfcMyrLqTJfYyapk93WCBxotlbECM2keiQdE50i6YTp6ZrIy1t
fqAVpQinGaoCnFjY5BsmoR0GeQ3FuiURvIEbRvIQw564k/uBiXdqiQ8yZh6GDJPm3eYMdCiwFzIy
Ee+MSBsJPn76ymlUa3MIjIYAj2n6NZEEGejePT2IhrehsmeaNBQJJEE9Vv/WY79RpWd5oqy4nUaU
qGG7fbtKFkQv+Iphlu9TyBxdwQUj24t47NL27ACGOGK3ZPDoN37JU6JeM63AbEgsqFvPEjjabycK
zQoDpBv0nukkcF/ib9LXJVwr5lyuvnSiNsxEHOYxkvIgszAITL07cpNNq3/bzpcFRzdzJFr5xB/1
VtRB982apewLutgLD5VW+J5FgCQFiI8fJPuLAjENKsoVnO4skbG7vrloRhQBp7ZyPZyN3CPrlctK
yxk1mO8d45i/Nldnl3rZH14Zu7OjT4UbvInpDAoyfPe1/zClYMuuW6zacxroHm6vXLIAZ/CzTDEH
drwboUkSo8P9/HC2MaPDGq9R81JM6j6aK+DPM4jObuJSAoViSVvfy43sSycBXuh6RRxmQ0tce0lG
8wqTYzr7ger001hPTuCUb9l3hEmYACw9Gr6Zyxo9Cg9RwWSPaB35tB+vu1IjSKgfKNUosOQknerW
g1y6+ck8YP6l0W97hbqmOYvo49mCgs6oMcXuFoqi72Ge0YLxajBsRRhZeIweEwpEFGbQtPiKKKIg
Pe9YhAt+LfOCKdsRmb3pWZPIXxpaCgdWHC0l3D73/jvoBBkPictiaagZ2IKygzpKFUFEZRePRBNA
9TEkMHS/Ju36tqvZLtC0lrH+dFVVW8PeaXZ6HEHfYCDdt5vwAxDghiSYPjgmwJ6+5jsOdA9H8MBl
DBpQufSIAAr/sTT01NXUcYlSJAcvDqmBCcEsgIAfRHwUl7+jJDNKwuJdO7ThSovuLmvZPIcwx0QO
knQFnjmIQHasnrMy5AKR2zJuD9YkwMfbUxa8QLUJoKW0V5IGxHXv78IqEQOYnmsqjIrGgWiIxVNI
a1RXIyHokW07Tfp/GykD+X4dcT5A2d0lDh5/pWc9pRY140CQYpbLvFMpx0FlgpZdqxbHK8w+6EFl
rHXxZVkEUy7lF7IHb/GDEI8UhsH4w8I0ZoZogREoTbgcpdCMMcO8JR8L5zDUBRR2kE9VnTL1+BjM
KYeYky4mNGlGJFycKmKUFV+ljUVa1n+PB00LcFalwyfVOjDnhjoNoFpAKr3SQ/lDOXtWLyyFNPJP
ddlpF1DiU1YPHB/G9X8KgmKhnhBksXZAW2AbQeajGvryQ3ggnvDQUVoDKZ07Obf7K1Xuhbjv3wHX
AE1GnnmSEAifQ74aputYaIUHJJS+YzY4SEi0vpP3RCZAn3lHeZdY6MNxLsjafVgHvxXeZIu3/K+a
DEIQCPnUpfrWhMPJGMG3FV5xfH0SaFk9THi9B6ULTAzteENeZptjUHIZTmwgUNb6jfoNkFGTUAFG
Ufr/nrrfG5/ltEqe0PYDPWAor5PPG3JbSEMGtMgZn0jWI5bYInm1K8GjKFe2+GPSh1TfL2AAcvbj
t6MdEdC5vy7LOVUz7njQxncBHwylDuCAr0Z2BiSLVG4cr+nXTIl5BgqVFiZlYA7IsaKouyIw2zkQ
n8eJolNdp/PQHgo51pW3tdsvMl1Xyc0Qp2CiBrbj+qULEkFvXoctziunRROLSyoIu9EHhn4CwGQl
Os16YwkncgX4YUHcSc1Hp1wmK6skGGhCwswoznqer54sULZzNNij1PpPmCtuvKF94KtlXLu6Hwek
OKstcHU3ySKHu1mXwr0miP2py6qx6KQoetTg1azWa1kEEWrGJvSbG2iZwQOsHB9xs1onWWOgQTtS
aWU4B+S9QLuWH0ejetIdmmMVEOJS4IOlitzNzX4EEJP+D1LDUqS6JyFI+oLs0gJ1yvCl7ZEcg9U4
yot63aX34IloJqVfHsIGHY7+u5llxxm7E7ET28D0fpgbQ1ofVRoQ+7CZFO4YO0LkbxdoVEv2V8sL
nBXyiLBJ/RdYHy6M6CkLnrYIG6l6c1ja2pM2iZ/ZozufboElfxjypoWLTXlXGyhQyQT6MGrRkI7V
4rv+LJdXgBuLap9qYMC140uNFRVag1o2JCaoz23aLiDjEVKAcTai6uLr1KlJ5i0RCuIRQuy/2ikB
qFoslYQX2ryHi4gI9+52PrPupaKHw4JGq0DhAjahSMeV/cVkIiRMQGivcDHZTZtHPEq6A+9F1MqZ
a5wjg/FSPcwpYXLNWiQshFMAJONzvYZQMQOi0PDiK6IhTKWVMTv3Sz5hYYZ2rNq4pj88mLgycHtQ
8nrlDdchnP7OmW0fKHFNp4NdskbOh1Quhmje+mWw2uuPr3XRMZ3lbVAzjoraONcIvivF3apmGlrL
UkDQgXbhA4G3GgY89UCmeZXRtiXHi70VUUnA64RTuudeRDPGPXyu+nmclqbif1S5+9MR3bE89+eg
yl23Jx4m8vbm8gJjCWrd2gKCjc0WUt/sZVjC5sXP59s/+y410G8YEnLdPLWr+1T+QB8NcsddkIrB
cegfNbDT7zlUV7Z0B7pmenMoi+HYf4BQVZ5R29bNQEFExw5C61K0/zKH1R9DfgwNaANuV9VKW6RJ
X+c2apqofLJg8jK+cqtv7z1b6IBOrJjLTP7Ws8XNDiL52uo0o4bkv31gMN5VJLT6yWu1TUtlJyvk
XECNZEAgZhB3EXoK8edvPa3wWLvxvRcYC5kbWrm0V3Ad7IKp1bUHlpqy/ILFfUSSTf4dXNdM+kye
7i2X4Slpzu4+L1QmKfyt7sgN1Ai3rzIDsU0CVFYK7H1m3bmTY/M8nXPnpvLkg/6CJeZyZvjvO9rz
uOqDUNLJkBC1IpLqN+j8k6JVIkw/PyVP4XPvJ3j7J3q2XL4QxhZzNgIICDjC4/JYAY75igxHCt2h
LiC7MkN1f7LX/sRcK7f/dlqU8eTSAAaBpNRXk/EuobLtRwUWR7izNSRUFO9ExqgxLus+R4wOkKSB
lg/JYDtA17HGpJvrXk64vCXnj9X4UI8xYn+aRZMNIfiGtsFQ0NofKlIZv8rG/fnepJCIa0GcWY04
VLAZ0hH19RttPXEsc8ZnA78l2PCAeUBUYvc8L9LppyvBgtyITHZc39XdPqPBJZbeLRSdY2W9y4/U
05vPnKKoZZXcaslBpw2r8pOYDouENINnozE+zVm+Qe8wxwHQt4pYaokLodqvzpXYplXEIGlpTDqK
vTj2bl7uqWNF4HO9fFkAByDAm6htTuF/AhiRioOTWz4ZDn0wQpN8ySVnqgoBWOSU5OxP7XUEypxv
eftyvjXDU40CpmWhSl6ldchuFXTerKRmqfTbzJ8xtw7BG0zAk83P77vHTZKfNNoHIL146dCdUxLH
lLxf04oKVry8x7dEtP+hCkzOZK2V3UCl/RKis/GREHy+rUGLAmO9IKVFbxEkB8oa7QovrdycLZBz
l82wZj0slTnEL85ZEl0l+/Meci17223dtHup7zDYdDXOEVIGZ5r0BQ5jl84zaxXgLrh5NVPUbIcB
G05SXkkPIdPCscx4U06Drox9gb9UmJpStaPSHTt3SQ0haAE622FjG0X6Zrj2WMs0rpLvKeYvnDF2
crkdoLUJtwxTApl0eNVrMUUTcVDhE3p/iaIdja3JI++CJWrrQYNF1up44BQrXWXlFqPiaR149fCW
7hNz7ptRYlXBJgCa7ecrQoQfn+gUwUdHWPAOLwzkixCsAp+T9sfi6pXgoJ5c6/+p+ueQTvZ8bIwa
q8odO39YLPoOml4hgEX8C9BZQuwJTIfis5+fZg0hlrHDEFRCzoAkLmVyukHKo5c9LXc0/QT0kPuy
Uad924b+xEdAb7CD1ZT1q1i/2h0PV9RNz1ZfDfd+ZiWy6lfOKrUY8pWkOzvQtgkyWx6QmyjtMt52
xPiYpGJ2h1zmRyRijjWLHG6EUTu1uG9agyj1LrzJqOdeDjzmlaka+Hy5wRZkSqOMtZ1aGux90n1R
U+QU2NmS+Jf91heNGmcEdHlsuxokxVSYLTXFFzbT8TKGwcYqkMC7+STDQz1zw8fux4FdcXQyq0Q+
AiTo9e8ZYgPzzBJpMoT7BPTieiL7wQRLIOi9/sSPpJ5R13R+b4b6dSEvrQFU7OaxqGpO/1YhjOWx
GJTE6IgI0ZEVcC/HaeDb3FZ9Iv12JxYlm0Rhg5sFAzfNQ9i9uHQc7i/CnONzchY4BFZSn8nMIQPQ
VgLmzh9K1grtWx8quzXX+cLvSbqyC9HufPNyyAbehSvOs8A+e5VTE6PcjSZ8i2MLosHlTArpz48s
7uW1Cy9p0Pwk9SNHcI/OY+81cGJMML5oGjYd8bQYdO74U+/o1ohbH6LzrN1YLIjXB939WBm1Dstu
w+FzZvHu8EIy/LIIEJ75IMCUWXi3lm8EW/uwQRhQ85/qV2GUVJZBDx7JMNWt0PzOk/dA+R64/1yK
tT88zeRmQ9fAZC/ijZtSNikonPYUKqD1HV7isTsaOTInoaRNrIW/sxXBZUHB2Nd8p/BbRd/4OhR8
Lgl1wZ399bcrXYe5dGUZo3ebDWM1kvGl4mlIbWhH0IDzOuA8iToLReXmWIaYzzhFONPd9hUFY0Yj
80W0n+x7eKhQq5P4o27LN3u7GURf6F28yyPdwXTYUSvR3eVsEfVifjjRJJiHTzEV6U9MCKzpzO8s
VY+ZVIxT7GaSLL1jLCbMgEpYTK1n4Op+PCvw8+OLcMd4U632AXtdALcvhU3ach6F+aVtnmK1/x9D
ot6zKGs3I6dIcI0XgY/6bmeR2RBKdFQGFNtCqqimpdUYOtTtgeQaJOuvqqj5/gbtcIdMq2qM23OH
hr1tJug8DV9ZidgkUzbAcU6r2vhemst11mRb0NeQ8bpD7zKzFLVsQbyD36s5j3jD2+xFTqqQOIxT
DntsEC/FPN1IvBjKs3tWFEoWYfZX63KK3hit+yAGZoadmiIvFst6hfL36oA598MS1LA/j89puNyI
gJv+THqRb05sOcHCu/cOPeRYQokQlPRD6iyDeQ/VzHTehPMOBIZ3R3U0Gj+v9HZFlWcvqaGSLp7K
ZnEPxZESy+Z1BuAJK0CsvRzVHuSOdqRd8HaYE7CzeLa5Q9WrJR8OlCsxIo87fyw1q/y8Ugs2QUAM
rE6wIzkcQZM0g8VCE/cwB+cX+WuFZ5ZrhN4iWCOA4jgiLGBkurbReXg0PqGu5SceEsNK0aSYenZu
kvTpqzBd8Ac/JajHEJWpzUavg6RXQRA0biWDnOaVzeESCwbPN0r4xjY2kbk2JJJlzFnH370aavT7
d4k+8RVb3POFNBeLJKiHJatn+qf2L5xuWYqTiucFsKLcAbDzxWsnIb15mzE2ga4jCKvObcfFalSG
E/y+UulveYsBf5RSoMwueSop+Uvrfpu31IMOkp9yQ8VQQFwb+yGdBiI1sqt3POhs7VojWkruEqmp
SOpm4RoXMoyAwRiPMfVjqxJEcIWGXFzrGjUTT3lx4iemNqe12GM+9w+Us8ZzDO7+S4vWc46snEfq
jwUC2J2LsDryOBe5w0sccMh4RVtMJMRettjHquy8bhRtSVq64N17Ww1WvuPThM5wvTiPvoGx7ErM
+DIqfth3cB9TNccY3lZo4LTWqZT2Q4ToqiaahMielCQgpzuYeLMGSHNU1lfjVj9N6VzfpZiyHDNm
3Bm8t95q/Bt6hk9Hy8TnZJe0o3uEPA9gVQq+xpouCQTFDTW9PzUJVHtRhFLuB3dwscC3bwLam9uT
QLv0poktB5Kx2diK/zwOvvMXdukubUZQ4F/t4VnEsSvYbLdAccrXohguFch+52mZB7U26Svc+a4a
NJuQ687v+zE3BlOTQzisB+uEKSDeI2pnFoo3HTMPK40Dcw7ZbjAY4RCDI7M8Z5b5jJ0k419QeptR
o2Q5+2ETx1oxEQrjcHzWOevbvRMJkMeRtVZFtCtHIGRwlTOo9o39GKw68gLs6uBoC4qEZPCk2I1C
nHZD7LcNtyxz10sekoF/T4KiTR0fV55WbjxvJBHB1yDorRqVcIUP9HDMXI0pSCrJQ+xVBVjhNlSN
bMuEk2Xdow1nV14JvgjbDq3Adtm/yOMVw7Iz5qTVsGb7lyXH3YYCqKvt3NGO1dnEr3r9QCPlKzlJ
rmM4197YnTBp9Ltn8gQI60jC8zMIRxn9auxp6x+sXPmH0e57KESU92uFko1pPU3/3fY/6XxI1yC0
+yH3fI4gWyYWSZUY6l77brAc8FTPNqrMRWiokxLsLqDOjM5mQCs5ojYVy7ClIOQryauzh0R4kWUW
/6W2IJkOe56deJ4z3kLNiNZRAhLYu40pGYIf+pEHKMm0i2/6FB/CMvEabCO9vyBy1tsQy0C9rRYy
dQf5/BJIJcZqoc0b6C8QOpYjtqreW2KfBgVmfWDFmjtjfj0oMl4b3pga+v6LDhx/CHXPYwr9eH/T
Pj0ztxk5byv5vUWsrlWgyGXRMF1Z5bzSZWyfPZ3Uvba43KmjnxuRqz5xexROUR+ft1IPi8jWpKkh
OhFZp/v/sAxQMEGl3r992diBcaxoXEXlxqxrzbkLfp/JmUcp1H1jCEsUciqHLznQDvoWdO4haxW3
rvH0+v0/WSmtX9xrgbx0trt0U+KOPDNFTyF60hj5IEtjUqS34mqYnHv47JVBpLR/WLL5bC8hfJdz
eJo2BLe85mmvDAkZYDnchkOw2A/4liTsWbpNaEx1K0lLYsYfLcITptoMcjFCpC61aoF0A2PWqcYW
ipnVpeGudPuDcAJOndwSZWGOdLIy2vHO/2HVPDcF/YcF0U+pyd9Q88MMo/tzaR/jitLfCHCP0QbS
ZTXiZVXp5MWmgZoS5E9SjBhyNXFIyGYbg5PRDXRsuwqjT7zyZ5whsFPY7vW2su10SfAGpJiS+z7z
ABSw6AbMEMul01XZxao/3RwhfVWhWp3WGbXELrpM79sku0j9IKfR+hXwLzjmD78SAXwGEzfNZS50
nYTMj+M55PF+IOcgULZHkFviMOM2SJy2LVjpiT/kAgtknjcCYrC+hoseHpeuvmiyIuPt/NsUuYZL
be6RQm207QLcgMqxglT8HTt7l4WZcqAUHNtRZKJs6yUV2D6EW5Q3EoEUon7FzhSfbupvlqGWOB86
JGqYKOz9q4aRZ6FGXXz8+Ncpv79z7v2umOJw6u2Ow79K8PViSxyZC3l/1M8BRkqYsOANRpN93RRC
fmUp6DU9dVwDd1sRmysbqGOgPTA3Y0Py+9TiBq4qoULFQLipvLjXx0a49RpbZco2VaztD0U/jLIg
8nCjw56stQq+xHX0zYuUNJDwTfJypWpCflEJ5ESnlMCKg2b78+VDB7Boo3olKQv8NXTeDb27K86K
2C1K7yYWuzlFrr2XL/mdR3yLAXh8joP94+7vwBLbW/uM2nFOjKdAt720Batod1HD6cunrP6iCRlH
nc8G1FOWNvbiw9PkPC/SGqkWnYyZRowSigXndsWplRLj8yoWbmH6OqvgvP4KJehcYZZtl62dU6u9
lsp46z1x7c3KjMRG2xHPR1VBIemKaoULFgG+LRarp/eHhMsqeL682z8/lggCsMZyrEEVnF5KEeGK
Pis3jgFKQOVbYMvoVyqkRFiTAuWUO3LXmNGSZv2CT94cKLrqEfPXW2x2NjIgbcuOQfGSiEUX+O0o
BwG58uzRUvsntrTnybT040B234lUlyZequdfe4vyHVftT0Qxk8YBcAWrX16d0i3gvpHMHc8tNfiq
s/Buz3i7EmajL/kJBeNHJsZy7geaZ13SkwLwyFYxey1ZpjfE9yI+YZJF40Tt/KHZHsouVUbWFO9Z
ExmMPgXIVnVLUE/PMxEK5pLMdW99H7rQ11br62u2gjngCI1hUQQNGCnH32VNYyAualPl3tLNGtqO
XXPIGWYyUcRZigyhdBWO0tcGJoW9fnkMjnIEs/ylPuueiy7lIsPAObsukzgID5mBgyqPBB1Tv+6P
xLxinQpX06xLybqs9uIbIWn7u0ULyXF1IdR4/LFJyKXG0OCMBy75KUfc+7YMXs51gGNItT+aH+O9
jXj1t/3WQGmD9C32YREpFWzOtqupLROyGSvM67LZe5CpPNCM8htI6TmW8PuWWg/TCo2uAmtNU3Mj
JYN8hb2mduNrrRrYSzuA9YuS2Ir0Lwve9FIhBBARwtezqAlLl612lD8+1ZWRDgbt9C+gcASN/3b6
+uMSKdsLtQzzM9besV6bDy69fxiIXKnO4O6WaShI7P5/ZMMJ9qRU0AGUyaB8HKjDngDGa5TrZjqY
K/KzVF4gMPnH2sSh6aznnHkfaiqLSfXXfJN1pf2B5+aMehJ2CtVBLM1T9tDp2V20Toh+6C3ReRoP
Q9+9W+lkSE26Txk1iFyPAWcAyWMfwfiWp6IKcfXuh0ZtLgQNdw8WLSTCUYYFCVH25MUXzFYvG9hZ
/9YBg/4b+N8W1wbutzyEu6iSfEcmSQuUy9U+U2j11GOKy/QTYXb8ZB/GWvKF4kbK8LQOp5A8J5o0
JmuSO3BdScr/MyNTxa25JRljQsKN4mKmjKuKJi8mqRV6HA0cs4Uv6ICGJvVEVXgMmHhLfn1EOTyE
G9YJBBLtmF6HW+P5FSs/zTUYhgHpH7DLMd4BpvUzfAFErrLQM4bRhD5XLFa+JHZOoSzdET0vG5NM
nqK4BGWVAxzT2bfw0Irnh8iZzq/cjr6CeecQDUk7k1cp7GAZHuyOr1p8Gq5bVi8uScb8H25wM+f/
R2N760QTEfQIoBd5p8ogN6Uqop+2MUOPv/s6hMwQ/+hv2fEvxpKi3P2FUIpdHuHoTv2riczCPmj5
JOMaqmBN92bXZGqNEMLAtDxAxjfWbSr1tZGLfUjVVIvBW4wz9O7oOFGxADdRReCAy0zWi02RD64n
W4IhidrhsO2GNYlszmW4skiEwt5w9efb1kSR3Mt9ZAVuT3497XOWY+Ql0cwsmM5FlneDTp65dV0r
8A+X86CX1M3UObQJrsvz7dANsWnAIL9lpbXydH9ma1f3FSt3KqmNILB1Bt6BwAEAzskPzw3iZwhv
qWHSVw++GTvmTcaG6kPjG5r7YhqJdpuZYHszj38Lls39660uNDLUCCA/iUnnHqu3l2oxpw/ay4nU
36bS9xKXP8W3AMdtonEBed+McNEgngCWSESTJjv3XMIRuG+EnG/2Mgtb5gUrgGj3eQcgdcLUUWJ4
JoSwwqow9XThX/5SVXdKOl/6zDlwohdrg6H0wRdvB3GzY55vLirldW7fEXn1844ftwmDTHYCpmS1
VzlstFNXx99cx8vxOGXaGrseY9cu/Un8M4TA2bLcbnKVLrTL9Lh1XNXsH32YmZT+S5D76AVAbsqW
Vnz7TobwIsRXrw5gnjKAUQdI5m9AdIxLFWh5IS+M30Y09uaFZ3j7u9eNFNojy5oMF3Nypcwul0PB
73elPOdj+TrNtiS4IY9gz8HF+yGaGbtqFkRS0IdCVF8WXsghsxb07TVuASCoYjBTM29hkfcvL0i9
vGJCfsAcnPYmH9evSb9Rg6+Suqc/ktP/KGyViQSqDFu7eJVFxbxmI4R5m9iXue6cn8Se3PBe6OGl
4ZX+MyUMGA3msuCiSLoXeX9gTlYIKt3WwquBDnx25dGVJpOjNAymUBvp57bcvS86F/PtClZkWlOL
4Gpw8btasvunOx9eTKHu2GGHmVgnFkHsJihhzeh3D0kjxHP9PAR3zm/fjLs+Z0jC39sCiBcx+Xff
pUGPtLAAEygO+zW5ZBmytaaoj9b7UfiqrnbMpPs86+O7IMoRf3bzT64TYt6w+3j3Zsyr1NzwgqKf
GgWlBybP05wsvrFWpXhK/Yaq2ZilvhNwTD7eTSd2K+iEbn8bfDaJiikc7QPOmhUdqYKMe7Bl1Jyy
6c++Dey9AfAYVSAHnN2UkY3NJZnTBFnRWtjVE+JWoMS6sb0yvA0JudFjWeQfJn+HsPuIayestoQE
KvMQ1jx4+y0eNe/jkAjq/zojnv74Kqi1t6SmzUYMYHNqHLd9dtF2VQzj4ZzkPfRAXB5D1PVGEaxg
pQW8FK3Sp3XTfKZrhq8zjbShPO8vR0VWUJXzDP5mpcNMWFDvtfIJ8iQB6jB64fMq7Simj1yMWLJ8
QtAi2e1w0HgXSukwmgk8OpNcepNuv+Bjp91IOl5gWV7vHsepbuCzUQOShmnQDGOwzsXeQPblriNk
eLiZEgFS34W8/4Zg9kAp08KBjeB/FRHIxY/h1zbzjGUSkkELs/vWJnNgGJ22R7XSu1ZKoT7K+9Ti
IYXKiwnEc1olct3qrwSZCphhYFF0OSMiFsCEKJy51HvV0+5YNa1jTDbu0XQQUr1FAwlX0VaLUKCB
zoW/sYbwHcVhfEgEoifmJX6hnTEmUUu6ODnvtmHCBLnXosoOafqiQgy096HcUWbVX4GST+K1nqbU
cIjzf2XddldrzzX070f5HxZS9zRe3onyaBfhCFUz8Pc4rkjNFI+qyL29TywKGATJDmHc4VjN42Kq
CoOna2b6lKcwnTfEtwuQ6QDBz5SaNCRR38QAnE0/bgW4/mcQQN6nSi5AM7muASf1iwk+8BYhhduf
/MiZc/o7pHG+0x/+ximMm8CuWMwmkUKaziluX5sEA5xyA7yVPBlSCHFYUNTu0wcLA9ftXQrRiAVT
4dqk9UrmZMC8EXgQslUxe+RlaknzUHySOUaSsfKCVcjMLZdk2Rr/YiIBOknmtWgU107WDymsmz/T
F+aQUFGYfwZo9KZ4fdehmOv159jxvvUauUCBAGxhFEREFWTJD3mzMX1Zv20ho87g8jRKd+E7Y4a9
m7emL7fJ8LAUaHWk7H8ZJbzIFDcurduGfhnLN6thl9TN6OzvbWDpNlBETzKd+A3HkulKwGqmtA3g
UCo0Poj9HOumjEjdkbYnC7cjXXjhvwxAzWAntELd2huCTPKxWTGMiQ2rAa0KoZh6iwSGly+aGWLh
2tB236qdmjVjwUYAtUpMPJIXCd0wV9BDiV4n+NZpNOfj1BIQxxIp4TcF8MGY9ndydOkrpJ87Jupy
lPvkaiLtUHBL1pAGhM8vnSvz35h3ufBobKNheL0wW5R3hNo1r1QATug6h1QSWbMAj1DqSfAP3tDv
fD5tH11cgVdHbwP5qlqxWvzFtLk3NTUDxzPkmrkKdzE8lTE7ReYd+a8Zk/cPJwdTEhPfiItsAffK
U2gStB5Q0KXEFLrJqcLnjNwLk2Xf4+898kWmMBlwdDP4TdWqh2YlPnFd1Mp9HyQi7bNE4bxo4J7v
mNMMytExFMj513DGA7j7knMY8Z7SvBngpaY3scn3nmVHN74afH2b/AVOAfPjeQhJbflBf0GIT0xx
f25PvojxRfY8rfzlUJj+1xkXUEa99rRNLoFgyg51d/Df7YtSQelvi4Q8T3vBggO2MpNRCbCdRqR+
b1awrbzphJQ9XZnFHlcFB6H2+k+5OOGLy5ubeDuu66NIh6+b/VoydN4HqHiVR1imXjogDv4TviI4
NPPMHPH0I4jWB0sK0CgQEnSSdrB3NpKDsjt4SmM6cs4R1wm15CWWRfCbA05tNAXdqk3PfXnWhQlA
OXG6fMbwzZiTWepGuIaeKGVdUny9dZkfehecTwdhG+l+6E7Ki7jYHVvrU3J2wehaB16pZIaPNC1s
gfd+ULk4uoCYOo1R4sRKFA/3aVVu9VuJ36YA5aKnN1suiVb8dBkhX4fSlAOdgnYN1LvY1I5ythua
3QFFMfSkPrDWluf8Y3v9gWes15QRVkMS4wFaD6bSdvYKZ1u6sUAH3oTiVVPYl4jKg6JIqekBnt3B
RJOHRTVhDCN4n5xYtjur/oJJCtUgxHlNOyjiKQROD/bL9zIEDCVWINyg0E1LLUAPtBUgMgs8x9PV
kXU+Aco10DDFn8VmvQa+j6t8qEaWMMTjzh6D3Le8C3OYdZ/BigxZpF5seCgVuzQTamuWmoQEspeQ
pXR5ZxYTw+LoaNMdf0YVTQLtlYHWfAGWQRmm8sr/+QgnW6YKzbkp15dCxRIVk0Sb5NNfiRJ0w8q9
3sGgHzC2kS2s94bjq+BmmO+8TACfMA2Xq2qjoFLvWw66cWk1nmFUgxT0H/Oezoto82uLmb9c/TG6
8Z67tTtLLwOctgkAYBz6J7IrmrMWIDpEbMaq/tZl6IkROuU+8Z8R8kMuNaxDGIcL2X+bytU7kiJs
A+So5IshdB+B2Iou+qpigdk5W2dBZVqKxqTO0pDwNunK4KUMxFwmzQnYm+mg/nimCBRYt4/hSJoB
WdeUgpFxKrW1FL+v+zsm5LaTcERRGNDgJzh1crVb+HpHrUosEEEC+KQTg5zmf1KlSqpKnl6aIZQ3
FCKgjmklFqfX+aL8FN15NB/pqQ9iluSQBXtb50EhpisNHhIwbBCywhDlJT0YVYykdm9JVfr29Trm
wPDlkzcC8UtT3eVeNQniGjDh6r8MxD3elb7gHYdYeidWeZ9LEXQUCggczq+IeHBSO0+RckUjoNrz
K02mB12eFNcWjYc25DzbV6W0t8u4u7FbMc5BvAetrcoDbVKJiR/qYYtCEK6URyrKYtwpplKRI0uJ
JiRY3UBMV3+Kc1gWMoLU6WN7zm/Ywn9De8DyVl+pIUgXxcbMeFHkj3I5tJVRsF0dvCl/wXjod9LJ
CrBuJtRDob71LA8UFMEk9ELIF1OONEU3dnIqN9ampS1tmVFCnj+ZJIaiFkHrmQurAHW4y5Ems7B1
FCiqws1Xjz1IfDOVyeZXa3abjpTnlJZrqd3ApiJZHlocYDM10mnLY/I9zwPnzaVlCDV79oV31MvH
hYXbvYEJAg49HZX9kSpfbWUKSsRWmqP6ntYZMLsvCX4bRgQTLLOREzbbt786tHWic8q24tPs6qPM
rX/d6pYwE9fjAZ9hRIMBr09QDUo7uAXV02ef0Ys9QqGaLe4jXQrOZTWL0vC++kU2xmsJ4VWgrsOW
YslbQNW3KuPpwbaay2qn40atCOf1dOeNaEYdExTUtBa/wVjab/vHYOTvWFEWrpTjIUz/jVDM+V7Z
qVrNNf5s0W5+FILbC2OQUQEq768Sv+vWQzc5fyM1COAQU9Cc0KFe1rjMfCMYEH5kv2WFbQBanWr4
AYzTyFCXn5idO5J+yh940xe1kwuQA0sv4dCR6o/tLTHK8R1gvUhZkHex9hMLRoZdGrg1lJPP22Og
l+9Z5krd9rvIhlxa2yoYl9ppEPVhyR+ceUc55Db1PEuj9INCfFeSFEWcYQ8QVChtAo2yIY6Bh7aj
Kw9m3w/4HeJRm9HkLZg0wi6pUaXyDoEvnaoLfeseXgL26gkOJHJ7U2qrC9ltpMFfCd89UOUBDxEu
+5V5ghAudUrlePeq2RB/UCOAnomJL/l7uD8S7IVj+hlG+n0VER/fJO+Ps6GwyZck/IxJrskKmOTH
wm2zGAzLY7v77M+jNfdVL5cNcrZgTyS0fcf19IgiU2sBFcGGl9ck0kOfXwDl7JLt4s9WxECm5bhU
dp17300fvxmA9ncxlifXfei2KQ8lniCKCTbRBsESPtR4JoYD+P6/iMHm7z722kuyh7usCVS204pe
zXSjMOzi9Ne/0l711Pmawxd1O1rTcZ9JbW6HV0nuGJYtaxFfywoUHawUHniuwwvMbiIWbZn+nrtV
vGOyT8TbjvwZ211YSP42HSOYXaVJEhRHVcJ6982jZ/DeBjCVPWAcaT2T3I55wFvF/XxO9U1Urr/J
Y1At8C4HCon+Djrdb58MQjumSlCceF+jP11orP9ZH+7V1PbTjTdiTMnrHcraSdOu0i+AFLBXAY7o
PXADrbidq48SJLflhdqDdWK2vmuFjvgLvMSxW0ed1K6keZePuC6A9MpEaEjjWG5R0J9TbE7mhrQK
1rcEdPlVhBy5wWfvzReyTe41HQng44asTD+DXsSdNUOZnx58oFhx2VRYfSc+5/BRMnEG78Cm1Bon
gsDs8bhbUQzQ8pRLj2fiKkCGJ23n7It8OGL4wfg8P0UgpoNCgs/RL1KAxqbUeGPKxKKGWKpLRYHu
+MIiHIPI7AxcAOjt5Ecs6zlBP2HWKfIdHooNBvNicK8PkSu4Yi1bM5VSZ6qF2gmpSrxK2ZNkKX1n
HTa2W0ip4MlFAUr4ZqxQ+oOdqvCv9ri7vGntZy5iiecigR9GfSPbBwpuPLQdhNY1eLruFRC5rCtW
MbNLByp5AcBdCIS62tHZTX4D1FtbuC10OAkV9rFmXdUfUTbv7Gzr8MqdmJWV3Bl7vP/oeBjcF+16
2vwrjrXOFh+4sjrCLONxwgVga9YK/Uw2jMeDpr8rfKAeoydwB80ewCZLhztWvpkG6wFHQIQFkkVc
KJU5Rbg/adgOlrFuuw7KGUbGfvjN0o1hycPozrP222Fc0p2sdBN+tOgr4WIA1bziVonxtrzOWih/
Sd0vio44slWU0uuTCxsiIItx+R4FkNiJTAGzqhBIQTAjLBtBZArQk3NLyXptN9UKkohPce26lJiQ
RPx35NE5lNDGrfxoYgrY2on01+Y45TNXPWGGqVykBVtxoCu4y2Aw4XUqgiVg/WpKqfgUzksmNnVz
p+Fz9trH58qfhX75yiKxdLgoI9RMMXKPqSbQHEcTv9MkI1cHTIynKe5APBrdxiNiQWBEGxxzu0I3
FfNpUn+qHxZ5hfaok+T5YGs9FAFqj7hAXLN62WYEfZuemZLuZ1Qq8KVkHZDnk1RBQEH1fqonGain
ONXqQ0nVTVXH9Nh6Ca4dvdQKLN8UG7ajyFiuTyC9dNKog3b4diYj88QeHrq+qMkrA26XiZ/3K5cU
q20swn/tDByrCh+2YCO/nv8RFUD5zwCaDmS1c+Pp0LavkKzQftltXlgy8pZYO1vSh7XMG6jnJDZI
gdpewoXTGPK2UFu/3Fqcmd6QZSgZeN8TVr9fmBT1qCLNRsrPa7clmLqM0906CTbo/OIkk7p7ALla
WVEIOcKFjkP2O9cwnlvOt+H1VuqeyXBSmGw4dM6+cKNxdibYUqJs7z/96kb5K9y+DYV5VTaI2dRU
GKftT2ld1JMnNRgCfLDK5yyRVbfAycIHlZjebqv7Rxzre60lURcHwBMXhhOfRv9ccHuo943IBwmH
MGY8D2oHumTiiK5aYz0Dcc5WqIq/24Tkv+bAK7Y4ZlJsLaU45Yc9os3dE2FZqLdgDbQ6hpBmFshL
vSeyXSRLNyUKK6l3YKsbuoYcQniyUEhceEkYoNJORoYOP933KDoAYk1yDz4FqC/yCgqNU5YETuD4
QD5fqu1J7EvanTC5DpN9dycIM+2BWZhtZNvzvOgnAFSObOgCuiLGniu4+Kl20kWQt+nDD2lUyVgC
LsQzx9VcIXWoEBzIvg3Pb6t8nnKjt8YxjpoHUgduE+UTUiN/lVK7aYREkAJIp9Sy1puYLTFNYkz0
tujyhvfUwklb2a8HJXIGDcEbz6LOJ/gpJVbE/OTM3hxYrcu62twlN9A515qggX219E6MF6jua6sS
GeOs/T0WUOz+z8UYUvjiovtKswoi2UJfQOyeB77fdndeOAq9rVTwBtJ1LaoTVgH/KUcaC9RZCopY
AwEnAYtWihHIMf/bZiIiluWVlPLqoeoHLiTZpqP1IDGAjJY0Da4nmBd+4/W8YiTqqvY/Z7nQofnP
iVOJ4DJgAjC+yMeclXtsriGVZlATVw/B59WiD7id2ex+w3HLdby3lryU4XCDXRI7NbOJnpbBWSR6
h8EoAEiKmbX7AWsMOMkZ7UkSmdazDq2TwMCGrymZkHlD9zlcocCgs0tID1sNsvgSogKCrJKuTG+P
0R/ZkfSOU14wal4gU1AW9JRhHOP2LEAhtFcTrPc2zhfl6v/BUat+jETEpuVqc3Xx1UHgLHc8aGjD
U3BCjPI9WVDRxLtvN5eOsLEhLSp5hvdT8VKB9CK6nMA0C+DfXTZLZ7HoEApqvT3nmUY8yB5HwyYh
nwhpjMEcRTLopBpX0LngS90dCv8EmMfQ+7Cyk3CK230m9cGy0CC5G229/p5+Vo+T7+Nu4m+8oRJP
CwNtC3qeTmKEM4v4uj2yvjCpicQUqC0B4u1aYsREkIE6EFFyDdDnRidi/utXMuKP77LbKDoY5ChE
2sF960EMXIFb9GPX30lBZ5qQ3eYLv11wY/ceBXOfy97BBuuEeuozbpvoJnLfdTaa06lvyBtyvs+t
tr/TcwbL1+T8fbVezRm/893J0ixIUVK+Zew7gopgEQYxdbYJlZZ3HjGg/AazLL9d7BAlHZftlQkN
+DrBxA1pOq0gF9oF+AikEY3UNvWLGDpJWEVZsbxHoLEfMYVjcRFdaF5HfefC5fpy48wlWN7GhbFa
Adf0IrImT1Slaxrq2RqNZkCk3rP3bSziMGFKviLvxI3JrZYpRg2VW1VVQQI0jXy6dK4T074//+U5
0Gw2op7Rr2CUSLCBSEQ9EjFzTpZE6fSdBASBosNo5uTUp2IpUWj2lNh+l9WVKbsnKN5pHMDYnkm5
PF/392RsUYbTK+AZd2HQVPT0cYZ+rLq3kOp0qq7Dro5FWwBIL7uzARB+M5Y2Vv4K9BsYoZppbqEg
wJ5gd2mDzFf4N22/d9lpFjW5BtL5MzjqxWWvCt58ky0jIxFZnALo5RG3WyKtMLoDk4v5FRoNKPbC
BvNnsbHyfJdJj12UQsf9zoc+Jb4GS3aG/iMHauGcLxZAvuDAO7wLXMJgPodTnUAc3fBMH9h+p1WO
yR6hlGASelly52E1ieJzlWUWlcOEFYiq3Kebn507BR6BT1yJRr6ySfID9sXK+mBeph6j6oWDRclE
F5rWSlZK+I2iIJCGj2Sd/3FKGDaCCQXAKjKnYN1cFPBxb+sKOwntr12LK2iylhcd/t/UgkJ/5tqh
7L96OqvI7o8nkum0w4JcIO1sVPaytLSdRmaJ4R8AC8Pyhd478OgcSr2GbS1fuCCzazCWjvGVmoFy
4hcr2HeZRtnBnXVeSWA32FaY0usN4lZDuv25+FeqoRpecf62w+Dx45O6oTQ+getwjr+7MIjL3/ZQ
X1/gahv6MDPC8YWg0gsJVRroElLnMw21hmberKuNqDqOyszqkv79vi9IWY8hZtGHCoKTpA0evgI1
U7uzqb5CDoqiU58boouzGzMlNQwePsHmMUetRLztImjqM+jKTJRN5ZoYmEvCZ2L8LbRc+hB4Zyhx
E/BvBG6rcnJzwFqKiLRKkBo7ipLBMrMFlY+Zm1SVtHbvcOU3URT8RWimcfo7mnEQvBkWAXqrMAU2
fMgKWh22K92w4N4Tnqa2p2JX7VWayUpmtiwCleqPEsmNzSWF2F1bJY8bg7MpVjjs6ff9isMsdk85
ZhOS1TSZyUevViyr1/4BUgYIviXvmOU7Sje9RISinxEZfvsozesfj9wtgLYn5SE1/hQDO7c19UOu
YShOfkp2B7Fz4EI1U3n0t58ZN1l3jlgsRPCwKOroTpCNonNjxoQkKqZPlW41zIw5bULhLIM8JCTS
LHuKwUQN4ZgHBokGbAYrEY5WKWsNxpW+M6hEDJGYw+RXt/qq02zLJ5u5jf9+AH6Ct/QOrErpSqeL
y3ho7rJdaGgebnSeaMEFlQWnDHZAiQTsDhPoN5cH8UzICqvvNMI2K6i2MO6QPkDRvwxlAnnH5kLd
yVpFGEar+WbiRP6vW8IPtO9enfhyoKCuq4NpeD5cfvtios4EBDIV1scVMeB/n6hJnQDV4+Ex1gZ/
Z1rbWpPIClwVBzOdMk8hXS337FWUgxtpsGVqdadTVhsZPf9qFwf6pidAGmLaBX+zg0kLYU8HuHu5
Y0bEqjE+b9k3L1Mt/EXkp+x5ubJdvMq1sH/BxbHI2jJozb8SxRximc6LRSJQnU+evGIqJwpR5aDb
zraGDHZQ3sBfZ4VF9qb4rhvxl4rRuARL9SqMpVq9hqPflEIQgzp6oO3OMOJ4229x/FnIWuCNx/jq
nJ70/jZxMZ/x4ZyQOJ9F8yc2V9OccX9bP9EqCZ5suvRzi09evN6oA/wPfn28jdDBKNYKI4st4XN7
nrgzeGUoquDJQwBkg6C9eY8zuXF7zvFwnuhXu1jUQuOowRx9NvyNXFjos7hEc7iWJ6LKn2UOZpln
X+s3DlRTYNtx2OQLtAvu11YYdksT05yv6kUbj+3NE78e9ug4VPqd4UNX98K+Y8uuzKQuksYjQJQw
mlBAlmtsaEWO3TpP/4+T4+zDIITJpio7Cz9MXBzE96mHZ/9PPju2wjWqxYGn39ppu/28NhsDuUjY
Mt7K9zOZZABCrYd92i5CW8Nd/x8BKwa4L/9NkxtfLPbDiZqewTM+iRuLM08XBSVdE7DtzySg9HG6
IM3pXelqniBeiLKaXnERzCp8GEzumDNxZ/phCDTSNCPhRKyH/geB5wItX/o+hm/r4VypfptP14h5
v8kXljhWQY1pG34spTGM+sbr2bJC3zbC/Lb09gk9Z2wUYd1RGn8tOMA6d17GhuvM2VYZiH3a7C6a
xqDNHItRsjimIKiMhl27tTwQg45ra/806v7mGINJxtHQiI2oMYF3mxgQj2k+ovsxmBGiJpEsAZnD
5kDvSXI9r8eoeCBK5Z5+0nR77MFIKZIG1pk4HKysVV/hYR+8wKuw70KQlijp6WeXW7wNPMs4VFPE
PA8Tcdd2Crd7Y9RS3oesLunWlTsL6kl2WRLO8UwBkGfWl9QJv4RnD6tVAKY/LXCtxQomMiKS1ELL
SRhFLM+Vew1xLbEc5ml0OaF5TTprkBApHVkl+VONL+hl2SeRZfX2rIydUiwuVc6GrJOe1y9T/hBm
qpQU2JO/PnooR8L2L2eDobV7fEMn+30C8SNranm1MOEWRMax9xDkHSvC/u2n6bhGMmTVaf7Umr1Q
EUamOpKPxPlZj6pdLuNd0zciegBNoI6gYXvXvrzTLqGOlOeOBrmZRSxVBm57bB65aAFd4nH7Z6/Z
BhjVXfIfyYLwJptNcn7Q25vG2U/hSQ57WSKfIceDuFc2HhTT1sqj0iZ2HJUIJJHpIzwPaY5Az5hS
s1C/nT5K/XvRNlxOQHFu62QwUVfqFif5WeNmdjMmsm+59i4zY/P0Wm7TiSMjQCJmggaDo1BEvP06
qkoXVusXxE2C1PwFgOims51qmvIAxHa4Bbu02mKiuyBzG20aF6EuTIR6qW6ZcfaA+WlP3kI5Bc+h
1JGt6amxbYcYKmVnlCdRiQBZ2Gynhdk3g1u0vCt90poYB+zJNA1ircOy5iRlb29lRdf0GYmaao7l
bcgz9lDldFR4xrnbkG2LBUXq1pZ1LX7OjWvkIPynkIXQgsILy8f1MOF0YKfH1i03qeM9d0PQjHm3
xg1VDGEfa9NqNT/jWA5N4gLIKVE1UPdnxV6p/jZHZZBm0lZDA/wiBwtL8HXNZ9GWARASbioKE1TJ
O2kRwdBslZ4h+WzFGMWklyUPewXAQ1HEoXulzPMr8o+2Qvv4ra7VkZDE2T+nRse6nASjbp/SSMSw
w1DUdqB3yKOnGk7rNDrGcBrrtSJ49qfriCijrduHd7CiOwvh3JOipZoS/oPEm6qBkcBAb5ofFBDG
TNxTJUDRKVPZ0H6HJbG2+tDOh+mYIFcIphI4xpElGqfel1zxGCKLb+REwOvrNRFu8Bbervaslb8x
7GC4iMMx7dFrmtjBT2V7rV90K/jp5AyD0CyA3h9sH5J8mzgI3eoMYfshkxcCW/EmK2mROEE82v7y
6q1jpFuvqsBdDamuNICfvzvue3ZWm5pDX/XNahHV3uzrwxeUzbMJrbHnC1mIfku6H36Az0xi0mEB
amMEa7CNv9ZlJEV38lrlpgJFnclUoT8dgJoCjsKeGt2ukD7He3Are8NJOaRT4OOjyy4wD13Qq8dX
2iraAs+GoFqBs3Q5X1UZpBPoS5LJYSrJ448F52wZPtXKg6SelyYkl40VtC/+gZD/BD8wyQpGYdKu
Erga1SRE6HP1A2gf7Bs+mERQVAD4uUr4HougGPUGf7LZD1J1b+b+FHCQC6VVR3tu0isNojGZu7W8
CGgdrENX0MF6FMazU6UwsTXj/rt4qwsOqK9XlMWbu1z6+CpHpbCZVzVkB0iTLr+nsNr7MzrWabVX
nZuwP2Z6ImZZzsaykIvynLVXgmqLPMDsCLD/7X7d9atoHTgcxG9Y0K/84KD6y3SQwoPMKkuBfYmV
IA2JQsHG5MFPp9WDaVjBQtJmqnf1+kgkK6DiDyMQnYLc9L4Bybfxpohuncy5tWPhkqmuPKt03jOm
1nAoTbaMmpp2J8OHktVKRD7UklIZZWN/tL+kqGrBNEhkzXmQsv5/cgjvqMoLrl7tUuudyf9QNPn+
wiLIp3EjH2wJk9Sp74naFmuwjmD1ac8uEluD13g6BMc1mLz/XgbxeihBW2uhVdU0hmCulFqrdf1D
oOAWV/92Xh6CcFKiRcoAcfSF+Bg/uLDmLwr4Eixg/Bv2DHbn70PCs67Zhw5F8Ek/mKToC6O0mHfs
pIgbwWfFZmT2LomOKImq96oCo/s1C/bnf/bWDp9Q3VF1HyaCPJT9riufEg56kvfly6nD+gztvpry
5C3BBZsh0jKsyeKS0TiNXVZ79jTqqtjrBo3xWTbm9zN8udo9ghDrXetm8l9zVFrr/Ij1yoHu/TnW
xAAxrAjo61hfnfEgvZeMjcAskCoUjh+I9y+PPXSqlQnnTbL/zVnTIk73UgKwicdQll3oaWd78i98
pbsgIBTD+8UehGYvBabl9orSBladDJ9m9tsv78jvtEn4ZNmljf30Gu8G4xw+TJrH/koeN/MTBYrJ
CHAGNCwrT4h69QB3klTooASWkeGvQXCbl3PcQu3b7X6BwEkFzpzvxwMnSqmJ23qTfVB0NCUfc+jV
xsUF+yZSfxAjRMmHmNCfqt6uqtLmer0YBTcFIJCAaYCP8QYlh1VfWhM5J1Ces/aJcQJirXUpqpCq
yPgXqXTL31yo1aJM85xJ2utzOCbrHpCXgcgOd+t9R9KfBy2TdxfLIZ9HaoT+0bMcFdW6XzTJFvo4
nV65dezigPPrlRaRBg1hvvBrp/YGpatZahQ0Zct9sHy76LAQVjl6sNQCGzyOE90euwHMqfe3ap2z
nx81aqbjtrEQcH6PcGfBweDSByvtL+tKh4tuONo/BJJoKu9ltfnZWFGt23PvHNghROZd14bk5XkP
QfG+qfQQMaRlFCda1PypBvd6qHH45jGMtqHFV4q4jFPqkLVmKdrSgUzvUW3OogfPS0UuMXSFZN2O
+IB99KzY7q59fk9TJCMpgvL4rSRX7KoCdaogGNwDIQ3hDs66xIhwGS0UBBN7NleRnZ4xmJT/f+4A
/Q1OLe8ZkiXiXNGqC92rbhr8eC8JzAjNlFhO/L7lgzrkTJDGLRhxC+IPbzR74ynNSZS1FgVTa6Fr
zC4i3MInnUyn/NIxIax06B5wKB/t38nxSh41LSzdk76DPLjztu31z/ye3RWntb1+xgz/bk7PmLmM
pwuDn/k66u05roYo+pvbhfd5lXv9EPEQSHuUAJoJBJAxorkxTJMfr/eNOshqD5JHRHclnWU5T1MQ
z5Kvh1pClbn5L7tdW2b4Re6Xf50XdHOMQsA9YA27Lv0/DMKtql46Uf75DVUuxd9mVWeXTNJUoCQP
lsmxqPxXvQTVgJKYhgDg3ByZr2R7YzivOMRWNNgGuyGJIpi1q3mu/EM/uZmTX7UHnTyx0TC1KGHI
QMjwF1XhamlNgAzUHz0BdD65FcsNbTNKxZNtmcxRNf0HWxQq/RAhZHKC6/4Gbf4hi6/RdKBkB6kK
GqqI2LVKQc1KEiBf1buChZbbFeSRxAQdmp1ruzFJvo0fWDop8n0Zw+bVlTaadKnNY6EXhn4EUnhi
7G09QdtRHJiA+rMoZBHV67PDcXxrIBeOSngP6SvUuP1FK6umFTqoxoSoDx3qDyrJdFuOi26dPCUB
YHnjEtopLRrRp9F097S+j1C64WkgPfVVkbxgdYZGNKaev2AzKq6mRVPlvJ+Z9k8dLXkEm348+Bv/
LCqtDsjlwhvgixAO2PCTzOp/gRnukggnlFI/GrPFq4SRuzdhXAB14r7RllDqzFWTt99TSRLhxTtk
9TPSqzNhFEY34HBgNCIGM30SwFYlLAXRm7Qq8BfXf2kY92Fo0XqlQ+wEyqEqbdVzCRzYmjh7SfrM
KJi95fxtL/Ac7mR09vbnFN1KMn6N5uZScUW777+B2dUEQxkLv2nvoXvh0NsGFRIuo3n258Nsjx8K
FSySDaCmGsIZSl4fcOs3ihprpSS+9vknBUKa4RYhNlPKISEGv67e03vzCCpV6CbDokKRJt7YiRHw
gwlv7RuI4+e8bcX4NmiRS9VLu+XV89eMFxDEx/wCrb5dpyYRI1LQAhn+PhkBWDNL2sw+Sg47wCYM
tkEQDQYNqwcgotEyIUKN2BLb7bSc4EYDPDsOREMDwqUf3VUAuVXFoIPikz4OywVXho15UdtlVrDT
ycJ/+Nk2qwGoT/tuRYTIarENMdKzXcCQxt8uTuyG881RZKUupS/rik+wJWBXXSxLXCbzSjDWW32m
PxIXt6DZu6EDVnyrcs9EvTLnyBgV3KXYLg/2sjdj+zphfOxeVRjGl4bbzYyzhZOzsJhpSNr/Nucw
oPq82KbciyxBy+90j9tgu97XnTqSn088cIJNntyvcGwAJKy3tvUlgdgB0O9EALCWtVSWVkJMf2Py
Tx/Qdjfb3+/jRmvNM6XqEq5YLoJPfjpBzTv4yxjRjVL+Sat19viv0jGCZXFtAz7/1GNkJzpuPJEw
GlnhykuySqIDy8vDuKexvxdnV0LRBBK4L9Bvp91pht3tcbnLjbXq0IAw76PovdMFonp2PVkYK1W8
cuh9BC8zhqLR1pCcdTsi3X5s/D9Qusrzc6fJhncXOkLnkpCAbNskO+4zn24D74/VdV/jszgzG7f/
DleSQpABSho51Qdve6b9VBp1VfHMPMZuzujrnbkE0d3rrgJUrJpF6yzF2DlipUEFy3XqvCfEaBIz
0CCYgyctRVdAo9AXpj/Fq2g+fg+EGq6+hNJpQp7Tcrjo1z6U2KMUMUcMuLBelCLvqgmB49k0u/hO
WsOoZip1YIL43HLqnbc/k7A6Yacs63xBQ/EE9b42vRgsWkP0Y6AmkvYV72HS285YmF/4dRtGni/r
52eX8o5MBtDfns1JnUsKRuqthKF58Fa9LQYYtb67VLS5dNHpjIbF2zK3BuOwLInBamxZO82d0uUf
CGjmNp/AU6t5P4IrJROLxQ3Hif0sjJM65Evnw6heO6q0ae38xUf50icXNwo4L8WS/B+Eg5tAI4ls
rdoVV2mPF1EIpNS3f2LpCv71IqIy2Y+/V1p6knf5rZ5t2ChUYSdLc4PobMV34BC+VbPhmR2nJ94P
FI2kee2mKqSb5TzBKPw0IlA1HJRFdhqKZ85yHRGlxaK7ypREYy1/9foNHqz1iSf1XuhhE5N4XvVu
1EinZmzjs5Ib5C89C5jGn6dBCZnx6fShxSakWxeSUSmSIUKAssTzHXlrZxSjcWMyasnYUjo0fjYT
cASNrk77vufKovtiFbAhPIjG6g2Bwo7jtjfeEbFBWSXeNR6npkbwV8mMGZeOG4PHm1Ci3UBdDgcj
Yi1a/eBsXZhFA80TbITKVdG+I6hUpZFBOXJztTIBpq8qwidM31g9JVMwE7vHt87/oPac78mBCfI3
hsLUHSLno69Nv55qJ7YvSAHrJm2FiqNKD0lP3WgTJ4EV4uFHr0t1axl2Gr4iRwdFf7h9bTgDO9gP
wgtMAHF3AgR6jJK3MaynjnHmXhE0gnFotBNSXadPJcQ2IuGDMZbaAn/xQqo24RK8Vbo/Ch+8tWBV
kVyEwQCIVs7oFH0zUSZ4gIhbufrj6TLim9wMuYI/bvYfVlnGd3ZRzTmZfTVZoMx3T27ZRI6rdtlR
8siU7p3Q9cq9WcrkJUpoOE5FPlvedLgXkQrtaFQLUlK8hrzgFiFLkr0zv9OP0G73mZHvCeTDwndM
OE+hWKdkLj10kGrVJ+dDQaEuTXSrqKb0FYbyWgzxHDo4o2xvvYnUE9MXKMhIPVu42knyZ5O1jGDB
ArdcpH9obShZZ/WLy6KyQ+NguhGFt4/3nYCD6K6vidBL8KdD/KT1TBKkopjDy04B+fOCnGfENEKC
MkvPCuqsBwEF16rWbRCvQ7DUHyDhHCFE73qssc2gnkk0xbDkJp/3Lf7IQobRunz13vc95yy2tASu
/2Thsaqo6Eg6xuiE73WQjo7gQP0Xn0cvP0ZSr3si8/9MDa8Ei02L9sImpQJTuuF+PLAN7Ll/F94W
9T1draQFwV5K6bbzoh3moQZ+LTCbRiNhNvz4OWOzpI8LP/RohoTYP4PEzD1XW2Rsz162N9yeJtDj
dnKXUneFYqeGFBJbKMFwYvQEcMEpEe69qjocPCCTEXMS+uTyuoIk1sVcsQh/X2iFUPIchBALqER7
eafOFbWRrR46is+BytZxYDlFLCwtI9q6U25PzShbFF2psXLsa5zZw0f5RCkAunowQ82g/xofrrjb
W4J6PdsxeaUAzV9wCwId9Tag9C+sZB/T6ULucqFAW0NVLSplPuSAICpM9wglh7ZXdZAXFPX9Xr07
6X+RwyMRI2lLd620dNbig51vrdO/iygDGnUmP4UAPs3SEO3Tq8wqa0iqw1ACueLO3cZn3SZZl0si
VBHBEonfl5p2rqwbLnMwwDKDeKYKVYhg4/MJ6maCkBfQrOBjT8nMZTjkObT4KPNsPDARww0AVAVU
pEXVBjXFHqXoEaqzuc3tMjBujDIiIPYWg0ywTeej23dFyfVKN5+Qp1BZ/w03uL4JW3t7eF8m0fUa
ngAzkDCHcujajrFSTCYQu3PXhlb5QnQykkrWug6JXEozLOwi2W1reCtkvHLGkP6yDTND9t7+IqOd
lmdtOwDoJQzV3fA89fXPX7lDnjvOGbDPyh8yyInww0NM5r9mE8PS6XFBZRHqyooxNPHvAqC/+zs+
B67LQ4Ag48HkqMPMaDDnE/POAUH4haSAbBJCrPksWnQD/97XBNP4teML0u1wlTIWqSJjNFzS8CcG
Bf/c0iRmesvOq61Ige0+zRe+tyEjPQ71JCioWDcVUzVIv2Li4po1Mox0cdoXZTebSSQyG6a7gMc7
85R+mUlNIs4gguyXQUHb+XHMZQ1xtEMKvJ+Rug5KH8S/StJtFvoRMcdtHQwXPohbgg8BOzqrZYB4
hZHp7YX2gYzFk7/tSwv6rhgoYkBK4PUlGUgTGjkZybvFOV29Lil34f/zxo+pOKAcSM6jSCO7XBgh
b6sa80SLeqWGZzUk5rPM9zwl5yI9yYsCu1mW7CffJsD5NI7ekmXrYzhSespstQe5fvhNPdbtnbmn
MxEfOAxdVoN2mElyz7qQPhpoHEtFJVV808RISDTpoSSNpyxD0wl5YxbhQYwFTZzluv+XLS8QQmlR
KjAX+JdAevryJU4Tc3A6Ws6OErxVG3wv7kZiECr26TOw+8hUXCoRWLi2EB2ftFZdziHwN9C7SEgi
NK1JOa+VcNzbGBl5eYTpxGtcf8U8KAKoyxgk3sP1GEThhOklVyCfnvkMBLXaYt/pwSS/EPIRm7Uy
EoEH3dVpQT3QhMAkljc5DpFyqY3jq8dhAdAZFq5BccO+gv252f9OOekxGWg/mDbFk3/aptDRrcnI
fbJRKWmiTCF5Whwlv/H+MkCddJLXzg6vc+NjvVRWUJ+IRDlx+ITPTY/PtwElmllfdhO3MB+1dhg3
WwPfKoIFtAk88HYAkD/yRkstocBJ54asRgB23xEkj+EyRnfwsuuLV0QgvAe/hGUtUZWkgYJdAnuZ
1qaFMRYC+Sr7Ub++bxXyPADXYSOI1w39SNzJduEfERsPucC6PzSXJa7XZ9b1XjlOUgdbrsORTzO7
UvSbCJX6XGDzVD/gWyUFSo0ozWshDRtxpROx7cuC0lUENCB2c8KGTQMeCPTWW4nPbnBhYDvOzbVE
Rf3kjO86rLR5VQiyY4M+6z2QRAxQ1J4sV2VqVu5K8mOD+BeI98f8mbcaunM3++N4RPx1CrYPbU+Z
oWVf1JO4dV/FaaHE3s3HS5AxiIh/nRQtqsk9HZkEkvy70Yo7Bc29LLKHuyR7LX8ujbuQ7OQvObNs
fCHrsMcr4ClWRoU54k4Dnw0u17gHxCr6shcGwqBJgu980RMzKwGYyonT7d87CRqg1LOCKQN/xjMY
wlljqCzcWfkajbwAz6uXVdgCYHjzh877wynra7DKFRv4WThX8J1w26fpVRuL7l6XWv8ZEEjoDTLn
Vuja8ghFfMdyy+fQk9ip2K0kzxp/s63rpQ5KvIJ3VrJimOI5xtIOYWIjXZKYVdWSlxiu1aOhThyy
OXX+uOp5+wIHNSFUYOyKPlAoKBGU3NPGhiR1kisK4SUIQ0pHMpmVhVd46cWkvdvQLK5xY6dZaeKt
hzY25xCjuY4ZffpDRoX3VYJW9UvkZbYft/DzNar8oFTS9UKSIOa6staNSfwg/Mqxa90JyN2iS0U8
PW4jIaLyS7WYNnMoSPxfM+b8z8lOxZmGLs+1oGa3aPZNLhpaTUjcLLztNagn+H20WouE/D7ITgul
zhEJ72qttHF2+y1C66+PHi9GbZeLY1hECM6XRcCp+R/GSMrrH3gVDmSWiDFZXi7XZH7dF2sW+p+C
yNE+LiwxmVWhEIfY2KkBPoCiZFzKONq403CnNx29Xfs69t2NekhSrqQssRBZIqvLEp1IPjd2jby8
dR22TD/qXAd2VLytAHcnZ8UnoFXT0pTScAv6xmhLs4O52eV/NOgDZQV/SCbE+VlUnL1toLU+hbEQ
bHdvVGjhAA/pL5Dy3NjHn5BfNNHoGydzyum3PKXaeurpMWU3QZmmY9mgocblXRzi7N4IsUuWUp5Y
Wfl7o8ZnxkpUIQu4PIU8TedLOboMsCuFP58AASZGEuUACyY5TJZ5aI5DikESf+jrD3aoZA3CqLmC
/nI8Gin1JMqa6kndemuy5yT6EKYqVT9faMymO0UipQuJWqrKX+SGwcy1EN8U7pPzSYuKZzzHsWzR
v7N8mJFoCl9VPgGvtreIqaLs5sK3NrdDgeq479vKa4LHFPC5oCzLAnmtDl/DcBUbRQWbE/Dytf5K
q+4AWqSPnLgnrSUT2eOuU3M5U2BUVpPZwfFSaYvhw/hnYo1Xc5MUHwKSnTAzTOjO6i+EBeOXlUCO
sZYKVwWPRqSBN4lnHhRnfXHhIH64VIQFEKbCLw9tWo0NhpgK4wC6Zi86d+GauwPk/ACotAtnqt8J
X4Z3rLFREvbW4opLdwaL5uOmEBki6Zk2yXvAJXrO1c9fP/OAwmhc47QUE8UOxXn0scWTTG2XJF6/
+yoaWEngUb4PE0UfLZMEcYK3eqxe4BJ4PlMx0pz5oHabrK8sN3Yhi4MTQcXLJGjexmKol5cKGUsT
rYXAH3C78Ys6l3mtd3zwJEBEtn9Hg/ir7VKEX80c3cdIWlb+TCOCbB6vgR5KkIzsCa4S0f/pG1mD
NZxkVVSTGM7xXRF7G1zkr84hV2UG6LPJN7qApRqe0wyMACnNQzOm5EauZaeo2JR/M/9fCXNiS7e4
N11e+B2zYeo7WIjFaVAAGEBXKKyCevz33+wr4/KPzoUFRKxHWR7VjheSMTw9mwQPB9a9RvYybo+8
WqJhQuso0eaWo/R1trmjNyMNsJP2DNZMGgdSRAWKtIbnE7yM7A6uG2ikAzye/pzb84HdKge3cYyi
8lXXcyglMDM4kvopusRQnWM7oGwisGeFSXTdQTopRZrTllhUiD7gBH8dPhPKUCGW8H8/ajm2pTuA
X3dqC/cx74ITmyiGXQYyGWQFOOpbpxpqE7KkdjD2nphZ2da00q9kCv7un+8idVYAJeIDS3k3+TnW
V5pKaEt2iXUsH0Pr+4zUiFw5y9MgN67A22EtgOyR7r1p4krQ01jPSq0Jbtv//8WqRWmVGL8DSfiq
Wjtoy7pu8i3p/CKdA2WT/Uz/1HHBheVYZVB9k8nkpuMxgtVSseJZPUlJPg7VaRHHfLxujF2KUKYR
KYzPdMtjhcAY63uPxg8QpE1ho9ei6Owhf7dHOABkYEzYbP+NGUEhwiUFmlqaMmNYVBSRKsnZKUtL
t4iVYQBvnF0KAge2KhqevkKImjUhPDkVV3Bxt1kc4fKNoGsq7OUZ/2YTVNHVaqaSK6A7nR7pUT4K
2U0/HJ0Duo2cNQRpNqIXP2TdzN75Tgi8+pWZzLIOEkgYqxzxw8OstWhWhXtKUc4nTgQuE/vR6Bu3
rNf6E6U1LKBnYdw4soak8MYqCUgjLyaovWwTvHrBeXFh+ZUQQpB5WUP2ZcqBWtPAQT0RkbNxa4dU
Ulw+8IWfVzSAvrvlEnYbOR5hASnlKQfrIgQC+J6vdCPab6QnrlpHQSJ5B0RtrD/tHzCaME6Jn4EN
Q6qtfUs5yTvIR6ivQvu1WUdtONR9jBIYR1Qf04KQgKoeqGnjLnO8bzugdeLEh7L0959WTiUawE+J
mqLdmSkQ16cSnAt5vBserUE0ch5ir5wA8xzwIVDl4z0Rl61UpZM3hixGZwDBnV9MWwF996t+2vlf
MTUqd44JwUE9Fs2gBvbYL57Pmad/furgutD/eYW/9DA7BA5Wx/ZjmVFTZ4hABhgaNH45TDbinMYg
Hc+n4J86ehJTJvcJDhkLCFEh/aBl6ljFDdIhBve8WiiOHM+DuY4fQA7haOwNUCV9+JOGTOLHVevT
yDXaSvnAttVBhRrGNMQFHd+FOPKGl+OLSAPGm/ooe5v6+/aDUDOMhSDCkavu8htfbyoVA852PUtm
lbfGTLcY4jmBCdnwGXU2ack6+L7y6MTwGs91veJCUcxRlU0WRGawZFqrEN3JW2uhy40K9SsayANi
ZL9QCtBNNFZth+XejRnTf9raG1fJw0yIW47xK37sp3jPu9n4S7zde/7sHEaTVcqSGWXC6Ed3APX4
oJG3SBy/iAALl2pw/wCXYk0M01UFDSmGIXTmpuNwbJLFXxG7gEDTMHrES1S1lOkOEmZtz+78XcGs
MY3KFPVsOgFHxq0l9S49HV8vTrCEIR7frv+jpfnI2lSP3I0+gCm4j3jMdtHarJfYYjaTRxRbswVJ
TqnxSs6AYkB09GUfptTSxTRPJirBloomy75/Ru2tOVQk/UeUynK9BHHrTr7HFVlqG+5t46shixkg
9ID4mkn8ASlyclL8WPILNqRX/wOqdrAmN52jwCOSdK0ThmBMykms0JJ/z4P+hcxJSsL6f0fMVQpX
0K5TzohQlY3ohGbT5BgLw7kb1yFkl1Dm043YJUsnB108qTOmqZBVhngcFkl4oNoIuxEqvQrxO3yw
ID51PtZakmBAdMhpx7X1Nmax9Z2gbeLL6lqJw8O1TPUi/l7X/xymyDJQbU6vEGLksV+onyQxEi/m
bqgCaOtFX+YkOI9JbDnPofjJ4CRssU0pYS81pYGOUusa9lUnCrzQTyvC4Nqxpggbdm6vub4/r54C
/jyXypXVFzNHZRzAMDwRjqfq2FRMy1XNMmP/VqjVPKFYUPAwla16e3vgnthAKxwnSDr2oCXK53ls
86teCscdmpitlphBRwnfBzDnQqwhixuCPz14CY/yzyK95ZgZvoj387xjftI6v27Dim48nukBvaE7
FgIbHtIIAVhWZ0R87El6Mhro+N1RnwguDjurC0nd5lU4VeUVfTjQCstEnuyi8eZu6fyx069mo4W/
544G57Iv7ssQsM/sZE+FofWCBh4pImGszwkuzEIA/vTAwwlf1M19Gufe505PSsZkY6ubQyEkNkS2
GMGFquYtc/Z5Xi/56I4f4zsncASMXnzJqJpiWovOktccjLh1aVjTWNZVundz/v/yLHqhG0ujd0Gg
wcGAg5LkiRrSWBv77ieXptBihSexK6ZwFgxXo1hUeOIswkNt1sZkFgvyPVeF8KoTeqi8J6V6TeSN
Dy1JHby+CUOOjazOSLLpaFH5PC5SabvOetvRBGQZgmtuCOHQHhafgJCisJz5kYGGztjrvPy1DTKI
zxcio44qaoPyiJEXinjuqSEs6dd38kvtvDoa3+ZEOiulaxO/NK9LZTxfiJ02v17IGhpr3ZXkRE7+
f0HxSDwey/KG2clU4cL4gWkFw6dfiJv65eXsA3J8KYWAkzzckxzBvc85y+GoQ6sdbQ1djQJ+zorf
iURNcm8D76pWrD+HTHp8RZ4mDwdFacnu8D+Fx+LbFdElL28OdSFeVmmXN+QPH+XGR88yNy5I+SEb
4dNb47IGCvc5tQBaUVMPZVaHy82F0rlonvyF5atXT3RFPJe/VpzCPqm0igkzv9dyrwaAI9Jpdc6w
2a7iQlRDzvbRcM46or8v+AVOYsbO7/jKnkJKf4eAL3gwha5aukXo3PBmcrNeHEfl0y4QTzMqDBpW
xC03SUjsKmAmV4OnMjTBX01a/FQZDad3dmTFrxIsUsFaCbPB8BO0GSyOKjKBnJXcM/n/0GPCz1V0
n59vPhr2qPO/RGx53ST/BT9NPuGAwhCJHuHzh/UPu812H8QH0jHWfb+kSbqSZ0rqCu0lSXHmTAj2
136v6qXe47DmBSg+skfkBz94VL8Y6loaqbfW9dW0EBUNOuLx8zezrL6L9mU4hOmONwZuYk/Ycu0/
v/T99I4XoZABt+qiFekI44Yvsj2s81Qbar1vpc8HCBDfIY9xcXW3+nniwzpPqM7YnEwVd9c9XCzz
DJ5OAS8d/6E1QQwZIL+As34/tuuCajT6tHiAt2uFloytr3NWxmXuFXbOK7dHDp+nflqyNt5sDu6d
gJeJyk9I1Lo5mZBNeKlQ4N9kFBkGyVCbfcLBjyYl9nGYy3V21WYy4/ux3ooljTApPf655fBsSgyN
TsI/WrORMZZaJ+uaK2qdh0jSRw6C28qxjnUehiux+4i84wBkt/JcfyPB90kZ23lFBcgPU5XOE4t3
GTEoX5GFJVGeNUwt1JhckH4YkO3L6yez8pixpYKqmZYzNSaFhPil7HcoesIM97a2jF1xgNgQ85oL
M41nlaI21pHw8SrxzlRYYIBPcI7bYJaRNLxcZ7ywaVsgWcfIE/hS5FyRmg3fW56+b3G1mrkXfByq
ke7LNzYt/hXfzRMV2WYVMTBufQKQ6ByWgnzQ2NIL+MVzHAvBeA+NGSTaQdQhBeHbxLk7oiRMQ/fO
2MotIXznwCVPim45Jzxh8rASrRXKOuCSC7cV88URLakPWTFy4nrOcGiq5xzcznpmS4c/G6dwI00z
+skj0T7lJ6zN3qKZLfXuOG/Itt9fJxk210p1s0EfsOxz8jLUa7KTkh2SzeEiFy2K2sCCDDNte+gD
Hw65La6TBF7uYkqe0WA1qemSQ+TuJirkbaCVSQqY3u1FKpUTgFC/jLjoDwpgikL8rS8r71BawH/c
8BrlL1CNL7FyZqTngssRRHJnWaO9bddU5t6YviRnMPU30zNXypg6y5jCBUWb6CXfqaTRE4XiLTsZ
AClgk9gKamgFBe0wZ7UDmNsx+znBkF46G8Eqj80uzdPX8xyiYn/XzWViAEmjdujhN3HmjIYq8TP8
H9RrAiyYH356JVJK5qigHn9SQPm7U+ovL6HjMDRa47s8ZSNZXWiCYCq41f4VQZt9sGrkcYTWiKyK
XpuD1jrrNpQqWj353ZyJR23ejjoft0io1+vNFxgR7VIS8SdEzIT0lWynTXNA0EloBk+PISyIxIWi
87KBuHfb9TSDV84OH+ShqfWz0PyneP9Q0/9DOswPSl4Ul2OoZiCpLKxhyeMHohcY9wK/r10bAF0S
aYojFTjzfhEAFdxsvwnTUSAyQRqpttRS0T84KhkUzOczVO5n/ndmztv0fIa4cGG5+7d0WGC9zxGU
48g+sZielGr0LCfCz38pjWg6DeTpldiQv4DO9XyqmXX4LWGbwa7RHvBT3RfOv/k1KNfB013C7j8q
wHENWHBEMfJvWFE5o946ar8NvVsd55MGcKVBR7ZKMS82XbpSSvd5ZRIAGej2yPKd53/YswvYDYTG
zAkVqAg91qA7LspCqVDc0PoG8CaDLvkDvcS1AgNIyBbDvlQymwNfVqFinmDvxxFHOriSMKNe4buz
b2n6U3HPsFiaBJttC1ddLGgELYVBhKzZA3i/puSMjfyUNQDVFRH25BntE/YObvAdTWPsRcJdoita
NiNar7ZJ5TZbnUUNNN6PzMrn7OLAUepch1qUmGqualRuJQP8RLHy563VrdY9pF5Wyk/SpqHO1wlA
1JFh5TO9wtE8TXdUQzutp7XtflBKFIQnFqu07wN/cex7QEJQWJmGoni9oAJKgGj23eytAgdK140a
hmlE5VjXms+tXJXg7YU8dBoTU36Ya/DDH8e4ADSr8Qr0+P/n74+wy8Rkj9C0LsrqYeyijCkW+mUP
Odikwx9bKcXdGuco4Y8U+A+iFdE5jMAa7HVq3Y+RvQbnOaOtnM/OX8Ql8sGESySJhv1LlaGbwW+H
jid+Tx4ysc3ZXYYHXEUniepLYrkhJm/K62U/1BiVrOoNqGYbdrBCkxLP52il6Oak1OdEf3Q/XLfo
Iweu/Hw7xpwq1wvJc27pQwGei/AugKoj5WzURUnuzv6Aag3dTOLof7g7PuIrwfXByV6NOjo4IhSF
2r7+RC6VrPUhDbVGBAMhsDmJMlDsqfJ6HuuoeaB21a3xXMFUxizGXgbF6N0vLIZVB82Wy4eQWqhF
vIp6hyZLnZptH/hpELUN879K975myW4Bci/vwXAS6NYK83Ta3paDq9YzjxVV5aM8OgNjYHCicEPB
aumgpYe10aygW8KR5vBanIzus55W7KwsC414Cp/FtqS3/EzdXt+yaYIZiKK7jgpGBxZj5+Gj3mpu
EKIXO4Z1cC1IyUlShzUtdaRK9PiFOWbEkWoNoZ3KREIlDjaLu/WWdpflzjEGubLigfrw+dS8H31B
s1ZFqPBunNPw148lA15vQj92yCMqxIPR9SMnGmLoBMlK5UHC4GfsoguH8bV4MwEEtE3SqldyvcRi
g7e0YHlRbQRg56SsVfo8/wgyOhf8R9eJhqDnz6L25+GlWgMVqOLX6Hbe3EgCCR9YfZR5mI+zXZND
fevZFbvyXxJjXs1P1P4BpIO2WOa3iejjLaUNLHd/30Qlt4aWznkKNa1ogaNtjs9GcaP94qMWvUXp
WYMlDV95KZh8+HDQHKukhHbbBtn0MdZyRgLcy+AI4AhO4vFLMRQVUl+EHVr87in7Wo6ZotWpd13/
YZhxc4i70c3pcxyLAb24S1Y2F8foew9vH+MqwLV4DJq9q353o+0NfdFTa3ZBUu2nFLHQ3X6+p9Ev
9eLLZjbbs7hdp6elMCAeAwvSVr7YsE93iBNYM4+Ay6a08r/5KYvjkMFJvXWE0FfWRckT58qYjHUz
fsE4YN9BiX0R8krtf2W6gpovVJ8XPIsg9bfu0izMw9xtOn0Uuz95GIIcOvT/ecDntR36Ys3b0tz5
/dQbHst/zqgGA5YoFi635+62kHUcZ5+0h7afg2WFZsoOMsp+3Lut0fa7o1OCmfv/ccuZO3H9Tup5
onZqIMKSPx8EVJsSwotFuR/bBRth2Oltx1cR0d+dv7fKSsq4B8MOcP3beKjs7x7Lt5HtTbBz3ruR
71W3Ztf8fKDPSpaV5QbAK7fSLhoicl5cw0wXcZLngB25JyeNRBdEbf6dnJXTTqP89OXGYiQzb6pw
vdvS6pXlrOfiuUOBFp4Z4nzZWTlM2OD2gMrCBOuQ8tBIaprAEsr83P0BPHyOmjrXmeQ+N4K46Mri
lgRokiqf2yzzuBqlFzfumIEGZSxsu8P11ZSFposTMwSS1hThNPWtZW2vPtTuq82K1AYnVMj4qbkK
3UXlilRtty7R90dAs7cNe8skLc9Sj2Xt0kGDIEmKOXzDQG1F40WoQwQna6PoscGHT5PMzNI01bFl
YPwGwFeqL/grEaXZSocSe+9XxubvP9E45KES4UmxhqpHshhPLetyqlhBkwLu5t3fbjrWWdW/5m2E
yd5nAHoFx5kBkHT2OC16q9ybp4W1dTU5wXfqieKanFWmhwCfU4/ZEiPGgUfoKI+6kY3qDNlKNTJO
rVfnu/ZGXFfbYK3rRDktT4Cg/LWsfhvqVdZyw2OMi4Uhc4MU3JvT56HmPstgrgLQdbMYVYyPeVP0
QTZD6Z+NvkN46IiUcVf9YI8a1igkYigoFJa8az5qg2WNYqxycTqmy/k2iY2DPQld/rIFZhGp0DPc
jy7KlW+9yD8lOGSNsa0KcwgPjHVGsIlg+8xlojQTk6dPSsvxP8Y07YM1seqTjmN5MTsLjW2HqJn6
qFvwyGEJUTSf7HqKGZYwk0V35SlDoypOSm3FOkG40yO3tagHJf14kpIOw6KZDh7nZrg/tsVozBkt
WwiHFtvyyMfGjhmUTojT8StOQp7bnnzJs0XqRk2A59jj6ZiuGs5ivASKD/NOLnuxj745w2HZruea
L3pODdZDyCazkLHAsv86dF9SUrAz3S87+UU4bitruAL+PQEuct+vdwLWHoLKRveeqIGqpLWAf8LD
M9iJNpHBxzgF2J35ubdvuegoBrmdqg0ukKtU696XaAvjIwHqvXt13mPkFiw4lyRoJYaB6ouj/U0d
l6WKHbk4gkXp+ZErJ1JeoszJqoiUHKmri6FCQbYiMW6i2JHxlcSa635l4gbNe9WxfFfKo/8B4ZNv
7FV5K3irMX+wiJX4yVA0lTeNA6Y2375jXCym1f/551yvUyXOrLPNiJwfRmBDTmnAbNwPmJ4IWlD4
5wufnFtTyN9/gKuhwcRNVsgy23naDYJ1NRDjXV7EvwxC+/dAADFjMfXLLEJ2YLZKlsVKXD8CRMxX
YoQ1uuWVriMbq3zKcUMz2hDfGvGjv8/5kLgugW+Qk1KVG6g/VETP0RHyb+rT+0KK2aIJNwUubIMD
6D4ZAeVP7nNQ+w8IT77ESS1QKYtJG2qnEkszAKsnn8AMhWCo3Duft2/kdspMu9d4CaNtt2ohCIx2
YiCnVDbL26A3SU0q7wFvMrMx6PhEJcF+ZKsIcoxZmN3qRMkxdZqhcsQoSbKN6DmwNgkja5Hg4o4L
ZM7tfS40hfvJT8MZtRZIwsz6DVkt4fqR5S9XfuEMbmkw0Cj+mFUsBRg4vbGRxJmXgmDHGK+JYBlv
4wEm+RVQO5mYQHi9JW1oWkXNAcT1DaBAd3qelX4i7XYtwSemxJ+tdGAh7qs4UA2v5iQUFdIXa/Om
8cKweg2b98fhI29KWbdABPO3Ky76gNR+A3dnbV71OfEFnByEKU1KrE0/afzTott5CMzN8WetYa6i
1VUrJ38fhJY0WLAnQq7NLY0et+YTRXPZ1Ikxf+O4FumVLWp7Avq7vI/9RtfASdfogKBwYgMk2+Mi
PLEj8udvPEj9Que00OSjeI1vvGKoUcSyvk4IdRxSwQA5Lv6JmO+GHU6oN9AVZys70t2HyzflQeJG
b/B882FPKpbiDn5g9TFdq64IIlDV54e/nEyF5+br/X6umQNBpyudktj/lKFTvV/MM8mI3zgABeFQ
e8Ux1QvLcmeBL5WUFinvPm4GJRhr7705zPSnasaqLXg7JhLbAcCS9dlAYkF4KKfYREFjjs0lLk77
elWFDhmundpwx26akAbt1/aKw185NEYB4zuVp6ETDuU1jkY/I5+krdInnkgfrvQwJ5OBQNa7XQsW
YVJsOghdChNaYKcEikskGCBglfLB7iV9MAhA5uRocfayLB8Tn60df/A05TrI2Kpvi6Y4zjJRcAtG
pzwNWBj5+5/BrJqzpvexIKHkm+qATMAeQC6dNrsh638GxeZ3o4wXMKI8TTWEN8rn8Vw0G5LE2N8o
bZmyRt5Tvsd7uSx3Qi6/Y5rLRJVNZODna+h5hwFMrLuv8VyGLbzKpGOXjdehicnaGYtlZsr1AOIB
OmchhbxL+lx9LeluLQF/i3cqRwOYeT0jowV0WJHHCDSBPxQf1/VXGi73z/Rokct0gaej2rI2wh/Q
hmLYMxYVgXZ2c71WsWYGLDGkR3g45/c4sv6YxXApXqclr5hUjZBT67aiow4lp4SECFiGptePgkBS
aBDxOs2/J21oFPJv2Z8/u1V5O/Wd920cWbI4NkBXHg+6/bWRC1eidHWcP2McQHvb9bdoBQdhDVKX
q56gx14iYjh09CwxMP5OesckNIERhhtaqAKqXY4eo2QKQOYxCuja8XU8a3kHPdYP53WuMB5jI3Z3
sXARplkCR0M+flPjYmGol5shyeIIIMHMl1aJCxUjwWqnq/r43rYD07gDt0pw2AivZpODeB5o6G5G
Ux6Iux8I+fIFSkr3oBLTbqSjg/fb5yaWaVZqhxQJBF1jWEK0aeRTRdkDt9xi7tzKkrLpkpt0f6vH
U2ka/aZqLqxTPlCCp76VqSq24X+lOvmM1T1/ej3ZpHPAcOTbfuAltRwO0VhwC7yE4inQIoFie2La
vKuAqSpArmYh6q4zEXiKCIHom56mLD58pwQQksi5c5lG4giBBuNNCqUUy2bfQVl2frN/H7IMyutP
JUpla0+CsGps23dzM/tGDX64GjJj8kteGwflexYEXlmFykYPjZqoVWdnBKHFA0Yv7L1hDE09wfzQ
Z/zsO0+ctB0kPO9JF8NWT6MvJWAGZM937wqyrPwX/YaIdXPQQ3T7Vy2eVx4Jw5FJjoW481ZL3ldZ
KOylEN++MF4EIms5yh/BlmhE9qnqAgc/FKY44AcKwCQ3w2Nr5bJyiPQ3RvGb51rhKQ87qxPJwccz
xRcNHDjwgKP3jJXx8J69lIJmBBiEY1nkax88YZEssLHCakNBRhDsQBZ8McER7A/YjE8hQFsZEgbj
npo849T8l8gs8xD1KF78T/gglbovquijZWZADE23+dqJb3OTT6FpzyNqSiL3iRgtdiuZQG9dh25N
1Vrdk1ehSrwME2RDESHaIhCcpws8ZVS4OldxoBqylCWtRTWafreBR3AwY449J7UdaW301hkG34oD
2aKHxiXasjEBegMLbvxaGxXzP7t4QrO2tHyN1F4hHIfEylohUCUWLwHV7AejBjkL5ub4aspp5awF
b5SINNcNGq9o0SNNIcS43b3Bfn+HPS1kFsGICU4kUk9wK1rTlcN7vB0dC/lfslhyK+nGhoAf4U8X
OWY5kHbD0+oAisREfWjfhfsZpEUEJbrx1U+ALW/sjEhqJJOV4xfX5EQ6bmD/BOD4U10r3j3simud
1I5QpUCLPl0Vu+Lc2SuQerKrjAnrfPEmrFZ1ePALk+lyiEJq135pGQ20fgqrMIKZTSqXFyDoAX2u
xcSgAM5q2e3oLcCI1epio63d1JRUypMv178GocwaAp+S0SFKaLum6Lfi4oCLHgFLreGALNP5zTPu
yp0JKFCX4Ef0XPJ2gsfrHM2JKZeLjqxOUcvo5776cGG1cJeoAS/gItah0QNkdzZ90wcm4C20uCmH
O8GlPgXl62GrSnmtp4/7RI7tE6oTFeSW4za1RwiSynmPxY6cej40qx0GmmFMFjc79BY0wufTokQL
RqB0Ba8YwWgb99WA9ZsmoeTx12Fvu/7qxomS7U5RGa2utTrqQvlbJRQyP3bAQKb5ZyV+lCOF3yb8
CxBfvy+hTCNdx0wXb+SCDLuUw519m3W+ocbiglZdKjhJQp7IeO/BL+7eD2+lQfD+JnMlNPXlNGDt
oC0aQ0TwfUg3vqDrSv/RyqHHsOLSXoISLVe6HmNRr0M+YzETdO5zF0CgPg5Ks6iw8Io0Xxx0zHuL
fFQ7sjE1QLafcyj76HJ3tc5qBXlnqxph24861aNN91EE0BOcBXBFQPqQ0Y76GCHYxxsFG09obDkO
3bOTrFqXpGv1j/cn3sj89MbFemPcd9Y/fyiBcPn76gqFrBKnrM6YrCb9xDjurplHhjKx32CCPioR
JGPcNmCQHE+ckQjaaART43T5wbPKa7mgYh9AfUhuu21b9KTKZCw8TJtvKKOa6CiE6pith6r3XJRy
i1iyeB2vnyUIdunPtBVWc6jz+B0ThGSqNHMsDRCCISGS11rqtVEF/r6iOG0rPvgGV8tiT0kxka11
k0Ata+S/ZB1zcnfIhUEmoQ8Nbpl7IC9h5BPQpCWPYNWL6OLV/h75H28nVf3MXzC65tklNmAF4b7i
J60CuH+YJMSBVGvfrUBFLU5XG2D6H8lOWTzV0r7R7VtF0x0uOrV3KEUtjT/0Ja1iRWL37iQOEf4C
VGWEQcvNF/fx59TysEfnwIXhwfffPqV3kxepXncPtW9WEcMwyOMf3iU0sgM/uC2ZYZM1byuD5XbS
eGDugIY/lXwt6LNNU+V3spVLM32QrtAcXA2gC/pOmU7Jwkz5GDZ/OINoHpmuziXKu53//sbYFsaP
qm3wJ7aHoWf9ec9EHbZVSts8u3mm0tWcHkQ59m5DrvhqtfLC5zCE51OsJ/l00hyYrfKuo0VDXAHd
CM/T84U6IP4MqNOtRVkEOACSUsV18SrYBA1QLdBSu3VS6mi8HiK3KTR8oR619MPfQxcBmss3YRdO
OX/l6yqgofcBFwucWgmPq7GHyAvxld4Io+sGtOcxH5WoqJLgbte7rMmlsnh7NPMTR+f2zj90abce
le746WfnvZ51XTXihZqcQezYlCJ4KMuxbG8AR73FT45F2G7AWetAxARdAOJFDLE9TQweJkceAgkE
Zkrjr/E17MHg9HY/hR++E40z7zxWJ6t3z8Wj9wYRv43+Dy6FvSdc3EAfx3T117QnrWgtlVN7DB6w
fksMmogDKRxw1i3ZLdjzp4mP1Nrq7740ti3jjwCVEeY6Aij/BDS5tQZD5d+9jUXI02fGwcr0Lysa
KsDaPGNoejQSYNhyDkwqiO2hgQdhcnwusvhuPpE90JpLO+KnDhdHSxzp8mG/EU9IER0K4zvCuUAJ
Ix83vhvqtqNlsbWkcteSLzSkiqN4i7TQ2nf01TXFJD7vVkvMt4rZJDALG/EsJ+VOE+2719cfQk3A
y489kk0sjL+Wo2ohCxtuEXg9LCgx1xdZ31tiOzVxGFNNN+EfPVSe5KCLBJX1E/jIVZVBRezLP2pb
aGhriE3/1cNuojpZ+HxGW2VWWgBiW3ga1a8pg2enujgNMPFo2t1IPa0bm6gipN2LUF1w0kR95kQ1
eTSt/Fj4lcnNt2RA/lYCPrP8gd3WGOJjdgvBEgmY87J5Vzp3TUdphCAMNuf/rRhvKwlO/7HX3URH
gZVHWlKNoagTLoJSyva3WDANjhLHLTOawDvhMM1CPPCAPj4qvjzDQ+1b44GkI1owLBDNfVDhfx/x
QXui4h6/Nbc6fTqc0BSygOh4ZpdGmPoPM69+rVu31ONZaTTcyfPlWroaTkpxPlYdLE47cH9tfJsZ
syxU/t2EN3D+Dq1LYlKc87sgxsGu+4s18hirwyqL7lbbuyd+EwaZG+8n9YZh/AVXLPSZZ6JJMwxw
87DzV2GF2p5xfD0ck4diXKD2spdBImdaJuHMeqRheR8xY/NUvh7rV0QHQFJ2GWzd0F2vSDywf1DJ
vj79QgCGpFiD3ixiRMu7FtjXxD77Qb0cUmR3kEHjt2Hosjk4DxsD/9xYuURPia1OrzGDHtoEIw0P
RrZg1PtDKoaE9F1crRkTN0EuxORu7SpCeqvhZo9OwSJxXbK1Sdv/1QzEst3yTlQc0I9Uo5z9RzXC
l8PO2LXk3PY6Ix/DjGJtpMhoaMOdj07wfwooDdvUujSHewFb5uYZnbshdmv8tyNmEEKqzZPM487A
WOLCYm0Sv1apv20GZahEtDfI8j+ArZF5FzReGg7d/DOcFS9mFSHzKLiaSLq+dDS6iJ0XWbPpqZ/w
dksKGyu8rfsOfljUYuj2JRoNpglhPn3cZj3sRVfD6P7IWWT/N6EqiD4WVP/Mb+t9lnQM+jJ4hSPX
4Fbim6Wf8noOlcQhajo4rpT4OF1r1iW3sGsJWs6a37gLTJKkf4/9N9FzV/VORdt5dj0XtD5QZYJt
W/IQdE2SiWawVmvgTF3Kf/P3Q0o38o3xRbmhOLrAvtSZ3FEZVfFV22JGGFr7ZQnSgKRkcfg9wSpM
o5j8Sx4ymixyO9P//nqmHHhfBi9cq5pWjvGv6L2dEeNJEWtv+PRaQNEq1rn80x+2DNvtsvUZa6n0
BKxHplKYQ00m22oJoQj+LE20SkGTwkl9gixZwnwUJo+8ZP23EkCxS3ix71UA0SMM03y/rPzqa/55
3zfXMgCgRcSTT52WMF63pPQeSZZUknm6lq1yfl+cA6Bk7H7z7HHyIyVSbzaY0VXLCGagAzzSXTU7
M0e3NkNR4EZcnrPHr1ho12BzfFYavusa2Hz20CZiR2fiky/Uq/jb+Rau3hcyBaw5FW4a3YRxlKAb
7k/K9mGG1exNeiddZe03+M+q4a98H4LaqDh9U6yHWOj8ZbNHTHaOtxOGYG35ophBkWHqzKc8OxpH
A+qiZWSseGShks8vFSAx6yD1FUoP3URRZIh6xCMTl0YB5a7iC9hdhhE4eFJx3C1xAV1n7/fEqcBl
R8b1vKAOME/jfd7alrQiR9K4JF7rNEWRtnnlNYIAQzjcZ39Xqg+mt05tRGcZSoOVPsiuzcOEsZSt
PQryPHh0xEx8gT8/y1wMfKwig+VSOOsj3fqzviAZmG0myOWUBsDV+f0RcKs1OV31/HX0YVLsJpnp
pvDGGMqj9vKcRYE20fKPCKZ6GdyC947SfzyfJv3gmwPqjsuT/iOWjlMncF2QeHKCEu+vYUEVy6vH
u3HfCczRvm24pfllGBvG2cCWcqAtEL0rdCEE00SGc+i2FSqMuRkzE5xqz7r32BtOwwvbIceELdvM
YktaiSa46y2sc6R4ndp+zLme+4zykDOnijltZSv1y9Epea4GJLffU9wcCFuYX2epWsXYUAi/xi6S
oSUSlofeLJcrb2loUrkbyrMgdBMaZIteO0iKht+HolJogO4uMElFOV/Dwn9t6J8rDlslOMkwxzBs
kDf0Joc3WViclutGMrc7cUpci4MjSW7RCiOBYj6tA3zMkwowDvz8VVKY80r5gdhQ26dTiy/V31b0
e9i4lAHLLh1paEGeZWzlHNSJX5Vma7Aj7/fM+O48o3P5H91jbpD6D09ABFOKogJ/yhkGoeTnSdtk
S1k8frtz8N7n9aMcKf2XZyruP2JEWCR+D5Co7UuWmEBhSDDwmTmjB07dps4ESjaN9V8QXz7Fhys5
yi4Xy1Gz+J53VhJtAAZ6xbUBtio9NGtg7FQAiDQrWNV0Mmp8dTgC2N3DfgyITODfJdKKXP5HOL5G
vvHxU5KVx+tD8oYg1WRk46B24hnTsXCZmI0hPXXhTj/TGQt3nD6Fag9FqAd5FhtcPxHtFDRwPcxL
Uu71SYlUZNYjkYilYY1HwWkPJb+kVdi1O75NNLXqnjFbSh+noeAr1HCEfP7bxbajLY9FZdCOu77w
fUMuecq1qg/bOoO8oO1qOojD9FcfclyJD3NjF4hVWff64GENK88Td+Z8FuDwHv6ueT8HJdAaq1sh
MWaAGLDtvxfBNTlypaYeBb25s40JK8XEaFQiKtRzz0Y/qOVjB4IZtEj9A2VJzRmURuwJJz0/naL3
tfUy48iF1l2MrUmgvyO0xgnjCFQMV/qlEdcJ45mUeMctu+7/sDBWfELuEKSD/DdtZ65KjDKpJVw7
ADI6iS2NWVXSf+l2bABel6nzA4hSBfZSArlfs4a0bhUFMWIflaV/9xj1rrlmgicvKfp8cR57shFl
kqvnmVeJhZRGsStFKQjzz+JfdnCXFwfCYaNfulaQQ+fP41bIyU22JoPcRNpynfLMbVVkZNR2edAH
iiLb7Yha052+S3TGM1sHdx2ZxhIazfHA4SALL0N5fowGgx5z/QxgPAnvRMk9ARW1VfVcfEXiQSTt
dK+7f52FAf4ssBcwVHoEMlw0kBJFQr7cFDlIDFljuhqxpC8/84DUhc9t/8A1p2SAZZhcsHqE3nsq
pckHqF6Gfs19POC730dXO7sKZe6E9w6xJL6fJiLrHNvUkRpAeMz5CnePuj7UqJjP2QXesCHWhG2V
sqnFWKWOUxYfgtFk2vb8ZwkMggGJIvyYBe8D088ugoonkHn6lw/thBdtstrWhEYYYbTGHNNEwx1n
Q89UDyi2CR3lg/L9WosS2QB2DvfXgcfh/OdGwIL+rOEWuZuokj3+xnr1N9rktCI0wYhg9cxemGkD
qbnuShq74luqnb2Khx7ANaXnKnZAVcp5VHWVPGffYcl/0e44Bq9qvN6IbMAi/Wxq+vizdBrsxpHO
4dKSCMzJNr5NBLBczMspvL1D4zMOGNcVJT1kpR3luYpKk5atVf+SuoIOicwbPXtDy3uTlHo4rDGF
9PyrEYXPXF9BQykC6/PDiZ8Xpz3eAK2bitbQs208ZP8K2GVKrY2FYUiwjzZ9TGV+rP2dccJgsnH6
Mp9NNwJ56um+jS4PaVu8dYwqcOKZyrjoiipcAV3JNsACgI/SUn0uEvMGHm/JcB9Yh1Di29WZXWGd
XQ11ksDOZV6lLzMYr/OMFO8JdA3mMtF4alPLXfHUgWLGzmFHnVLrBrTUf0dxonvKCNSOGciWHuAQ
lh8JPTOdoT1zFrOD4ZIH883hsj+19gR/iQk09YBXywaVv37+wcwzHN0UE/Krbh0HiIH50/s0tyt+
Mi8uFG+pNZUd5uJOT+fKTUDeO62DmzV/D1yPiMFiOU6MJyYiGWtNjI2/1NP9XVz6ft06/rTguEbt
7MiWmzuAbZbwWjTbZBiuYAy8U2HkmB/yrNYaaMLHL2PAUH1abECBslF/1HXI0llzqufgxWYhzMW4
yzauv+IGSUJsd35MHjBxI86efL2Eb7GJIAR+XBzNtYQzX+wLejuUcJhD2SQ6M7Lv1RhHJvZFI3Cp
zoOv7ZzLlM0Y6ih6Ofheeg1eQFSUBTb9j2SLpjOwlWornDjqNILM2XN7LMD+1td00PHv4AezENnD
y3O0Dpat/3pUviiv6uI565KN0dR+mwDDmCW3V4SYc5h2P6X6ByyrkzdS7LguxRvew8HVrQ4cYpxT
V86lcZy6osOtSCzQLmfx0s7W5DxDkPjqKzEceOFkEhvtyGFxaL2CcJ28Iosz5YBNMF2xKAOXadkb
QqOfLNLm9xaOszjcuZK0J6uiWBhNleT1OixSAKGVya9jSRUwSNOjhnftlEWisR/vIfeCz6lri2IF
gBOJ/uYUGL7XuRYZ+sjJePQpWTivI1Nqe9PNotcPpNK/zEJa5WBrkNNyj8BZ2VqFm+hfbdxGiNOU
yuk4zOPouu+K5r7KAZrvwdOYAXq4RJpRH9fpX1HECQjZFjEg5JwrIVxJFcCqqynmpgqgMjJAvstc
hFbDe8/NcxsLx70WjVVyYTLHM6Gg98an5EgmDdVs497CEjD/1yn38NPtNC0fuds761h/LxoDwojF
VwXRpm1EwAaltaQ2bNCuMgLfRkwTjMMr3th8eG08ZCrLCXvg0FLxOHhlfJWd5b0TPKjf0ikAhPd/
U7VlcRmRnd2t7L9PBYQG/GfY/c+Tf67wqdGnFRw6SUoMSqpUynhUr+9cMdUBPruwDhMFFlFRi7jR
XCen3EA7jbrsu3XDsRhtb598Zh3Ji0n7BAs8xH2/yLWUYyi4c3AUUDsVddV6sHwyji1ARJplTawz
6ddX8wILY/dnCBCaRCsjV3sv+qsc/Yz5h2mgOInxKYhLMheo6viSFFEpU8qLU+v24OtZ+FofUDTn
d3zj0vDZSTZidHXjrHktJRorU0ju0pId3bpN+XZPrF/voVLhUVkRAGfgizgXopUNl8AKjcg+9qe3
4ZlNJqt7xav/YO1/82x+sVHAuPlU7108en8u7tKM6RaJomJufcKmVO8B+bCQRVwtVMsT+hx8l1DI
9jLu6n+bUU1Z9qcisn+C3nM7WpyAl0Y0rZUbgwMCmWa4s3PwxmXaxbcErf/B5qA/IsD4b2GFfHtq
BSEDkgtHMWvakQ4GWRJtEM0Ff+Kz0Res4/mEYyQfiG456GEBwu3z2bEqbu6Ew+L89sjeWq7U8rWH
IirkCgzgmFQZpuK8U2g+yT24ZPD1sZUZjx/jUEX1jdg3+0Uh7DpVm/IinVHmwvckdxEHdueXR/PE
YnlmkOznRjLjRPHPeesPm3BS4ntGWA7PyZMgo1rPOPJp6qQnMAqaEgCdaQ50KA0NIxtI/z/7YCEU
pKnyYxxvB7JgBHSBLN6+AsRywu7kupx56Lr9Hyskq0cswJpJekHSpW7Cb0/7EtYJaBl4KegAMz86
MfKa45YJ9TesUdhn49qX+GFh+VW5hpRjjuofn4Fh4Ee1cqIw4KCxngHEWJu6UUvqKKDFnSgR8ZgS
J14qbapZ+IR/hNeP+Kp/nQTihoUzgYNK3WRCsL5HRDo4qGSEcjD/VlVkBlO8s70tTiZbVoo8vfzk
EvRHTghWrFXdLN61ttTtM0DtnOzcd4a/3+vKRt4dX0Q86xSpBKES16uvHoAr/CEwGPUc+cfnb4Ue
aXOygbpbLVeGiqxd/+J9mrlt6mK2ruDeyZcGnhvb455g5CuG3e3QjgLCw2i/PkDqPevhVF9AMr+m
WhelQ6IWflN4GBJ3s7vaZuytEg6L1NtSyfEMpbiNnTStyQrgCRRrsMjV2IsEeiiogQ40JJ3WMPUs
GisoxS9OBqm/xvmcN8Ra7EGI3IwqysfVQ3Uojma3FYDVsWElXawKv0ZO9dTAUHXLzVpZjdFRcHs1
yzmfwqebxXoLWL5VTedYTl1PZmeuvNr/b6eRNhudp/WeBpxp58jlAJRJ2JzIhvGNAPSZxr3M8mOP
rGC/WZ30G05VoYS2YzZ+cKBECC4IxOdvhj1ptLLjMN02TMDwdQmR+rgYExVwjGf3eQEGOzkmlZZL
t+Dk53gkSODDKErEs0XuTMLVGcPYbr2+QyqnQoApP6ni6XO6NMNLM7EPylHEDdhfNFzRixMVEwnq
a2k49RRisEMVZ/kzlxItSVVFbUZzA5NdqRxBPzk09JmI+FOr9IGXvP1xjiqG8h8qicnP4VMzBTUS
ycCosrOIpcpx0+BUQjhQjJarNTj6c26VkSNga+o4KflJ/jC80hvgkIrPuoh69UurjUOI8vygMZ1H
IWzoWj93GczD7pt1+xubU33pn30X6mjCWVBZo4wz0+PqkokJPgutNnHoeoKzjd57Q/L8dU63wXbU
wa/SQjj43RrYBHBnL5hN9JQ5lYJVDhrAcLIHoBHhPw/dv9Jlc0CkrGnXXTM7fBHEfj/iN5B34qRr
asBSCstVyaMHb+GnPmVvciVjY/7czbDZJXyKSGVz3RJsZ61qBQ0hZsd8iEnlSNwPhJj6RP0YdWXd
6tFz3zYplVY297EClGy0+1sHDEtuj8PuSdvmXJYQUjskG6RApKZsjak7w0jSoUtGNJcRwU2tYUgD
86MNnLP2/+BnpbqLJrCkrJimT5UMzEOW1UIYXDAsOkMZ0FNUANa67MQyNUcp/QOvD8wdDXeICL1Q
pUxEV3NJlGLn5aPhyoqBXjs70Z2uLhOTVSRDu9MT6dBLuE1hxd57YRW7UoHhHJb06SiCJuSFrkIy
D+FPo7nyQU0+bRtI4SAU2NBBew6GRaOulNsGk2KvNdcqXX1f5bGYYX2fIp1Nb3Qu3Mk0CjrcRWwH
4qdpYnhNrEp14BHhShDXL+EWNy1ZOoUmELsBhKK0wbWuJZi+BiacIEElogMIzxL4sIlsVFDMUHau
lsj2PkzICKvVnCa2d1iSLmvj/zNtaOaq9FdqOLRbR0ZpVr08fbClz1Ex6o1r0PxFlmHh28OpjJi4
1GERim4kKUgpz+X79KK8olQy4CJuRwelMMBMRKGv/IpoDltD8WaDnGfxHQX5/w5ZRhKAFDgfXW6J
SJBC5SQze0/ROnNpxohPdfec4oKj1sjUPRlkSCVDCfnzdj/rJw7lwPzGAG2cwWTiXwIqQCQY4EdL
ts1fldqzd3jfwLYRZQzC/E0DA0D8dki/+BatRdxxwdwhJ1ouEzcoI7JJ4MWiToEMw5km65MU7IJf
xETfLxTTlrPfIA8H2fYAfOSP/V+Lf6+R8qmcEE1ysr1qL8XhfmDUOgf3C2Rcu54OlIa8P66xMomv
rE4GZ67glKNYXQVc47Nzoj7I9Gzj/lsnG7r7c7XEfvRq0EuC/ZpKhlUKZfUJg7r9KZJiREPk7Bjn
EclIK97VC5VTZ1e6+QDFjcEmx05cd3Qjka3HaQ8PvopAqsZ9B/3p3FNJK5aKhuWZSl5IBrpMkbn4
1+h0bNgHnTWzmw0BBg57yySs0JENoJjAn1z4gd6WwXOEmV71yjwkxT1ywdh0x7PclV11JsNTX+MP
+jw7CA7N66kpvxXWikaiC8ymmwGaRNM9ns8eBZpFBQ3qxtnNWrm3x+v3NG/BqPaPoeYtcqS6eR3w
IKmCdkFHxCWjpvI2WoA6zPIOxHrsd/vVX9wUKFIMG1DA0FwkMu35FtSY9xbjSjfF3Rv498booZhU
DE3hWh+iLvS33to5R+ghDHBHiwdqWAWuXya/UpYykBAMcQP9VKnPfNVdQaKNfw5PpHSnHgvTZ73Y
FZA5j+kWAi00EELJY3QRRFE7pB0WdMpv2fDwADEbKFU1u60LEr57Pm4vMfXr0fM5vHzRAs/g1L/T
sz2sfarQR5d/mvx8pPCONQ13eaDKWINXAMcqM82DFXCBoCyArg73P7Q/09uvIVzXiQZH7H10Law7
U8eKBCNVz9wISrC0JM4ZZOCeCFX2zsJagrx2hcVfj+oJaB5wTpDes3arS/A5h5xQiSR0Qx6vuhLe
NS/9bAT+E7by6fLs615FFVHHzlwnxFIJ51mmVRg6EChaPjV1IiqmnWWi5Fmsr0DwCMze9PpglqtE
hcIAyDvUo8rdP+UqiEtOCtkE7OC3l1LRp5lXJc/ClHqr4YhkKM6yy39fpWRyziL3y7ix+9nSyQNA
KAgmJLCXudCPgCQP/JbdJ0nrrQh10CjJ9YSsl3y1IASAYw7ViehheqzxToN+Zk+jYMJxCOklsGOO
l2lDy14UlJzZOBsDrk4kHGhEP241plRpjDpaOtFu53YOfJvqVRB4tPxhRrhXqZJq9l1Ol77ltZxZ
plKsSgsJtuixa3UPPkn6jCFOkX8L7NJckKtmQdWu0FeArcoFbZOPtxMxTYr5iiTCEkVMFGUSh3Ll
37F/5VXaajJD5mo76UfzKXDEmxbHoanKdT/+1ShRZs5eQZoyDkpJURGC/SMZah8JGCGkSAgZipME
L9tUx0TR5F/8rkRRLnmsPLqmbWQF+tp8i35Mp6gQhd98QMzaCcRaUD6aV0OhaD66sulPiPtYMr9q
RnowX8TgyY2FucfYU9EfxjBC5hVEMVsrQdlISDm4CPeC726D/Ic+m3dVM+vFsLvP7mOux99b7op/
TdGr+i7zX7v8RoYt7u6rHlBZzudMHcgstSoZ8P7DdIjyY2MDQ9FCk7yxD3z1gI5jGrmyqrzYV+l+
3clxx4wmFKHZkECTmwDO3c82oqi/WYQ0LsqR9vkTVN2gO+JUjMeFindv2VQsODJ2mY9HUgDyVJuO
NANdevfHTrmJmy52lXDBgBBeGDBvxKjeFEc7IlPP3X3DmNV5j9P9z4G2AxSuvjQoAAf5/ff4yBA7
3crj2ANmsZQHNp7DYUUNfqmTWKba9d0AXKq5lwK+2Tk3lgR7TVcLf6pY//ZFNrpurhVMmG5C86vO
JO3Is9m5FfPM2+ob82O8vEhuM3WVQ5SfiULZx1uEZRpalRhqhk6ozqSELqDyifMa4TleEjIrgRmw
NDywKske7xlfP/JRAz7E2zC+YuSEq2nhWFuerHm8u8F+anIedIKfclUFu41NaXc3LMzZ2WOy7XzJ
BnjlNmDa3M+CDRRTaKOUzxR4URr+7sXW+Cg4mGmCSZLzheZ89jDoO+ofG5jaXxb6yFBdDUxXfBhB
t8RMsBZ/l6L0A90xfGbVMSSufnNvaXxIMAgWT5TVloxVqvWd9LrpC7oMNmIkSy5LqcaTmJj5wbLQ
hoJlV2XOoFph1vg+sNAnm+YVaIm9e0J8ZuduwkmI/mJI22cSBMlUIOVOQ4EWWlcdNoYagYOW35yJ
md6DIwrsw6UFmWfgPHv42AUVQH/aoBRkhUhdp/IuOiJUkwUCUCHatCMenbOmw9O5gRCiwBVBn9DU
HQw+qTCZZjBhY/IQIXOiBi/cj/1kSRyfjHQjHO2G9ypq0kHBIQYYaDK24FMCPFWPE1AlaG5gb+R6
EhVMPH3wHRNlLW5JyHo9TCCK6keso7jIz662ADOKqC0sNVvJF5LWX9uMAAJl/oC+qmgbLlUL2LkT
RfmOg/aIJNAe+xlf1OcqLQu7FMTL79SXsYv7riHfkTGTDLCjgWu8KOCal3HP7qPHN0gkmO3ZGuV3
dp+yzeW131+MSy3isjSmZ3vWAbwtpViqX5wPmOwS1Shtt1qALa3PWykIKBFdzEAGsM3MqNv9E4kB
OsLm+wOTNwnsXxH1xV+169fwLDU20V/i40IWZDZpjPrrvX3erodz+I+BoYZihQN7W2y3zBzVDRUd
UntHsEQBCFtir6yUDeX67jG+3QwVrwVC8SkB5vMsYFjLUw8lWrQeAooQfzKW4AbOqwSXgu2AxLaw
rWHXD3n/JlXpT9vcsuUkTslRa6pJrf/Rb3V94CcRdM5i2vgVlnWgr1QkE6vjNa1Ftp17RUlzFT+j
XnASd/oY/zUDyEkQOn6P1Ky/asM7qYN9y7QalIpUyJYUTLPcmRJNASDyWe8HiBn0s2KgHym8ESzO
XwS1yFHFcQ0b5Mo0Yw2D9Zzl/iGSTSxx2j9S1/I6E5ujnMSkdhi/F01cGXINilXAvnICeGcpLbrh
eUmEO+NRyDEumdLE4OsZHZOchke2orJWgTfW0UZSZ9tIwPv6NN7sp0FmAytK6DrRcAP0cdAZErK8
Pd7SKGDAhUYLD6+eWM8xRDehyP0yjB4SzZckkjMygm4VeRYAFHiwF+bfI5+uucp8ruPo49Qxiw9E
T/M9o5SfSJ/bVuGih7nxUcEvZQ6xxO1lYRADVT80ALtg0nFgl+X2hZvqe/Ent6AReKRhLS05jetq
u51uyOqj74DQEsOA06CXk7SGtRYJalcfHjJS3MjJUHzcNXLSm9doHkPD1AlRoJ39z3wJXtEFt1/P
a+aTClw15HXfVW2gqMUoT5bz0TZKIWP+2e+neUk8W6UQmQIu7iLvs4yt3OkdWagbb8+P5QrY0sd7
ktuTEgcqtujUQ3Nc/tTd2Xr/uU1cexvk8RaNgbLegohxXvwWrxu6JOKGQHWwJU3NPj3ECNPpf5cD
Z5Q9IRoNzpiAoGFxJIBOFsK7j11L2bD3FLlu8xo3WXVcucfKpD0oQU1gxFCuOELetG5toOTx0m5I
hBBBXiH4p9CbF59x71H6rHYCRbe2hTr/pS/87wOQ+IWruLwzGUtVAC0NVt2Sl86OnkWOJVCPdTO6
4skbLx7V0Ua6TDGUAlYjDTTXBxyRO+lrJj8pzm7TrqRPbpwyvG+xRGHsIGS1k7QjGdK3QFB9OvvB
2b7M+9XeprPEWq9gPAsa588wdSMGIubqFAEjq1adIHM82k3ccqgKGzwkVLpOHv195iqUeuMDq13h
bD3GK5brBpNBX42bopa0JLMPK13DqbaQ+1qEPpQupgWqErQ+p0ga0CS8TKWrFDgVSPc/qv+vzRBK
/wgTX9G7ion3xCXE1xgLBidsfaWrqDzOjR6wH0KteuRxL+3Jgku5eOnYyqnw8A447Pgc7jdQ6kIG
4cPYH8qXkKT6aJVldngCgc0it7qt9U5Ij+Bb6ggdaARDNQCgbJZOy0fefoq+oXIHXiuMWpuIKRHs
WTS8DUGYbOzSDma/hj3jSy24Mc8//WJTHiATmfbtSzOV/qgIj5txTlsgyh8sKNW2fyQ71nyLrC88
uIzQPglPv8fdv7ZLgJ+RuLDA2/RnMygCyKodcKY6QlSRnZPYRYkxLSEaSr7L3AzT+HrhHS96HS0u
W7QUdC3IVjuggvk0n2GsfFnh9w7ezJbSrsk9xSNM/HCEZd2Px7K7s5h2yY7LKotYud5txfE8wuzK
8x7Z9m5vg7dqFUnwS9SXdI38idt/zNrrrdR4kOhDbdUgYsAA5vGzSDghMeKVBapIwlIuWAsH6ny7
9shKoJPz7cfxNUN2l1UpWjddRXLr6akc7kmghyFf67WODDcBWwc9zojFq82MTQeagozaXdl7SwUI
8G8zp7U6xyqavGF0Yosfkmyo8YhBKdJ8XJvisrKgq5sQXgvE+vuOAlVXcC7DeplHCUxRoqchhN4u
vYzxLsdZU8LbwIlWmogF+y6l8GXS7wK2ozu/fSS1M5dPdoyZElg2hStUQIyMV24w7IwV1ziscpRZ
knhrv/P0wrROUlOVddwBMiMKpGWfLsh5s+yD0JiIQ2cKqcppuaFe3jP1ZF68nRCOK/vsLVb0eyyx
0jNpeYKgMFlwFW9Stg7DwlzVzL5/lDZxMRkaisEGix/4zmxU9QXmTVLqDtpFVCR5VrqNOqVtwsxZ
hZTk4SHksBROJkNORwuQI5Vsb+L8Rpv89H4ceZnov/8dqpEJRreFyM46hxJlnpQ4PB2/mgqgk0PA
XVT5zUEoSnko35Pri52Q+nQAudiFaVG5S1dGPPKbo921KLie1glr2DTywY3Dk9f9yvhzKZRdNx2p
WUZXpPONViJmCcnwivKMDqDgvfOGpcjlg7GVYuiUPinZhjeLtupvsyLhyFRRrFzxxXkQsMmJ/d+3
2GR0prlqDdOStQYtfLEYo1XNqOWFqsCGnjK0AbLW0alCbpwf1GJu3kpo/btSz3FdkVvOt1o+kGji
gizEeZsfMp782Pm5qd3MzeqSjY+W1OqV0FKMJRVkmtI1Vo3qoVmwfZHfnRoRK7stiiWh7lbVc43L
FlTon2iaw51xMmB/oPLauuKd67DlUMjU9r8KJNvM0zGPQO2geEyO8ngEu62KzAINBeix9YUc3fS8
RRQ1FZFsDHbs6c69y1RxSKCnIkZ36L4VJXI32bkShJws/nkpKPfNOKPUlPRND+p8IQ5GnGjrfPdm
bjaLDBXVyz3u67p5t/EpPPkeamZUTjM5UOSprpA7YsGamIeH4VdQZf2kGrRd9S6qXg88RE1BRe4S
5JT6Iwdl2mr8C1Ps239+6aHLgb31QJq4vvAn8H7YMiih1q53XFNJFDnJNdO8v+/bYwUPFJrlrP9W
HvNg5HfZxg17BCB9Ki1TkFM3wIslR5zzZbdxK+oZBxc6yZIE3x0aq5tl8FLKY7dn5VJ4j1bhRTxs
o+O2HOqagX6dCdo+yRmidZURPDM9T2zrjChZOa16k1ZLcij9Amqb7pyfMryt+nq2I7sPfVRgmAti
TBFaRxhur3FeJ8cW2c6VKBIrCk9Hpq4ifmHu7gpignp7heXsehJbvvDwujDYER5wJp2UJO/AIqzr
XRHsMdhE4u44Qqv5GqkofYa3gW5H1hfr+84tlfoiaGP3biNXLSzxSTyoLmy4NdRMBj9ZqyKejT5s
V23Hgebk3UZw06I2fYQPjqg6mES3sesmBeC3rqiO0JOs+/erwcuKK0VTCvmM1ywsU8HurZukddTf
4qPDGkCWDGKRwwu3OemI0Kg8iMDUaEj6wE84f6Fl0r5j56YEw5OdWlswxzauPBootQZDrnHWKiwc
Hpv9ywqE96xSxoSpMzfUJaviq4M7tKDo66/RlK+ywsLImKIohyMh+gi5/SxcxHgFx4bHx6H/jzsS
8Lh98XMAe7nZawBNMwtCgp+bdfdV4qZYWDCNp+LM7HSI+gL2HcwIeI4EGySnHk195HXG1CTquAmh
5LWc8x7Yf+TvG85JfYbSgshh7S6y+Bnu3dOaIrEWimS2k5MZWXyvFlmlKaNmXKtM8q9yIb0DNJua
GbFyup/GcVzls8k69eYfxbkxtl9hX+39qxwUGu7aDpm0TQMYkeAAMblYu9h9qfgTvvpqOkOA52nw
4vRFSGARKGvxhs5ViNKAAXlCFffp0WlPh9OEpfCORaYSCZPKEfUZRGaPPUZIF1N1a+mvj+/XW52g
FToCbSHBofeOmtgmkKrzcrFBQorYFqvHNHzGkr9TO7wLSrMy3zEglostwxbwDTsm2Z40skpimRxb
MtQBweZETG/woxSG6DAKn0KbEAoSiXs/HdQNmnGdextZz/J8nIWnRKFlBWux2wGOGI15HQ4t1BhX
k7nJKcSvcX6ByN4RSfwWufzuEwamCaQieC6HiIqs7ltjViYc8QVgjNuLm/5yRp2sMb6VzPPx56dt
Gp2LGEeljdJQRROOqhu6MIBTc1BKcP9NlmUzsff8oWT+BqduUmSfaUPL0d79tHH7gsDdJs55EXbS
Q9qoWM9i+30R3Z3J5k6fGXQ5/+PadOOqq8FB0PqapUAUA8A317GPKLu/ZVB4S5zuLrKhfX1uz/AG
2LWzMxyzDEpwSntVNDSF05so8NHX6QNclQc0XgejNBhisR4taXoDVJKtH9p+GSORKfcI+D28EHfW
wKD7VlvPajSnRJ+BFgzvhLSqTQrua6S/T4PXZsw7hyAmlOBtIbyvrKlYljrNcXr1u0G9YZdCx5Vr
7rYI4M/8mkxAG15nTF7m/lrFZojjf4KKN+v2nojZkBXZKqQ3Vq6rmujvW7J45UUwD8nYeUE7JTbS
s50bkZ3HELBPP4ElXydrFabzFNTM999B4EoGMEuq98oGEw0DRXcgcouYK+0Tx/yXmF4Ud3/8YFOR
NaKwEEqS5WDJcX6dsz0GYR3j9s2zRHzb280DFAnszAW8rhsRvSJ2OXeQygTRYfhDDFRopQ/YdK6Z
YZJE9SSjO0HAEpxjgk9fSt1mtlVw7PCOhMP8Y5V26YGZAU9UG5/z0o9gJGSEkRxqN0T/f8MMsrlH
gUZQf0SniyWD0tUlkUGnlikcKdBNvbpKxRl3W/ZhCW2NfuNMsaTA70s5bG4lN57Kt5V41osoT9ij
jcIhUyP3ermKU/5Ive3iDhyw0d3uK4CB13ica/tV5HzHjJCQfjPk0qtBSF+Ti4PIbvKB+WDC1zZt
CClCPzREuHulFiVxNnjfZe/nX1ts4BOHwnLoKgNNu7CitK7UxYJUXvLs/UFbZp5YhfQNu0huNuQL
qcDVsX4BboFd5awFglPleX/VH7y3V10jzG69jc+/vs5A/YpuJy2nqDk4VPclpiLdbNcnIbzZh8Q3
Vnf/LpNjjauLmfE8zlHXmineFhm4A50srXWkiSerJeI3Lo1wfRkl9HSC6diTyuIibeZzgdB4d9h1
/5ECWNWMviFwzypbTgTNkhrELjkNj/RMjTk/DCc3L8Mm65yhChF1KpwKGCj2v8pb1b2r695F5kUa
81MnKJzK91Qm3QQ1mBZIDTu9JtMhn+lEvIydvSvCPRObJVFebml4wF8EeD0iP4sRzlj/5hEgjo0j
DpJn5NeqtFgbmvK2zSh9C0Lkdo3YEJ5xmHMi1b7MJTPZ8NDWSiHuDCes7f3vD6S012GshhZXMDSM
9JQ2T6IlJ89kFfFgFLqoP5a+WT4hv2meRB7byJR4T46nahDZp6q1hUXzxN9OSqXQdwEtgBkRO2HO
hA+brwtO2TjsYfgOmjPR1jZI65SzrBVt1HtXCH0iCCutqPhDnnRyKFvNttSdI0UsWezOOY35nJX1
7+8+Z1vSSXRVwVDYdbo6t+9TIGLP+A5jc/i0RQADbZOiRVq0zqjbYJzjXbfMfdDEpg43Ecsajz1a
hMv13ImXHG263GeMDZJjZiyKF0Cy4TAJ9ufg3C7swS3Bys7HEb/siDAC0wZ8z9clUzUV5uUdIsfO
zxjavDzN6H2qB41kWE39utkqlSGVlr3nFf7t5lXYExlT89M0ISsmVDbqb5bNFHlhZlH2Fg4YoZmW
ozQrMqerdV8d91uBoVI1njNUd0nsQ7jgcBbFPDVnyknqklrylC2oY8fDUQV5fbJcGrKdRbAMe+2/
+GhZtRva2ST5Nd3mY/500H6EGO+sGvyQ+hK8zgikUU/DeoY5iPKI2Q5Hyh7ZNcK4uzluEvPfY96X
PIjsSnUZNaFj2Ts/JKji5xIZS6qzQh22k8ENVAAMfPHTaak7/R/CelXWDRbC2oORTu2g38pzm9Ze
p1arVt7pd7jnNEv5UMaigflRLzXxWl6eqUk3bCjrjTCDQMWCKM6545HugYjDzKq+mjVxlUUOtD4P
rXS6Ivz3m+rQDbllqxDzJgrqJ6rbMIhHjDAIWMrQmzrPs9jbgXG0c3wgDaTSuxFxLwJi32rR6K9x
SmZdrByucKDRxTjzTGzuW0NCMcP66hdj20fF94aGCktUGMEqYcaPi0+ufiPa0uRoY6U7OhuhNw0p
hgDNw6IvR2AIL3jyd92wqiYdgzo5IwDufBol+H6BrKxBAWBwtQJCNKM2rf5qmht37W/O/xJZAYhj
qWsGvca7tCbSG1v+dIEZWS009hh0qnN+vfdCqNlXVzQty/4aPSjHCIJ3m0pxfj3r0ByDucvoOQLt
2tWoA5h6JMsMl6lhQaLPiu77p7PN1NsNPM8zz0M2+/hm1GJ2qahKiFAiuwW/1YRGwPW8qKVLI4P3
THt4zWbzmykrZs1qhQOQL7zMb9NvWXitl8MLlvwAYv041iz815ZVWTFrku1kaTLO8wZdYJdX4qI2
F9qeckwoIEBZWvcoFv0Z671/LcsCMN/vaW2grBg8QS8rVHzA1Jf4+wqdl2MqFxarJHrUa3u31Ph0
GahwbBfljytdvWuyqUsUAL9hwsDrIuOKPCGOkDhdhwgsNHUHQRqUAzEu/ztsw0G7c1Lhuj+ql89f
60uCwYUJ9fv6z5CYZLpTtcLwwXLahlFtTa+nytAzTaMMZ5BoRi/iIzCk4SNJusYcy/oFr57djJZp
0SY5god2KMi6VL17vCTQdJMkGmeOOMov06sO32TQHMaofdZ8SLYDTNrUFltLm7XmB7GAPmkTueed
b+qPDtTU+DbzfjWzrqOE9FuonNs4aoIOGDGJCF2FF88U33bHqymZC9GdNlcvck26sR3oDdOmTiyE
vIuONLMROkYxjQKQ+/pgwSY8OPgskAUrKWg1CgWKkuogT/4PwGcTtd8ovoKaBEadtjaIgbDbefX2
+FJ0PrQCR03QBplsM1eguJUSOUO3EFn6L3OYhqOvraPWjEDpDwrq3Qr50xDJFg/c69+/zDlAK/BF
wFZAK8dynP1lfpCR+U0/SlW6TdX76cx9e+jzSrx1XrO5FQm8PJHpesUtGG6WXTtRkBiRCQbA2TZ9
mmmRvzUCSO3pdgg6TGPKbL8x8kq3FmwGMWnjnW4eV5miw9+6sZR3LgWOFg2DaEMvU5jSNHFfUexY
GIK4lqcinZg606hqtmWfzF/SucVO+5GyOgH2x2s0qEN5nZD1qHFlTCm6R52BzKXeDRLc0ADLqFdE
CekIf2AJXuvvompHmx3oEvCmMLBzOuJlSAmuaeYdYoBr7HJnUr9L8ZzstgTV0N/9/5AivP3q3uOm
nCFGsmutwtL2zLR1gupsB0nBcLR2X5zHfUz3hu4BqfRfq9tFgjmEmbs4VTlQPOq1sTlZdYgBfgNv
7AenwaMYJtxTu+EH4C17DbW1EKAQjCKDd0MZll8lTvlrPwYLKDQkW5YIRn0R8aNOx72FywlP83U0
HWDF8kl/IEKkgZZHmdWK4ZGW0gCtLlHKQnC4zpCF0Tt8bsPI9anER4mu55B95zOFZewwIZk/Fcci
bw87BEfsmvvJb7GIxIP7+32YxUQ2AJZS5ZyPk+RYeXBVnp+KWJyhNKWca+gtIgdFwdX/d/uzRtJi
alItMEJ3w9QeFrTLMNIYTc3vh3u5bE8jhBqhP5wI0cHApNVwk7aLRAIG7E1xRwEgC9pmoNsdDX0v
k++uRIg8tB601YqLQ191m3LUQNYYu+lzT/WTWqYpSNZEjvHggobT3DSoieNU+SOHHrDqyZ9jxYGC
/aB4wR0gBdH/70sk/0/6PBrQIHGgFe3QKR52OIM8yWyLq/pYS8DRqCWCGgSYNLsdLqOZW9hnmIXe
+llcx8oiK6M1pJaBGNUCxsMO59CeRhmJUznfxCOyzbHNyUAyTjC9Ni+ZNUrsD6mtP0gijr0PjBI3
lv2WtLbdmT13vHJ5LxxIWIuZk7YoXW9L+NYfmSklaYdrzIDArHUuCLsGThq2p+SrXfxLpj3iAR35
g7YZCwvLBgaDWWJApBgyVzHwTSfinLkTEXphm3uf6wUB66HTzlbBkgkQ29MKTB4wBHZUC5xXyhLs
8ZywuOAPpDF0/0glHKfP/8lSzBf2bCKCr7k9WALz4ycH2u4fBIYsWWiXjb+X07k5yFgUw3SNwBzQ
g4sZsFbsuiOubM8oshSAbapLuAvA19yBDqwneVCnfVB7s3WktXhYJies4lLuALolQ+J8lryfXDz1
38YjSasL7yK4i3lwIooHT4epLibJDEXCLp6XN/BLK7W5R2jR8+7VUi4K3SNTuuPeJuHRNGQ04kzq
PMYOsc/PN/xpkzLHNr2oGgk78KB9P20PAPUL1U8usXZ7lKssS4AyG4PejESr5vsXpEAQWDRRT2qU
h0zfTLu5la+Idu1dy+Y2DBVRvAmKyHKx1cfkClotGXRRv5w2q8YP47gHTQH5ClAzMdZ4QyozaGl6
boRtPeKnkMR1fPiAjRtXnb5FQOwuDJ0FdOdDV6PqGZ+p/j3duZ5WTKKlGDlJ0+AuenfMo1x2r9Y2
sywGwKYUl2CbV9W7S0Xmydrg1EgNu5h/T5beuIA+UixByK11nhqo8Bzn81WQzwQDNBbaGkjPMmpp
S38M4S9XuQV1vrkLzstAZJaXSOaBWULDIZKxt3kRyqDq06Jrtm+jWfN7rMfe1iTxEc8kppr48MUW
UZD3lC9YI8mkhSCcdiNthdWclsj2aDJfDhYW8ncU3ClGY0gkFDgR91Zsxtiw2ANkQ9zBhkeAHiE1
drfgb5yjZIBhVF9m6p+6R0t/l6LFbOAO6aOAqAjjh2kpfMz2BCkl90s4bzysRp0GeQKiLwoBjDIi
/UBqx3B1Vbqyy+k5DHoTWv2A80qPg+aTu67U88Ka0brhfIX3UOwHv/HF4B0hB8KUB+oMNzYrc698
liejdnF5tRhEoU5JsvnDf+iRN6dsc1cDxJ5fmijr0um1yFlg2sv9E9nAA4AIKts80Ud45gFwbVsW
kKBEWH1DKdYvUNb2c+ekukPJw1Z5SmcndOZJQGQlbIwzo+vlXtVwec/fbng/2seU6xmZ9Wxa2Vn3
9lotZ/DA1JICa9ywFLeK1FlRdQ/Qtu4hIhQq/weR+vYVvKo1PgGHF9sn2FTYmXYNMN43NnvaYZh/
Yg+yUnVkINVzTdKuuoBeclV5YwC083B5m3nHkO94TFlff5nw9jscGuyb0yYg2+SUJvwFN78fGyXz
ewGQew7KbN41i82+wdVb7xMs9MOKqiLXCelIxqlXi0/1KankTJ/WJDqj3088382Bdlsd3UpQor0/
s98zlHr6BEr5EImRSYR2EWJ7i2nZTefkoQ1/TMhBRY1K4spJy9CLgEOSJoe9kU3FiNJScCvxTnOe
kf42Ft/yPLhtuzpmjErvc4/cDxlZHEfpqh93yH+8MPRa6LQQTBpZM5ZCo7ouFyHJ8Bq9OLcEPoYH
FOZfrDGL+L8wYAPGS3BbBLYWYldsKZzCPWZTFELZSG0Zr20/xajgi7TpKOwp8XCE/TV7L6IR+FCG
Uv2Gsl2AomzanyTFaMngb28H7gzDLBwLosq9drW9OHnTLvev98/HJRdCvupvOffPVqFtfRB7Elpp
2XpZoo5aPI0I1FLljBIIQLJ5oEmp8sOTqrV0LYwGlW6tqLGcgbM7cUm7z0wsaRN6zf3ga3dYxPZm
ppMwgr5vFT+cBnd/ZKlO5YNudL1Ls1yQZOkE3DIVhXkvOd4KZsQvlcftP7h/+z+te1uQn5TGosLm
7gkUXCVKTp3Mth7AsKVfKjrppY7GGeSHAQwZ0apXe9yIDkNMwfVNLJljgZf3/fv54XlmDbL3DiaJ
FCoY3iIeaX9yq7kleMqrIj2bglW9wSc8mGLKrz9m3HZRhHyKw/nBMoMcxcrUAeziXWy1MhoWWOMJ
WgxljEe2l6SSo02QrakdQtuGDlQqd8Lw61xfaCYV+/tjh9wdZYyejTsXdl2NtKnZPLywcCNCj7PP
DMpsHSSdEW+yyy2/TSZY/SBlMUTTSzKEajG+EReQN+ZRDuq1LPDKFE3SM/jCbi+tLJFtMEUVHn4+
Cw0bbXkkozSvf8agc1v6ltURZSSy9SqtjJwmiQyKmiCtnmHCLimUR3G1bYdiFF0jZ8xwmL13Uyck
mTHdVgnc9RdXPrk5JfqcTXAKYpFpO1gHe2Xgx8zRub0YM/BaVftTxq0tpfOkfDBQekOfYfXPKmAe
NpmNaZvc3w1Mf8nOlygNLwqAR9u5ubJtuNA7nYFDEmmnjSfrlcla/BB+hoPc8Jde/0IfnQeyDnd9
pg7Jj1vZW8UhulvH77WIL/2zgbgsgn/Pcjd2tnhsqO+M2XhDGhQbqBLtx3C1rD35w6HTMglbLMMT
QehW5jzWFeZaIeDES+Qaubd2QpEQz3/07iaL6Vbbv16+TTOlc9x7ZuBhdz+2lMqcfQL97t3cnNYN
QxNFqWeRowzK66/ZBHZdmzpAtE+u5DHYOfACTcg0k/4GgkvOa9iBHh5cEiYxysId8OnOJTnR8700
XufEsQcUX/RKxbEQr1FSc3MIvtOVLA4rtf0Br9nYKxjBhbWm+nstE8yTBKzAm17HjHuljhZzedet
PNuU3ilH1m4LwGhoBcScuaXBczYgpqfzND6vTzEyTaAYLtuJXaC6uY96MdB4TcQkWbkS3r/WO0lh
a11wuHfKsnL7g4nlU70kH9vuXa5IV7kBb4I2VT0Iz4K8rEyNvUdsnLEmJLHwf1IMvrQduxBT4Zu4
vvyhXXIHCnx5A+tb1hmPYVvDwuSqTcBHKSKHRISONDCJ3iECf8DAEm8Vk+MEqGrOkGJprrxXx8/u
Yx25VDPbVySEhToBlMhzdd5VggRRsatLsGtzUndWmhLEts4XNAf2x77Sy5RNFgr+GeBtwbunWLO5
MiMX7eJxw9YrtMZiwaX2e0ElndWM5gumwHsEMXB7tNfaO6dCodE3MXtsDJ7/2V9oS+rVg1J6er/j
vErSh392uMOZ1+ny/TVXZuG02o+eQ3LQq1I8GhmRPzr+RB0N/oyUACjCrvoAXjMu8uvVjwpU05s0
jnbF4FM4NoCqCtsMLuAKvUuiuj7ojIJdPprlSWyNRf16gzdJqCwQcK43Eve8KDeuQi/WGaLtoEQm
1BrWSm7ZS94PlSzBDtDQ5vL+J+RiExCBKLuuuN9o8S1Rjw7Z3H3gvV8zo2T22zf4h44Vy+QrsuH0
0OQ/wcY34Obyf++sUy3HX6ELr52QDvwRILdiFXdvUxM6RaYuc/Xg/G7ANp0koezxZNvEwE+Njd2d
8ms+FmjNBicMwVdEdtc/hZqd4+Y9iaFh6jw1xeHvKvoZSF5OYRywrPT0Ora/UTPFhWOZilAIOyTI
bxvWiNc1rC2pGBHXF5qGP3WEh+QoqH3+dIodaV7c4u7WHye6PWVTgtvcsEB0un5nbg8TJvrVcJkh
tdgCxMEdgnjPaWrfoNYAlFnc5yRa+4WUKaou+Bc3hcmn7kXla+m7luagvMgjxoWxO1fMDzYNB3DE
uDdnqrnnlUpXBkNB3IUQ1gP50279hP97kcs88iwigFi8DWKnFuk88QJQE0rW+2L94yfyw0ST+TrS
4pPtkOOAeDMim0+LorvF0RRS/kxgJ/JBAA5iz5gf7B4JKJq2rvwATHfwxANDJ3OkRGIZ2UxhBxu2
SPKMIi2ipi6VyNJnWwiEpT18wpJSXA22MD5MuZtLQKojZDY4smYXbOSQ1ZtNVGXsg7FewVr8fBck
FroJi/a+CxWlMHEgjzXqyX/Tw2edDEfTyw2ce1TjNYuT3VODRhihOgiU7fbWLRUvE/n7ACZxU9DC
ACnibz/KIn4EWNhCNowCiyBbCfghKgORfK8IsS1Kek6d/aaHp/dpxVt4cqHwB2n0o6cCL4N4S0IL
s9U7o9R5e9cWYLP8pog06s0Wd9LBV1EYzPsqhs+4Xxvve/nBwuLhqbLOjXA62lPv3iceq/0qYmIc
hNxDUVoMznvyOtup4KrGT/Wd/lS68zEszu5xfkr4FzeJn1vH2PS0TJcXiFroV03eIzAFHSBgmZyi
U9NKGvb4CIT++yZJoiELmmQ1+xwMAyqR17EDFM+Sik0QqqkpumurzBXyJ5BkTYgWoAUrrOb7EIR6
4y069kxWWGLFI/WYqNPuilahp+GheE43IrJICbuJHyCGxeevic9FWvtr5LxF/Vyvym039PHi0U9l
zC6oYXP+48TBUZJ35Cdf4U1/CLvwA1sehHwIpilspwqowZ3NoHD28fq7WazDe3om4hyh4WvOeKNJ
5PY+0QoExHNFJ088dUbhvE2W8q7HM2Lh69Fb7E6hiEJXoK0JRtyjhFrAGSmZvczI35QdFJllQh9B
qoZT8bDdpbkcMN6vuN/QYUZiEDHVD45hNTx8gbV95kRMnLU4XcsblJlLiQZjKA5hnH8ko0jHBokl
AlAg56kPknaXAY5qGCt3jn4knthrluGDBysHDoyLfqF7l/ApO7fQpHJJfegg0P+Ep7rr3+5gEV6Y
i76O4xcKY+5zCzzrqXNyvstsaFnXvc0rhX8GbAtcb0V940Dy4KOtk9dWCk6BT/R9SuSTisp7wHMU
BC8OG/U8Twwo4IEuEa5pH3U9j/Rx+Pc4uY9lQPBH49qANFN6sjqU6iltdACVL4iNNqS0AH6HZWKX
7BXOFnhAk8XInI8iqiOOyJoV3h9b6vW6+7rweravU0Zd6CC14Gmz3EO6JZkp53OeuRG/9vFEhtRt
21TcP8Urz/NIaLIaVsCShr+1sLQc9UWQbj47n3EKbhVLXtmkRkJ3ZyOHvIj8PFrYPDoNE3sACefR
TsocW2tUhXfTAMdk9pnXnf/cdfkSprMt6nSqr6wlbM4b4nxhC9umHVsRm7TkDfi4hwtJh+t6+eqw
5r2Yk+ju+d5jU6PEPnx3oXqmojElnerHMzzlNMQ6FlUqSxusEzNUEU9mj9NMsDeOxGw+cm2wwg8q
GVeBsrYyy+BBCfejK7huJ52RAY47W8yNcB/E/E6b6lKX/3BVZOA3s5ErVrqc1eNUk2USGY72enql
J9uwqLxbLVpwVNGSxCqIhBDow3wxzSagOz1gPkHGCbNSNBm0BK94PfUXHzn82tlbsR0s0HqsTLax
8jfYNpRAU0rqh7pcmUET7/XPZo1ueXQk6fBwPV/Crb/+uaU2uH8q3g1TAlBIDZRG3ZqHX45+wct+
9HmX4/sw/hQWiuCbwb3r3VVusHlzCgP83/TDbD7WpA5gfE5HEPLWZWB9ebpkEcyHqNJURT23Qxd7
iiHGJyIyNnsGiS9kUHtlInYSSnH6Wwj66yyj4qZriW1a6PA8thTVHPae81AO+QSmunSc7DP4SQxV
ostVu4oIEgc6DjeoQZJ4+coC1TtYq9ivTxdcxxBoKnFWG4IE7Y+B7Xwt1TB/5TRX+lKpt06Un6i7
g5pIG7YhXHutpq5r7BylCBiFX5oTbpXlYVAkvBQWLnc6d2KqMkJusHHWoxBMAk8wAeMpYYokeC5j
EpH6qVn8CPNZlIuOOj3kCzunMtg78j5b+NXDoc2V1Sb7PnJT3yB1OWAH4zRjegYHBbwMMvgIsgFS
telCyQjzXU5T4FBg84kPpnIEo5xiIC4b+J7jtotNW6DMiAQ8vuVNRhOFxxKHRzgcwZ25FiAZ2qGF
fE3wBCMQOr8WLtRnfQ2H645TrCs5W2SJ+BYRA7f+tmjf2KuBzvIsOuw9bWwWFWNSCynoWbrkSREz
PUeqXo6JL1EppXaoLBhwSeugvzhIK5y7ACcNF8l1H55cBMejqvTHa+EuO5/4Fqt0DOyTIFg1JVU9
sA3Hre/ZqWGzpIfdevlCb+OoYoUfUMDwbqcNNYbG2pFdTH9yo1WUUXszCeW4UnrTfD+qqEsjZjpw
LaqgYQkK3AGuofUdFQP3nXzlV5VaBQu0sDYqKmb+sI4mN9dvMgKzqWM1idc//bns6MNsc8sklL6J
Muq0g1XZamLVxkwCbNGyixRerh2tV+8yas19UKjsf6aA8zoTg1l5OFBcwaWtckbrvHyL7cKvlzHH
rYn4cRFDsLOsw/6XLggIvFIS724fTBX2ba2+VS16A9+t96lMKQI1NdEXZWK6waz5BiKqalrGsv/D
DsnpOQj+PdmkGGxsD8o3sAey7fxVR/gkuN1Ch3T6wcrOeOQhOnz8NQgakMTl5f9gKeFnx6EWA5Da
FkSqXFZch42JeU5s7thb9xXqa6JC+HQuVfSjjlhkvQ0Fv5RzIcCOMjhakUg0tMjx5gmWsFsZ/kut
53+FsJhgJheQyBP3J8sKgX54eiCKww/KyP7pZapSd4u9yYpEKp+gkZhmOC4biIbHPMnk3X/qzyop
CV7KlEpGTIW80w5x5uUZlEW88KUY89DCK5zcdIQBoEfh2hHFF659FwYMrClhSP7xcB6c2sWblbaL
6j+thK30US/tyKlvbnVLo9NmZJipiRkg/+tfE8eKabnOlO2fBxOcRJGvpJYNs5KuXFpUKQV/bFqE
/U9DVF1JENty6BYXm7AWPfUD1WJoqzFhaUezlAJvMSNZeGfV5/u/06PosFpZ4YJbY+q7IlHAgul0
+yZTeqmMOKkLtdcaKQwrmfh/EYhGwisPY71+LRmQgx9+SpsmvUlEqWIjGvrQUdZkxAcfa0NuU94o
1PTqWBQC2rLsQeci0tnSm76c6uG7RGdrXROwpQg0+x8sK4hp2CpSnZ5jdP2IXCnVQt/dmiblrOyc
ZdVGI66xh+UUbT+8Ym7+czrjtpUodGOZNDKwTD+i5bHNNqjjxBNl+7aeBnPWAyMqd89cGDvhruC7
bNR3ld4omZvqUHhu7ataU6Bw3p7qPqzdVIcipZvc5JUBZ1OsHMbtdeqTewm5H/ZbCHUIY/Z73wTH
zVZKZoxfaw91vOjrRQELmhQT1CVBfIySupArLfJ+ckCMeF9D/XnC3oRibvb05wXFpty68otH52gY
wSFPVR048/hene/LP8jRXr3H7CVI9ow22vWAw51cDV30TsVtyTHuOxjXB9a6TlKk3+Zr0R1YF2ME
2ku8gQ4c7OzPZTxzX1Ib2VX1tSSC0OWVVaDxP3mAiesUCsYZCMYAe1tQHfYfoDvTdONmjF6xuY/e
cL7+aqrHlhUMei74YhbV74s9yFtqzu6tUVs6eruwLv8UiJERsuOyY/58q8ZqkVwMsEi3cOQPQgja
wOaYr0I3bFH0SLJ/mLsKbAgyFppAxdFxmSPvpX/0GBNY0RJru+BAEDbIlzIzSOJyfj3qUiBYWab2
w92JLh5h5EPJkiomwGETLeGyiU+qDO0QH2zYt69i/44UTDVCZSEjVrl9KIMPhQWwHhElU0hGWN7w
++Yj6LpTHAng++DpgjmJ17CyeI0rXRbkWuV+hrmt7wDjpLHw6CndKsy5H4fx4UG+I4wsnbbV+4Ge
TVwLDWzDYLCFZWjMl0lTEZtpIW/EBFhZxkas9Phxon15n/0YNzezLEP4ZmddEHuuV4BTOCoqnukK
xYnrzn7n6muG3d0h/xNaeHFzKfs7VfvqL7BQeDpdcdAdEWo51zdsM5W3cJnb0R4VJppP2yrLwr5J
tbmcypQvrtrgEms9haLOf51VHq0u7YzPxoWXg+/dYl+g9EZYKOD9OQ2sNg18aLi3P8mojArLiK1L
D2ulcUzBuI4Th/GA7D1+Kj3B05Ejc4HzlnIUl188wAb4V+sHONH9bX0m5xCrbC0hOwcdi48ACu8N
XTx80BJXtTE8Bw6dS1prVRy1lCl6bfVdnal5xiiHTiXJ3v7fH6gGBm/6vqpckH5LZk1txGi6pb5A
6imPHQ4TI1SMQaIL+PYId2MS0HuZ6HY5GGNpReLfog59FCkRklhi/WfbnbEriYVOfgE261D4hlR+
/fKVHHRHE01SJhEfuR9qqvVmJzku9jJlzyWfKsaq/RyKq0AgvT8hbyx/doG4+aSIVebCYHFuNhwa
NXZZEsDjtj6mmrRL6+8L1YRWbYQpMYnZhQhlnRo7Xj3Zx0Xzeu06pL9wXX2f/6s5Wn8tobBgBaAM
erwP2w2dfhq5B2dA9d7VrZt0e/LArbk7X2inzkLkEpZXiQ7rv6GyX77Q1C+rD37A0TFlBlfFfsPw
msKap7SxnZh9WYWUATIw7acq6tQmQuNSS6rAR9e2ElXlx7cNDgiKBpdA0hKOFKu+acxvGdL1tN6r
U8tMD2x3uiIRh2mycioBvDjE46bOCsa71HeEpAQ7Pqec24u3RgGqu2DZ0LkLu+69YkBP6vdOkbKj
8ljJ62n6KAKkEwTQpU3wMw5dNi8i0xJ9V9CAssdRWCj45NUKG1qdXXTu7a9Bn1ksmOOC91tNdkjN
RrUt2W2MSQ5WJ5sfi+WK8u6WfPMVFU2LsSRj75mbXv3HMEgBy5dU/qUCMA+yu7QPThG+OOv4n9R5
Ji2NnKubIqWdI2sdFC+Y4Bky+txB0STTnk/4IIMt7HFqr/IlocixM4NHyYRH/4m9JkZ7ZFatMeV0
7VRj+qIVg9crP/ONRtout11WLI/GvSVwiHnksCe3mESH21tcYCGy+xkMiti6FhiFSyADzQh30lx9
BeeJemo9I5/1PBrWHvh6CW2xB3taPglFSzDR5Kl5jLWasHfIIxXlYBUGUgaHbgbQfqYKUSbmHxr9
OmGHhbvCxkYXEexZpnKYD2tjYKYVsXu8txsGr2QkGJegjdxedhB3ZiUeOYJLWHQsKXJ0AftqXokx
fxB/V0jC/QIWh/NnrMG6VJU4/7jeKiz/IdmsRuqZe2nZSnAnbqTw1SGrqRidwohfqbRnoEsHwGWx
GsUgt4HoIgts3eMi/H8nhRSRXyiQGROtO+061SMwpEmkO8aXtNCCQEORgPdfR6GnQdpgnOy8v6Ho
Gv+2WrRWu7oT1tfUQrd6J9fcdygiXJN9z3AzVR7T3ancnjsnVGcM3BxxMqXLSwa/daGHetE/IcF0
H3GTDSJbM3DWJC34wUsrcO2YJEs8Q49jDlPnem9WHq4Xc/UC61x7xiLdhQ/r1q9arCjPylcLx021
zCtq+xQiFpWOufuEcqKfC8QauvfTk0iAMEez4UVK2VFfBs2/FJ246DVR3xRVSN6Q9KNUE/8awu4S
fm6A93Dz5drg3sJrY0m2XesrS/ZvTrG+rOzfcSh0zsFVPeTutNprDMIHmbgP6Oq5docKKsVEv+IO
PfXCWURlywjckvHLoHKD8tWxKdRa1khVqCXJ4K+rsvA/tXZ/WsSIY7IrduIOB2wnLVYI/SiZolc/
/Fh0jxtyfvUPLIIXadtg5wfW/AyNy5H8hVJSLm7ZkqSbd4gjjyDW9zNmqh16QHOsiQ80TTq+w/Mq
bupZ0S7hxEUR3TPqJ+HWm33dqjf1nxYAx4V0KmsAc2HTApjNkHZZMxJzrM5wW6nh8frbfnotNXpt
55jgb5H2XHBkAUhLZVx+208aSc8irWEKVpWWrNJjttQIA+QzoLkywstY5aXp2ogKxXOgPT3Bnn88
C5nUqGYM2SFCB3/e0ARonktyx+iW6nGVP85gj8r+3s1zVV4K8YPKK3an4JGkx8Bvw/2XhLOCCBIY
oXBJyu3/GYrulIPipJzoWDTXj8yQ3Huo+A6vUJmbyT8+RetExv1FHW62KrODL7nYq2h56Ls2d/Ah
B+Sjn90DGbSQ2wsQG/VhSnA3Fw0roOmMHCuNa74nc10s1HpdJaVBW3pW6RBRfj0ajVThp/ImRr2k
N062h8YfGfmDUEPgOZ1UKOXKj8rPc1p+g6VBSKJuI5dC9lgV7bMMFUPWFbM07xm+zBoqHi7C6DmM
vk12y0zEGWpA/gNrl9TDjSFhKiax5twlLr+z+BeHXhiS4GPTRBcRmbqM019ca3OLBdGs1MFHwa8I
bMp3q7m4dyGElxRsEkVISLXD9nm1xVF/mJD0wNR34T2nuSu/VQmtG42Vy0VoTGA4WNmVqdPyn3u0
Pe8WIV7AWyLGch8xuyt6CP3I+cYC1iMnz0f8DgdupnY1xr1o7cWDiqiwKWwaodRruN3dZHAy2EoF
uElq/WFiYm8JE6f5fTmWl0DinoTWi+dJwIY3+utwOlqGfs3AP75ZpGZNDj38uXYA4HTixPajr1yW
NcYIJabr7r9zF5w+EibBUQdpFzO2YcG2o+cfbyTjhXC1jtDimdRSvjk6w+BOzG3MeCLMpBJK9wLY
y76cXmElzs1az9N0IzUPHU1EoM3X4fb30BhM6e16jlDTA0TUVTZLtGzkgzJ8peRce2X8gAYTLUz+
9ak8tgOOYOvzTOD3Clx6IKEiZqRceIiCeAact0tPTTsQorT07ljUJgESrTk389BP0bYhdBdubd6X
PwGySrqR02s8dKBWO1SljSLJQE/5an9aQppzoZP6g7g3TBjsEJL4B2ZJe7A/PNf1kk78x2/vLJ9N
pVqNxScKAFP1Yb9GzswKxjfy4M9bkLWqi7MHzqdF9un8E4E5fAaRnnmSCLRq+72l2Wb2CUDeLSDD
GusyQs4Kj7TG/H1Lj2K51/6UZ2L9gFp09/okwHQYyBakjceS1tZxe9sF5tFB2kAwZ7n0Py0Ad3n4
IuQ4mEVlMTXFlMvfc3R7/yeAyCo42lWgyH9hTxG0wB3XfXj2l1fILpffcAfJ7ce/oc7GYuoxckFn
DOt66aQzpMJhxQpPH6/ww6YzGSkam1Vt5Lna2kSIgKe3nx+k6btVCwtvi73QJDeJTYs/q36BI8V1
lKPoT9dg+nlXu5Wk6AVW4w2ELGdu/EDqaqiU0q2wJ+xAq2KXKdFIF3NdW//K38WLYRj5M23pIwkp
qBKbponG3za8vuS0McVlYd+eo6f20M0bK49bE0nJsHGaE5RGEVXMVh10/chnfjfa2KjZtzZ9RAdT
anTwMHYiyjkX4OzRkSspj5vDuCIiClPkOlpiojuLsaMzmB9e03+Yh4nmIa939X1jNu3mH7jGu7Zr
HDiyuVfLS+dCAm19FrBDtNNFMwSwh2YU9CKU1XXf1TLnJvy5ecGl14Frs+uzLuAy+mEMy+nNPz6t
CX74Z0Z17+i+A7WUGud4qHwGkdHkjJRS1DwyniTjt4yomnn41i6m6WDvhmIwPEAL1tK+4X1thMKO
UMOvwKi670z5wAAuwff/hUv/ySt1uZkriwtocTaemdifIv5gwSioqMg/kDSDbkt5tygzQtPc/El8
Gx9FwzupDmR8nVW4rydYsUVnQmJsVscXzO/gRB6EtHWgZhKs+CO8ek18lpw+Ltq19fkKgSjDNBWP
y3edPx+SHrJz0zw+Xp2MNk3zK3dY5ms+ubSmxrdJ7ZivEA0siRXeu6bm5OaWVi9g2kan3blSIZMd
kxnJJegIDnG/7QLfJVZNLNU4lk2CklPU/BrM/gUZPZavbta7ura/o80rvYuxdPmTznXwK+PVAlPG
+xrJjiiq9ETnXfGIj18fVTAwLiIKn8UvGoTM5ojKe2aqR1tjXkBV3/uky1l44PhG61NRxy9NJ8gH
oToi9zwq+lvB/qhUHN4ZsQTQk31woAU5DgThwR1PmKmWdL9xHdRM/s1N3YlLEzWva25r+oM3Bfxm
r4J7jYfr/rT6QZ3drZUd0RJ3alsuYbAqTU6Famb9hsMY/L9KLrGAJ15wTSdhZEzwVaXQjzM2ah6a
Swu0sqCRlul77EIjJUJpLdM5aR0hfiqdVG3w+SrotpfpAJL6VtfzWol4D7El4auIuPskvZ3u7/mg
zghYB4HE5gkvrSQ0dF6qysRMLYGBTN6sXtq8A9DyvWZS1gkUV0lW/olUukrlBF2PGnBUt/kG+1mP
R6B8DVhNnpi5az1Vhlma+ZUFcvK3c/BN/Gfa8Bsf7RBfQyfeyXjV+vev3HRJHCzGgJJI0u4gtX1B
ZreieUx1fgxpkw4Zg+dQAu8ZGy5Biaw7agve69UpC5znQ1sA7uEVL+CSF+D4l62RxfsJY3BD32Oe
XbzY+BLPEvbjz0/LH093jZDnUCe6s4//b0TD0Yl+S0OQaW8DfB1joFncDHVApbfuo4738qXwMjo6
Lh4/YvYi5CIYrcvNpTfC7iyAiTPkj4qhsxZPT1ILAxN0Sc+kIQJtADmPKIdUq5h2YXRAN4znNYRv
STcDLPnlBqVc6Ic45H92UpVfhf1orHjaRViChAPXZ4T4A/E4wAaNAIhY66R8WZTnW/31rKG5K1ny
QTil96UiOFru8eH1K3ghf83NuzVhf6oJ76q9+4drqZOu8xHHN5RPw23c/ltLqV4c9LuFRWJYnh2I
lE4T5jc6sZzSwkIV14ts/m27M/DaDY0yaAklDJJnSNT0k81Tt4c2/D+6RC/t7u5/IcDugYZ0pX7h
TZya0nKYgsEID/tSZpV0Dy2V+kef1kv1atgTWXJCwVcAgc1gj3khFR/19xvySneFg0PRJugcPlUA
XB5XoDE93oFcDTJRQ1HO/+Ll+UeM+9l4O1XW+16Jhx+0TGP1K/8DQE8iXIzx9ONln1o90tQ6NcuB
WTq6kcIOF2InJdCqju4qotQaUJNEwslMqaapYIz83nJnJmi+cpTkcFUcrBqw0jzvUcMyRPzYEpfO
wrb+t1aBFHb8wVwjSaEKwkAnznX+haAIBcJSEzGPaKGOxEkFN9byJec2BVAVLROPaDuBgdAQBcD7
lwuXPpYs4VXRkZuiX/3Y7pjLLPQwJsR6xcljQK4y34rfiw8LBZlXIVFRMaxL9yBY6hgTQZmYFfqu
Kd/vLCOoa6m3DILVm02uyED6gZLpaM6Se/CLKsbDnoEhZk2tfZLjZP+S9WSP0Um1l7CMULnGMC0N
YTAtKxp2Mva7Z+w1xD7Kkm7SScCKJeNbVbXV0HaB/nWNFkREclzGjQYoEwrFYOlBJIo/LS+Xwi4t
ItEc47uOzR3K7UPr8V6RGSd4bkzYVCyOtvSSZp2gnp7paL0rfnZzvyXqaNfI/PAe9aZgFrRZGQ8B
hwZYh060Pv1/bbRtUDnTV89/SFE8q1jc5R6n9S/IA7gADQkJq4WRO7ugETh2NkDksfa4Vbob3V9t
MUMLAbzlHSBT7RBrKNXetqRUphwMhIVT9/j/PVhirfFw77Av1v5T/lTPXGWPy/ux5Agd1hNhp0pd
Iu3ZMwkekpqgwiFyPArPhPWTd6XW82T5akC90jcZrIf7Y4M7nu9KKqnVUTVXu/joAfrcj0YAA8rF
NlgX6CaaHJKUSDoEbh88RyURkG4YUdFffDDrg5I/Avk/5AwtG3haSwFhebQ7K8apsonO5Offmabz
yCee6kdFsdB7K1ndCuaomrad5pzbf2ju6ksFGPMh6qRzKw6Wi9xQlmeEIFMATj+oW+osp0wMbnhy
ZXNe4zvDckdZtJUPgaObnvbOvSCOtmwhvSCidiU+ca+v32vdAp5zvSh5cAGxrYX7weW0fTy9m2h1
Svp8PhyTShWS8WMJGyHtcJtJE/vMAIevUp/OKBWqFa0uKy0/rzFx34oIcTrEHpgWPCteaOjZKuSM
rVVR1vUyIp0RyGE9WgkQqWmm9YyqA32Xk84LE6MbuQojNNYzZmRsCc8Q4qAJ9RpHfQUNuRQEAfjh
+hH0mCZE0dbZHBz9W+86RdDSt8uvhNOblh3hyq+Wyh+Ae3JSlUajy7edKxzx/K/O4zf323naEc+9
hKbY4MsBM8rgFCXOumlfRI68Fdu1kp6kSeN9JkWJFN+gVmaNHLvtUX/hXglRVP3A6FNfyb4ekT33
o4r5sEtaWkKpG4utRCX5vw8gcYLeCGGWVS9dCgC9mWNPL9hsmzMYvIVf9G9sP3FLfEOYrqr+zXZn
X7tX55rRHxgpQTUjcQ9TBm8v+G+XQVe8iO3WeffBiKmbVmnFxlHqzP557EReEqLNgJUa5zPLqzB6
Do0CnmfNYFL1+CslUqcG/ynFypfJcwLXY7Azd8gOwo/O57Yhvjz+XFlOFRYMzSqvWChuPd9qdYxu
ohWUKl0KnqXFTzlX8htuE/kro6gai1kkVEtRYJff4S+RDvZaZltSuADsZ0d0j3Vm15DuUZTB/s4t
FUfOYablmCjGa26fwsx0PverqG8nDISwqlNWfQX2bANs9xQtLEm04bT8pbLa//7u0SL8NlDFXX0f
Y8ow7q6dv8l64KotXs7SuAZHqPn+m/NcCZwDsxBq4aeHcEIS1SLFHfsbM7oDFm9+ozA6nDjf5PgJ
WpMoixI0tndFDfOd3vuwbinQDDxuzir4ruWhxZXrTyRNNG2pzriBoqOV881+o+boajZKMM7iFPN/
TsacE2O4LntxVlEDKMQpWBvmyjgmBwMkHLO/AKtOaMw7DpV1yiKw331IO+hOz9wmnlWsXyIG7VVh
GLsd9X8wqm7RhXlRgqHuHLyBoWJVilH4rXwbUrSghe7EJNUvj/lnLhyThLrsk1O6RFH92ABznrtt
5QGcRYYP5kyXpyScL+c1PrsUXAYQyEJHJPSQhxY56HoQ4jdlfJeqrBSKlrRz9xKv/CNrc3fZZmYc
d/fjBB3jq1ZtwJ0VETvVtoEDDWmeh2foRKqpQaQocEZj28FE/KIGnMf2JjyU2U2W69NxdTRwCoHm
gyucXMqQPE4lBNoB1zwUFYdYITjm9YY9vLOKH4QJBV96nIaKqwR3LLWsb/+PtmHJvJ0Xn3Dh6mkU
X/VDUq9WurM7R77k2vyyrfsD1hGWKOXhJ75MRfhp5ydortGFkmyjCX5UMNsbR5fZalGT+9xCoVF1
MsI0sLLQVXKxHccqtx9nw4YUrueJPR1tZSkOJQNtf4m9nBLPHcnGOl9JfPgmHe8rH955clyFH4H1
hsFIz8uSGlw+mHc176BuceO9aFfr8mhuMB2xDTCOkkhEWt5VzlEOxOC8P505qjGAF+MEYFYlQKwx
iboRipE6FJTg9npb8qo0BeTtNjJ8ICY6j3vWDOKYb6tCxS89TbAVqxR7rPcPpDMQZ8XEVdItAaem
X/JnKSGROFkEPn7ahw+Y20V9s5fftpRHOH+HabG0Pm6s8OgkcUo4oXrwa/wfNaprakqcj765PsUH
s0VhAEue4Emq9Pucku3LqaJvhWyTho7KxLzs1pG23RTXfdeu05Ux5p/3HiSkW/naOSyfiFq4swOe
QYyGmq+vXSvLTXnfODNIML1BJkheMeE7FPyvJyTvDk+XzagkqHjclQ8/x2pfaDTLi8+Ke0AKGuQL
ELmP54MdeQtbxsI+5l4lZQa26SPJeevuazZ9bRH/KDn9L0aL5FZSNx5TvugTD1rq20TwRXswl5Rr
3D4gA14pj3hDc+Kzab5MGlZLe+wnhrqsJc7sKd2yYH1Ii5uGJ81gpuhf70Sm/rQ6lgMS4mGTxyGI
HsMuvLfg2J2z5Z/Gi6J+OqTtWaHzvJYpptVsViK7seMiiMDMFAr8zoxaGNqQbN/ejEEjrKYq8Pl0
5CtYHcle4tHLclSSgO03/1Jav7Tw58MPTj9QwuMzs14KBkVqoWX2LNcYGPWm05RhGuiCloCASB02
k6HoEZALSQwyQNtCqvhEahqXN+FNgRKubCQDVDcIqgSBBckncHP5Oc+P1NuE2geNSwm1mD2ignRg
MKtX3pCPL11kMNlWAevPACcvbZiK1AbSquqpbLDxXCKAR0oLYbLZFfuHU+/W93TasRumYwGl7toz
FPZBBKswstxsvwRUmWT7tYR5RuDt0SaUI5D1YwW8R623If0XGlvnsNFePzDMd4LtR3RgNgnTZaM4
ut9++OLD1FG9scgigJ2DD8mVIi8lPxV6XU2b3dI5XLD9mMYb5Cb8pRqixWQTml3/ni/54K3BkHXz
MgjvaDkizaFPSv7sSo5yBduBSJLRLt91XsOYcKuRjTNhgzBdUoUXTrXnfX1zx3s4nQgBIcLylZWf
jKG7uoNiwm7BzR3ZcFXl6Dwjf7WymvrYs1iutrXz7lsxgfdwx4AqkvV5WEa7747tndYimprLexRb
ZUs4c0qhvbmC78CnTMRsuEB5GfJRO85vYviJmpsZ/UMAPA4GeVF6CyjGpPzoeWiL2wdx9SdPEgcm
BNDwDNxY++r5SgLqk43gtkiEIsQCVd0kF5HuqHzWb/65DQzvElJMmXXfhHGwJvjsdPy90pC7Xs5r
jBT8uS8zep9IEqCsFiO545Gfve40sh+5DLNeaZoNl9WaSyC30WTAYyLggNCC+QCqz2Z3ObiXEPV7
9bBW55R99JAOL3m7tragY0RG2uF+Z6PzlFgs15XlopdLNWBQ/avQnQmahz2c0QyV0Fsyjf0gy2OU
oDnWiedOapVNdAguMcZA5bOi/7PJbP+eGlOCMXwcglMUoCVqQHl3H46s9iqmIKO/N4VheVIzIliH
xeQx9X+QNm59MyjjAR0eKWgGnpp+sCPJB16OoUtftfbr0ZOnmTcep8Xk638ps8YyaN9dVSm0Hu/8
aLtfGUndcr6Tf4xJ18kZmORvHMuchHL5zkiVx4l2cmo2BEPX9pUu+lztMkbAGmaZ6MJTIiW93jFA
pbbSJ5IgpHhTeH0dQVud8vju68MmwV4L0wYfHLIgwkRE1Gge01B0WsJjWhruk6N3AkR8F3o+nqDY
nLqgEEdj6aYbQiXHuZhoFDEXWv6rvYXaIEMLedjW3NA/IQmIjYccgZq6Dh3OHSQf8WBA5VOszD24
mwnUhgKabmzJ99yg41wlZGn9g3f9ngQUrWt58H7P0au5Xl2Dpu0SsOJQ165sBZ+T9h6mfReLkP+f
c7Br24Con4pSjLsCqzYjk1gTiUMeLz4k8tKlEEj1zTg6J8X9i5oirgMUm7MTlaw1jsbz98QKC9U2
cCGqygRqpfcfWb1ichjtqUiE1YbqLaizxsnjllTDamemb78WUNkrRIxVIMPQd0NckxXfV3YHv5aQ
eGXN4Q4++bWVAc+FMIag9Qa5RoxyhF2sWqbVgp2PsAbHBGT+ARfHt0h8Hv/sivD6gcJhQzLKiJWk
fSDJSeDucRsN78IBDueslV+HBLehP57KkfaxU8zFlVcX7SE5jBRfB1eAuSXLfuxfO4+2XMJKxDcN
6eMVB9mixBMTkxRsC2/9RctmQOfvM9TP6C/XXtGIk/o3eQ+TnWN/0H5Ytjyn/1Zv7XufnSn2J5T0
Xs0gN0/fC0RXE1o7RBPLFWHQz14uFe8o3Cko93Pt+lZfn0Xdsthec1aDLLpNwp/0+MBbynSlyHER
1bogKQatuN7/Mxi3DDSlESMIChzFN2+TBPmhLxQGL2apih0WieSwUqzqfkvT1o3/6yAF4MWlZr9t
GExntrPZ4LhwoYq56NU/G8v7zO3pSeQspq6OUM8Hq6dssisy4wwRey33OA5N5QghyDAhi/azSnzR
sgagpU2obB3C5RK30VDFX+QglWNAS2Ivc/QhXhK8TXDttJe0CFdHPCf0JSqfTr2wFy1BUqu8hpCD
JnVS0QeCA89o2iynFQPBzS/GKjDzsv0NfHiQSa6tjI5+wNuZ3jCeWX88713HQV7DpEla0Iw3F4GX
NIvpA/5NjXJPpudxWrYAI+ayKQupnRT1B8xKfcoww9z5yCRFuc3NfhGF9BA+aLFK9dkD/IFlCPUB
C4wL6uvvS5g/hSuvHnpdzNvnN9hLFX6xFYz7XiAH2OivGr2iMp3v2AN2VgE8dhLKGO+QdOybwR+p
x11T8MFm13C4cZFGWLWTm3nqKwgZy2/AWW0f5G3/nfV7Ldmo/MzD/axmtKAaDvbvrEAaN8Ra2Djq
eAGYAY40UO2AUMpuu3t0f5H8W0UCIB/WtIoXD1/4K0G9BzUajcREGXA9YO0Z0NwMQPNQAil6y2ps
r8c6wPPEXpE3+tN+ddA3AzqKqe/YUNzorcaq4pbDaLyoMXOuqINYerRdBNwiUEa15MuRDUtCVEME
h0is7SYEw7bPvK4wsMhh823wsdg9tjrBrmH1Ab73swuIZcM6wZpcW2Ng+9bQRM6OAdWmvIXqybQT
nGBrKU8q3plKH/QsbDKvqtqdIt1AVGMTL2cTK/btOr6G9EtZK3PVN4l3uIHZEEq/gLLZSEN/u9Nn
cX9PAk6KBi2hfWEtqWNTb+ur+NTXHXdOHlvbVXJDlmaeBfpxbL4SG0J4+MXMqAj+7Dz4vS8rxTKD
kIiSTRCamfLy0W8wm9s+K8WAd3xt2DzPwssCZ8wKZSFI8khL1pU9bS/gDBNNhKLIG3PKY6Q9+YmI
PsN7tGvcbii9w54EPzI0JXndFEtoAwmwHkhX1L3MMo3x9Oc9bla6RcuHzrBapZ4iSW/bIAoaSIvn
plj1XPqvwnMIucZnwXsBVm9C7X07KHZUuagwv6zrfKKhn9hSJzdMAZtX4UpxfMsZn0mVJOXum4vk
KwKcy9Gt7d4Oq/FmQkdJlMc7fpUTJIbqSfVsH6BFqQ0J9/3Kvu9xZc7CRIuwY8sD8k3xbrL8dO1f
QO2ZxKwcpfqt9M8Is4ZAaEX7kO9oXA/B+NSS65IH44E2i4dc8O6UjX97DbaqqsiGprjw9DN8ju4f
HDWiQHZCkzri/lGgcSUdb6YUlbUeCZXbwuBhdB7gj07E+aGAuaakrcRFFsl/SFdoKm2INZWtZgOh
8UjoFL30egXZMo6lZO3KhK7AEJD0PNtRBkvu+3F6LUkTDAMUDaX590rtEZ7zioeQZASXdOEjohL6
0FINmJ5euO75ifkINIx4RmSKqYKTWyZ0NXwfW06OQK1IYR0b22whs2a/teYKkg1/VAtc4g/1y/zz
04MGmYL08UwwNi5a5Fh8qFYXQ+rsfAyawWzyZ3Wjp3rzoHJFriFGZ6hFXKk+8DsTvZllL8wZH6Bj
uFEGg3g36KHa+jTzqsNNyKW48UTHC5TtotJK2fyv9QpQok3WJ+6VttMAFHHEz3u2fbZ79sv/Tc2m
jxjoPO+50YQpeP0pJdMghtyzl3fzcy4Dwqa8qcd43FHuExeLMAM2zaoH0NwO8qoBzvGlF2Ik3Mou
z7fU2bnbEVlkonpoPZqgHvzHo7BbKeTFpC4Aw6PJMmI9zpNpK5e4bO7yBvGOC6tV76gESD2mQiR5
m22oYgyelLUgEXMC9XWyF6rymZLFqAkMCNctlTyppiDKu3L0uecTbuL8ApTdVbZTLIU/GUeg18tv
+jp5BFYBeu4KLO/Kb6/rjKIupl3q1G9Ue8JLVvScvb5ickOhuEu7s8s6vJaC1Sh3V/VhLejfQuGI
NgHhWzcdKrbbSihMl9o9LZtl6MTHkDbb/rA40fW1GtFikjEbrIc3ghp9rtFuN+z7VzyOQHpwKlv4
0pLZPkelROnSvg33h9DJE7fVotFzwuXnMTjhC9RrqYnZoOi6lWt5hKb7DOVk2FXJY65PFpW8tIbF
qIBQuqp1tsWpAvdtS00MPN9wjPgOjczC9WxDt+dKsOFUvEg3p20chvRWTE+zEfejTZGsdsKkSGHU
Mmdfyss7IrJoXkCNM3TEzqWaRc0cy20W+HPRDIr1mzZA7FMNLM9VjiMT+11/FurssTNqw+yjr40H
SqquAG0+fX2xw2JqJyD8Cyz6JlkUXKFurnbzS0ryBBUWtboxcdOEcUPnCM8HgDkdMGC2W51GmmfA
U/voMbniKlIEzzbxTy+TW5bP4BTXeFUFoavjQxGCH4NoF6Vd1pDOJ5obXq0b0krY1tFuMtxVMjRc
rNA81tisXlpgV+LatWmLQeUmzM+6ooqM3r4V5tjig/2COFuN105HnYlLCLTdOc4F4yYBrjlyiEA7
JRkTWgiCVu8tOIMJhXx9OCaaEMbPNmVCfIc+fCAnIzSsUTJE5ym41CXoYRJIXZ1gucKQCOZK32pG
lfNhByBpcerbCLVZTmNwf50h4whRVf3IedEBs7M10xYb4u6cAC7ncTgBch49TGJg5h923TjiZ3yj
vzfgE79DxNTCcnUX1Sk4eZJ3JwolQGQaC2Sb+J3jm/1qZlw7s1KaD8fEOl1ZR/6PMdQlH2QDIVTt
vmZvTbrg3Wdlf74hkMkqaAqkH5KxGhE/pOsNiCBdglMgZtWbWAyBdDe5vMf1VLZvJhWmY27+Qd3C
JueGxECk3m9p+GO89zFEAKmW4n1hvjhTBpVdmefxRS5gI8vKvWfGOqvI+xTv4088DbKP1wT2fQ2L
DXGJ1UJJ9R8FmDrB/JfHJwMfCRj+dpvWLBa9ibk07vX7UwYAuTF9aIMWDl7AdL3AqksX5gIWqeJF
+Tf4MKvvdkKk9EfsfqamdCt4rB6AlMjjUzURtejF2z6CS0hsBQFWEoo+q1sNCZsiI69xw0AzzyxZ
Zgux9l4KwiBevp3p9dfoCy+NCqQjm+cfwBprNr9KaEIova8FGCx5Pskeibd3xhirDs3SFVsNd+xi
GnSgeZP7vvdnbc61Ol+K07MUGLxll/TTec7sJeQUZWtgyypfRzWqHS9g1BFbxFg7qY17pK4K3pwS
9RAvlYzwLMN2b/HhTxqPoO9uh5sxBb0v5hYM/iCnGNvCbIzaYqtnWstej4tPY+xh104qA8XdrAlo
cNsiDN6J3xOfLPBDTUoD/+BKihxv+/OSsUTfCvtISZ/xe03P3c+gYpnyj4nTMltDoTk5qouhnntD
xiraILMAgzzchjnyI1n9DRn/Dy2kV/Fe2PrBWST23fgUrKjdhAj5Junq9atgkOSbI9QrQx5SEm69
p+q+Badqma82UO6AltB7Vab7Wzt8LkmUOWVGvf+ddB2T4F9vyCiJceIaZlA9C28aa3EEwQvlBHUp
OD0N1MnHzGs1f7xHyIzFy3dec/GBbl2UvCi9A7mW1HsShTrx2KKJxhPK8seCvHE9cBw6PewpkjpO
OlHU5LS5lTmNu/Rt6T+51unPWcvUAMtLU4jBRJeXeyoJhQoiFfmfaHIdSWfuG++EsxOL2tBoraw8
1lXT85sy+qR80/VDMPmn/rcG2b096DailwDInrl6DN1CLor4L2kbSmfdy5+EEB//2KLiJ10fA1fw
KDZwALfkC+dZLbwLgUkVMTQ0MwwrKK9R7TshcWrOw4+I8Kt4QqsPJBkvJWHMkLLzEkTWlN3ZhT/b
aDL2Tv26W6XTGTFclU3TiTgLiYH9FTcm7PaUilJVQ77q3N4tryO4uPK6GbBEthyZ4HK8JGKXO7YJ
f7N6aBTZH6+LyWi7SNwkew7Tonvky3P636l0nFWdP/dniEwBCQrPyPxrSCJTf+3bfPhMnHFNLjyk
CE3NxZPt9fnc+SEQ7l9fRJdCoiHxIhBD9BMo2fGP+nrFN8i/WKA8MdxS28qPwBfKv151iS2DnyjK
nNoWttc8bWs/SXRMmPUuemaNzSN+dDGlEsqL3Za47KmjYVOe4XCuQaOTj0UcA8ODV77ABkVNYpZQ
/1xEtzeFwsIWWfDIbb1XLyKFO0M3MPJrMRcHwA2NPkeIyvjFqZGyfO+KBmZ0mdwplfIWbLdX4HVW
WSANGoeF+UQh9LqSH3S3CKlFQrf+91wsGF5oXEU8rXPoWYoh0Yv32gEp4XxBu/tJZGcXwCwDIDPD
FzOKQcUNDeHNrsTeV6vGN46VML02vjnBq6ppklthGLRG/j/45CGAEu0yXAsbu1+TtM3XIByDjXzo
0LFfPkEOBMIuH13g6pNSo7HhfAUNXHKJVJvf9S08RKxn8Q+hgmhRjNPqsiqkcNceGzs4HeKScy65
6eUp9wT0ylF7TwtLca9uAVlBR/BN34zESS8IGTH9B07no8y0oLIltR95cgk2CzBftZg/b0lxbveV
v4UOZQfHorL+Q8ljJWPPdvj0GUcQ/6mTHvH1L3brQ+g2jUbmx3ViMAP2gTxGMnIBIq0GEtA8dR/b
bmn42vzf2aXRMjGw3x4EWoeWZpiVzVEFpkdjg+Jm2KulONx40BXCslW7SLz7XMxcrWu0uSej+vM8
5qkVrVpY+vWHGhzsgwq78KnIF8e9p4NWeaGBv/bQBw706fVySu+w+rk6sTCcx3sKAfZwHfkAR1cq
BgyBSMqaF2u/9bhv+XWc/s7fNNNeDw+6wro/aebOgikD7HU3nCF5t4d5RunCPu4VapNKW+8EYiJX
+R4uyeDiSbSVHro5JOYoFj/j95hkmNLKzX4T7I7bc7mpml/C+TKRbjxxBsXufBC2XK72lU3Q4USs
gbHrp2YepkJDm1aAYXpUPC7T/V5HQX4obmd4p2TqY+5p6dpYClTl4UwY5TTuXjMm4Uz4YGiP6Aq7
5u+LsyUcEGY4pRN6OIrQDWRFcNpKmge8DxToDSqne/rz9mWsStEKF+56E1LI6GQDlZPe2ITwFZbG
q7pSZUAt+cBsXCjeZVoyLa53ohYW2y0KxuyyLpTpfk++FoGZ5RKVie2tZi3kUQUc1r8cjitI9uTm
uufF1wz8gYgEk7qeDWqPZPYGLWIkRXIdQ/X4pO5osgO3K1OaktohqmJ7zmV2a9WkKfRrZ2rk1FZX
tFhL0JoJDn4AeVEfbYpuplI3p5SZXvWMG29kHGyzysh5x4iwUw3kszL8hed7v/StDUV6m2I1rzfo
Rzj5lG89PXFPw//tSLZK+1qzAYvGAfAbouFxJXZyGeqQ18Mh+wtfNIqQB4xIoWFEms+p4n50yJVP
JD9Uwgbho8GS15G+coNpXtheBDRyBZvAz+gflSaJiC3iY/2nHA+EXzRfYSzQAnuV9KmsiwhTyFh3
WNjpwGiKIj8uZlTCgiv1Qf0RVXIdgt3EYU0Ai0jfNpcoy/Byaww4+tEA5GSnAuA3cfX7tJzvw+KJ
pvWGB18PJ0JD1fXe6W1H0IWos84mpFCvIJgJHImT8pXJfIQ9+PTpiufd3rZvfG34TNRUu0vCYiY6
meHa83OWogiWVqrQ63BHOmCykYQVG+xOIigMu8NOABJIjSjKNIGqsBldbgR7+E9c5tafIKYOS3Cd
6QfgzJ5/qtA2kIJ8xjIGbT8OIc7TFmmiTGGi/Zh10M+uzlpDQHFjbYEVd5WPI5Jr96fCUxaLA2fs
Xjo6OZkVn85A6z42PXYLsDy7DWmoUbUP4wqRZ+34dlIgseLqrhoGld+YABeSgFk0RXY98V5P+mNn
ia+8JqIDUBf+go2k7OBtKq0NVrFguDQENq5bz9CEDIKHZBrrf/qgwjT/KfxF+sXpfwugQJfqZqAg
ixDU3nfEgGacURY6rd+q/zJj9pISmvrqm3v20ZcftVSNMDpMiCRuKG953Y239TCorkcVFw36372d
Jb+ksBnppyQHl0HzkLKbAb8mA4if3p3c+fPYb7xY9DdXkMnA1b/uQWF817En29k+nzdJLAzwje/u
hp+zmETEk6hyhCaJ3He0AiT5nt8Fgd1W06iZ3Hd0pLLy2ALGAROt/4BrT1278pacEG040QkHdn0N
10AFl8gUjB/19vp/BoAN1piy674a/1ntbNf5oZp1KDgIA2L2NffjG+FkosobCMpa4RG+BboTPlOU
6v4xiq26sCaaE0US465Xbis9MzN3+6PsKdUuLISMEsxa80S3ZkytBb9Ax1JdPv2wFDAnf5oRpu7V
MlZ0fO03wkJJeKpu5xEFc8WMQ6o/JQ1rKcNp+8xsoiGdGLuf9HEk8zsVL3Gf8G0T6p/SKAucAn1B
WZUAI4pWWvTIJTYfXbF2Xgjf7W6l1qkRvKHa5GPNayrUM8TTvtzPHNaIPDao0a+gX2eat+8C7A1M
PHAa5wS3QaVpFg4bUmZE6Iq/l6rczaR0GGSTQlIAC1evf6SDvX7fOrARyhi6XTBhTdUBMNWovKvy
cZlmAj0sTlfsJzKeGib6IENKzRNT81hvynzG54s2Kfs1taaVjlMOqLfWsvBjueYNw5gKwpxDySv9
cB5Lt+eEDqoWoVsfyYHZtHqO5yRAYYZmYKRvkDStpbjLm0rfJlrT22MUUl24QheJFRbBjLL2FrCF
vjp9mn0J2GipML6d9XUImdqGfSdacfSiQX2T36wOMARThAv2B0uto7Az/tQ6CHdMkF8V1xMgv6ch
BOOjWh3NHTT/ZatgqG7Q8n1XeAQkR69xNTGnRxN40+XgwbxybiNah/WCU44I2hk5YXJdDr6IKXwT
yrKBor24wHI7b1WajXveR8ovI16li9oRQ3fFy+//DLsWPO/rB2+35wCCAko9cd4GQuQIG6ElE5BY
+k/RBz0bUpNQOs33v4GfjtxhsEOFfmJlXzEJbDB3EOdmHSnuuFLeojWjBwQqSr/a7fjEq0ESc0vn
SwxBXU/2/WcZfJ5PEEDsNy/wrwmbfmTBnR7k3YNa0yjweA23fOmAoHZ+uJPKNeOQ+pVt5/p/oZsr
rnoCVolO7lCtPj7gVKbNiiqSUzfNv95qRl0YmQNdwSJ2SSYL1FAMmd651uq1IR8i2uRryh5OEw5l
V9f8OVrqMpyC0HSxNYwpKct5Xvu97fq0qO0A6Nhh0OnLQd4+qhImXNymGpjbdr+EPkK0il+arrQp
2jQ+J+uMqPxM5XqbswIwbqACkpUkdYiIfn2cNWK30FrqBxAiW7HSYy3UztMhxWiTHtZqd8MNMXuw
6NTsqPLJg0/jol3Yv053CGm6d09sAyt/XKPYvXp7P8xzJogIZ19FroVeRj4jpMIjsg4GttBjscJq
ob8jZ0nlciF7tCtRUk5oDIHqTMES0JpE6kJIMPiuTtalcCP+2cGBKxQas3g/iWNcPvfLF9lIG9Oo
49sV9qEYmcvBpWmuorKzJcDc0NN0+cD219UYaddVQzNxYB3HxF7sG0KFHK3jLGRcSL7gQudWxcrE
fOLKVMRrwzBBFHO54xAnvvjdvlTg71AGLO1WcpYlqkHUaDXkcaluNY+pt2xPoIrIt5x/blN75cC+
oUDb+e5KN7u7TAZfUAmFL/qZPL/Jp5Tl0eNhl17GCxJPVG7So8nRvTnGwXRK1aaKe77VezppCDsc
ykqXtXUay3PxqdfIQLKg3vGft/JSxYVFFb+kQT6pWGkRZbock6FV2byeZeHYuK+8/53usyQhA6g/
Bmms5fZF9L3X4IPp6RjRSaOI3o+chC+YxrB8AEST0cLpJP//9f7ocXHVLknfwsTYxwGg/UKaopup
/gNx4X//aQWDq6vWG3kXfActllZsOoyswTla8WFAqs9I09p8IcDSk3WkoLo9gn/kfvUFrtNUt2L0
eUCcd0eIKoJ6grmNSsHS/LaN+SHXV3dpEwpzqhqbrN0smSoZ6JzGX86J0Gs72O0305tc6WxGJr0U
m4Mi+JW1fLKlMXfPfTJTTBup5VEXgSDK/rcIwRWdu3c9uu7kMUppDPERXtB/5zJNqfxeR3iV8MEO
YXLudGgtmDSV6GFZAJHdPLgsZREi+viB0netkK/9yaoi5blyUpm2ZxfpbwpB99CRW34VK8QQvDLD
LQ77biwPmnZCEjV2LkORDlyvdLPIf+lc3aZK2HTRlYcnHfDkAdINuujgXc+lc280nzmjmLM2UsF6
a3jDrjmByNeITTbXrvtk9lkBapVDaQmT3Y8Jh7RK3TSfV8YfOJsRQfAo5zSNzsVuoecJtRcfOzhP
jOGM/33F+wXkptNHTH2U4uDWAAyaWPFY7Wuj2VHpXui0EMHfocpM5GfzyuQm3Pqm5MlHfegQ4vBi
S8ERa0KyYRbw4Tq5Ph/CqekXfLvn/6eS/hGmeZlRvnkARuSpG4Ck4vKBNNSTZQdtwO4yK+DqJKO3
qC5KceM/DXNn5xiOJ0HTFTqkndbwm8y4yNRyIahxcYpZYsa0judDucDR0EZg/LknoadCm8Oy2krA
orUndodwqJAB3UrDN/Z0NNTbWyHRH+x8Gu8inyAWzaKlcTnnDJUOd+H89Al1d+x0kQLqP11G67x+
V5FNi/t5+aJeF7UUvK23SgRwfqlKmdqZ4LOZL8ETWRjZ0bP8aYmhFeVt4gqxfypAuraWJqL2llL9
CRQ3Me+a1MuWHeGykhH5dn7RH85cCHrP3/8HJABDv9ZeP19jE3JjwJut/llj3vP6FhvorMd0u2Jd
tpO7YI5zmJFSzKqTXlBqEHGA1F3RD/yF0OgRiy2az7f4T9MXAQXdkEFafgqryXqo/e2kD7L0N4jx
2rV8hq/9WBSc3xHVrf0rcbHlmgQoFPUt9dV7eMXM3AuT2phBLlqzi2RwOqZNSON61tJiXnUR6kmF
j2Szc56HzX8h9+Iu8Y6BeJZTn+oXExvQGGEE6L2q1/03Ynhmc8mYShDu7EODHNWz78++dMv2H+bY
TZAZxocMi2PIOCX+VB8/oj1btMvOZOZ4EeoZ+Xh1nM3Yd/bO2oTFNSB135fJracNrqffhIamp0a4
ttrnSYb5dMItHTtT1P4efnMLGkYxaDdxycKsxsHADOSfSoFVA8n3mTtdB1aQxla4uLDHECz1XDez
nf7TD/3ii/q1RYbmeZ6nYVDUAc6NzoZyfafVP5zoU/oBLbNE+cj3wL9+VuQWKPfrL+92KF60hiHX
477XyJhsTU0hKEvzmq6YkKair0nE6YDMXDz0KrYV41/myycbGfbvwN/INeORbiR6T2ixGwkkHqSK
PU8M7riThpLJfzbbOrgURXQyEyiImGGfILx2aMsjChwKq3arGFY6sM4VWpbyFdyoz4gOHi0ELxbM
9jLrIVHWkoigu5636RDPBWvI4/Xe7Ef8Cq4eDTMmlWKwpny5Hjqg9tlJLxqNFzzQi138Wctog/Sn
HALCRQtdf+cDsA+gdePccOlRsM9h9Aj9EAJpwX0/j4AArB385zDfYpLsGgqmTsdITyZCkYI3iETz
M4l218lQ4YeaZIEhAtbJWXAIgsckLhNpTCI1d11dlU3fczlSEBCeeQIq4jNbj9dmkeLtCQdVoRry
Qyp18FPhgDp4m4tC2WmDwQe8bjew9SON06kYk0vEOZKJ0aEfDzhxX2AcOPI/glYjwgm46qVG1Pg2
y61gqV03t+0N4JNHWZlGeQ/o/z7Ass3ma0TZ9hvFGJ4PzXohdgLjeMOzzw6U897WK5eFxyjSaxdd
JOTiHZDBmDBTFUvC+LbDOo/CSCJmeYq4tJqwCViA5M4iy73yRNLyLyCc6OUcmKLF+hOHc8xqSVjN
kCkhsTg+AxiEjlwwniYZQFrq1dx19sIX8Odp7mO5nQfpLU/KUWlZTG94aKdamm+Ifchj4vJoCSpn
6XX06QjT9e8F5HuzsUpucF1ACPi9ivbGAtLwiDy+9l7+gOjSQ4SfhHMg94Il4WR8Y+Ux4pItxj7K
EnVCyF82GHsvIJW3bJVD2llER5JMHjAqLJldVpy6WmgOG20yn52K4gRTNUvz9fTRAgRIzsDYOoJG
tNRB1xRzAZS7f5btZ2bmp1FyWWs2DrnfqCLfHTX/T8WAz1+MPsu9pMg+OCtjDZCeOz2aef7Uie+/
gMwaMYh1wt3tJmBmAZ3sukfFAoAlIiVbohTLvKSUQY/rlHc+vrh4LcvNvhddP1Ltti1L4lYsgXYg
cqGUkOM5GCcjXIxy8TesY0yZUqLqp9j/4w5gNDnauZecAHNnfyBw1ETtk0iciVrJ3yVQgzSARzaI
7kgIyo0NCC5AF8yrZkD/Z7Q3rx/lE4bS3/ixxaFT1+bg3mdKVHNys3Iu1oWXVgQHbPJOYCOnk4UT
CmuFOxu2TAKJBIMlG1YyO3SZSGtpiuNQBjEY8qScQJOuNC4LAusOsOaEx/p6XS0Itgq7E+vgzouX
yU2lXiVvCgmQ34f1H/3ZIh/Deo56+hdWhXwpE3f3hbMiCMvvGm3SMUfjwbkKHWnFk12EC+eFZy2B
SmLz0e00z5LQhEsceCCUROeMdrM4UxP+HBIVpswJMKUcpD3jiZcKi02BRF+OopkCKqrFctXJR9IT
IBvkP+lDD/mjoOqarRk7Ak+aX+Nu6Vk2sXfhCpMZovLH14o4VQ71nQjmxCXf5vUzCf53YXTDRKkO
4MBiSW9a96OAUnqlzNQxNlF+zh7aosmN3YUBbN9n7fGbR8DriHv1HZfPckyanDyWRyCJ2Ik3kQla
pgHW1MHuuiAoXw4M2HZh5dOZRQ7pdpwNj4wJ6/yVwSULaFG6rfWI9rG2vbDss8kBjYhsV4/agYLm
Qap9DlORUA/4I6tUsmOfWrXeSMTJaSV8IEO+ylhVc+6bU0TF6vLjY/a2BZCNaCB/WUiuePNhs4Hx
lPL345k3W+q6pIEk+dxWQ72UorZ/d9nAedkgg6nln4K6fFv0P2sfFryzE4I8jNj9RJ8XuIVmFUFx
u8a17dTXUqHg5IMSsUrJZglZHubh3l5LXtiTdf+OP6MveCRimdNtvYnMkkZDOaE9kbDx74YVHZcV
JxDneGpeemUlKk7m0m8UfKCe7HVbyPUMSvv6S4Q91V3nICa7jq/ZhfOsIpKM6MXUfpiLwd9URF92
wFqRVF/cLlvTKWMON8MB+5w992GbFBJ3H6sHPTiuW7IOGlvh1fol3HX0EFNArxczwzrJollJ8Z5r
QSINa890PYEim9O1bpcrIBWsjfETMWz2scV3CtXuMmfVJqgXGgAFN5LqXIi7FJiVIiD9vciQaO+U
pWkNcQqWxNYPBxL6X1bJyGMSWXSkdvSpccpC7T2aJE6W7fkX4VI0+ujR363R/9m54/lRR+wivuQb
zu0BFjR/XOEmbaQZIwy1FF+027lbE7oxSQntugU9jEU9+xN+vuvVKdmECsHZQuWXpWcXcqa4IiCz
KZvs/MG1/cIcHrIJ7OIrZYDiSApFzkBIb8RDvDPRPlGyGHLA4zYThL4PEfpC/8CIdb7XKS19iQqB
vjUAkQn+6cDLf5PvEfQvEBMuDSyZ3wB3GGUerv0gEvLUIaneKDSRQmOyjGwz+aRHC0qSNQySnYHA
TANdDHj4YF2lD82B6YK+ck+AJd/+eDDKFlV0hh24+9rCBxseWGGf9om9mdM2pgAp/ush5TkTXW/x
6XMIQKi+6/4xe7NdpcERMoci6gSD0bZXHrwCKGFBI9uNJBb2IUtGV4F/BEVhIXfXAlufMRkk6qFA
BV1gNWp4EjLoua1jR2x2jrBOkJBt3Dafll51jrWUnpjKwapxMpfKni8EBgakuKSwZ5pUO8sy2Y5K
BB7qOugsejhvHj4zLdjxBbbDlUJkMV8Zur45F+2RGsSIddlqavLY0jQu5jd6db9xREP+qVGAoTm/
mKy2MG7o+9yBrzA94hWwAZ7c2Tf1KfidxcTAQF5vUK0oQso+tdd5HPcQNiQoqFE25mPbCNQERQjy
LBtI/JiM3GeeUwEqXaZXZwMiLZmSyUSeBu7JdyioWHNLRXagSKzybBtFQUGS1i7Dm0qtHcizl5o7
kkm20lmAzOkI1LI7HSQDjGFP5j/rhtVwQT9tQz9lOPbcTWhrX1aCP2PAtxGmCTsQlDKbkBtaOiOQ
0iPLMF6hoVnbiLnK+kFQyCMrDXkx2lhlG7XWixyiaq+FGpD73tVLVEJ27ihOgn9X5dbrCLx4T0gw
0Wjox+5ctfyzept/yGOzNFxXxQlWo1ImPnNpTzO4/ZFhlJtXxD18lIPifY3/PNmkZ9jnGejeEAxY
yzHUu5Dq/HSg/d1kWmlViu9DANwb8UUfaPVc1d0kqjnbeYN+4PynyA2Se6yX4STJA9rwN2M6pP0Z
2/hhbBzWGMzkjiv5KzHnoOBbisNiqWDyGE/P5u119X3h8uv/CIdxUcvAuoibXNf/Z1VIR34Mhi5J
mQ0t84WpyccrVopYYwfG9HNPhLEKF7Fp3PdeXCHR7Oyrku4I1Lu0j2JbBAu7hbFaLWsWJFCt7qVG
iEoFFKaIzlKP6D4SD/u6y1/cipJlLrtvIB4qyrew2zk/rGDXecHrxHSiKBGb4FTUJPZOUKUUbNmh
AiUtxBmgqD0jT8K2HNx0RkySrARZ1I9Y0dJHsaCobKoEoETaYzs/whAsZsfBbkOKWGo47EYEhPrn
KWoeaEzG2F6C83S3veMs7bOC8MU482QoZAL6yaRKxjDQ5Z5LLmlXNx43HYXgT1UH0N+73iztJDH0
9XbkUrMOWAvECQuJsQjQfnAuB6O9arWLcndbeMnsdQH6TcpxtRyKjlRXjCnzw4jjY2enmZApOWIR
PRxnwc0N8vpGUQpMvZI3Rzv7Gquhp/U3np6nEu/ZBL0ltj4gZ/RUkEx07p0YNG8FNnmkR4xaLAiO
plYapqsFrSWsZetl3cxYDb/6wQCnAl28ugh6DIQ2VPcEKp/oRF+wyAagOb9KWi7xFPhl2SbsoA9O
R03r7VL9sJBF97vBF2DJ0v5jeI3ueDSahQMydx5j2/Tzzuyllg0uAu81S7PDSNTzCb4zXxtoc4HV
8bBDMzfCRfAERBvNDwsq6MbZkKZ3wFAEuTijCatKJGtBvXVUaXLlYi1A1pIHq8d+0Quxdk7/SUBS
nmAN19MNuVED1oPuT8b0wZpcgBvE9laNE9H+CMzFJPMZOjQXzGTf0XnOQrZ4Lesnwk0/urJl9wLd
2RO1esjcbvEILXKCSGVB0Zu6HKYK4fixVrjWAhH8r/ggzGFV//blETfztOXXXwNYhvMTy6FrdZKY
dSQ1a87OgMG9pTOoPL2e915wZBkMRqvE3ZXW1fRoHT/Khxf0pYU/Bazjh6sOmh1v0IcO35gvRrpd
5TeXEKVTFh09FvXWpgiFLbOQfo7DEHKFpCIwKr/3oApDyh/miPVY0L9MmepRT9msuNwpHNjTIsyz
YNo9Ft/cgCSzZ4kB7N0+0tnT2BY2Gc1//tQmV+pA9q9kVpI+dtUhDsiYXelm0GbpXzSizvUeUqaD
o15kO4syQuhKmlCRTEmwKoP5e+k9o27AKp+DOQ4Dt/o1uJKM3vJFI/UJH7xNFE0PZ5B57cRQj5zL
0ORypAV7dLBbMsq8jwHkflLfnBO2/FbpGTqBITJe0Xt1KQIIxq2XdToxOUweDXMvGNB7a28WG7Cj
L2k1eRwV1Jk39M4KJMyT776/EzK8hzot/vikVNSL96SlMmaI5s4NSvgYY1dQsh9qXSR+u+Oqv085
k7/dYejhp3uZRW00N7ODXXUTuu+YbV+VDMoCp4UqsK89Y4uKERO9gqpATew9wOGN/sIniCl1xfkT
PC15JjbAsmMfhM34Y9pCbeh3/uFv+zh2gbA7kftTYnX8hr4BtfXFHMjvp0RlP3wTM0Qx8GGOeuDI
jUMlZUalHXw+AfDmFp2VRNYIvcFtunbop/LMgGu5+hKUuW4ljOAh/S+II45IjZxRy6gGKs/9ZNYl
vx5/R3tP9N0kUWSJqDuM5rOHLnGnpF5jmMfF8XT7JpXV6nmclzi4NDQzH/R0XIkBNkPu2S2LYXFv
iCxz0NaTnAk0sljXATn2KJDVkI2EehTTRWcYxe+MzJdCGv4LTkaMbMHqn2oMVd9r+BD12YD/oc97
93DBFfRnwowzYvfr0mqKqNcIOUCGtFD6Daj/DlUauEOAd6SXpunl8PvRbpwlqUDiXzn/trRZ01Iw
T4Ef/9O0wHguh6zmCVpA/ZVlYzyXg4JJE+lgspCAfCS+7XTH6VrT/UfXtf015mKSF8kE9PPZjIRi
IdbfwOfPOMtCudL50OfWnD+pnL0jSl1oVZmeO8q9LXB/5Ztnj+Y/rRfJd4U0dKNVLRM/QK8lnSAy
Nrb5PE6WEqZcJbmbyOh1qxhO+OVysybrYYKF8e2BlWuq/iFPgAkz3F6YpigyZSRaEIx+7W9MIgk8
CohPrqnf1XJ6MKWIqLs4xQ6vgLjx6BCAauZyIv5A1jihW4Ay6+/qxc0IcyFdxTLyjYIvw6GiytOg
y3yGReWAL8EPT99zaboi2L8D6v4dQbvL8wbCWTVgq/q+viJfSGTeXteQcdgFIwm2s1tNYoJ1bUtX
76pLftMpWFXIjc3CxjUoAH9XrygGpTUYOJvcltNJsRFZhng1VEK7+/aWqaBSy7kSUDZxniEGsLlf
qZylg5jWm9vnpmGAibzgVCDzD7ssnsBRe9cUSBh3oc+1lrfE827gWq6YVVZp/O02v5UCYldI+WdQ
fDyaqQ77p9yOxosB+MzF+9v6vThCz378w+9AYspTZL92+d0sT7GcGqEIJCW7L6HV1+sWnnF4gIfR
vbSA3z8i6JujYC7P/CTpQ0/0qC2U5ejZQ2XbbRAWWEMBmyzZSaadL8TceLrVrgLiyh/uJOp3kP2X
8ZIPYOf7mjcDxXmfLBriridmOg+F1uL/pJbwxRqymVX0QokVheBkvjKy3W3+DJVqUv8LxcjYD6C5
80JW90uxkkMORx1dlS54xlQvuBG8lbqf9wAvx7jf5cNOt6/eGF92yhMQP1MknCzYiMY0di7YhLtJ
il+H3dgcM1suRS9fbEodKyvV6FzwkWo6Q3Aehf/5NFYXClYcQA9HU8JCZpOsJ8A7ICi0as2aIRUA
UthUo5aeSG9MJkombQ15kYwz/NndNc1pYWunXhHvdBEXO8WXckmjZGKFjrnh4iu+UtI3kneG7upO
uPHJ1j21oubhBZ/mXcz3e4eYRRuiCEqZvZVUT2XLMfJNtECX2ltnP3mC2WP5N11z9Ipu6o/n/Oim
CmZJ/7I95g0DRKvgPh+Ar0zK2BIpccBYaPIfC4qWhRKuULODrAPL3xdutzICTR+JNx7cV7lg5izs
OveGVC6s2GSuJN9hWMewTB1L/ahhM0PheAWTai/gFwhKyliWkDHAUqiDzZoa2mz7DXJj+ErPS8hG
ieh/1/tOONDOD/Rv5s+5TAoprn5aXGGokgcZ0dkVgz8jHlDOZGtqL8GtCDwTzLXikNlL7O+WQbb3
cvlUNipy4G5iwotOVc/ImDL44rwQ7gY3esgwIZZdV5zZaxsQrejYw6tQNiPjiResIdWQX+2bpmJT
zR8pqOAz2iITd3UxheP85TB0I87T1ugOYT1SkqXchkYyflzZmrDycJHvWzz0pwtodRSqOotmZ7Bq
oruPxDSxN5EupejKLq6FvudVEfGYh4lJFCrdOKpiddccB9Kw4Kk6fS1V9LMBs1et3pGKtTpvM5Oz
UCDZ49z4T3a402J2IFSwmT2KLIMHEMYpXXTByvIu0mxcOZAki/aP8WSoiFxQbtpmJ0xntC2FFMzw
VA/WFnZ6uo2vRWErdxNKby+zTi8Iashk5LfStVkWh1sSKTI48b7HmXUiVyYL6ez2RjXperpmVDs8
EDSb5ZpHe1pU0rDOGqDN6aQpbNQ2Qt/LrAZtJTtIRgSwqkFNRE9lzpqQaFgpIqTDZ2COymBClMHU
4q22tdmLR8tTrH7Mbdo2AV0owrqWaWDFFD4tTsF5HcZ6CoVdRZEC4VtvmtW1lDRZirKU3XbGsR+v
x5m/WDkCjiFZdGEd1wQdmFdEl6D0sK9HUQGn0rKsiLMo1XL93NzwHHsdr3I+xaLksooBeB3qdhAC
P+dn8nyzNVqt9Q4wRfS07bGjtK3KYgzcM/uCah6MvD4xONWSvAH2ozmOeQlWPSp1kaHTfp7CBmOv
4Qi6BStJBlGS6FGWDH6YwGhO9H4cfxAha4fPqu6gmuR97G1zX2dmDAvQq7X5vZridT/S4uwkAI2x
FP1YRgZjijFcvwG7rIfWbKfwq++8LAgpFLHHMTjeK7DJDgp6eawJ48GIJ8+E+Qi5dcT1SuBFnbkl
X/7Tj4/6wXWmtGavIvlpqwoyVWNvNF4wU881zQWy7jWbmqyA2lewzcnC/1UqLmzpL3kyQ3Ugx6gh
anTpuyHY4lnV8Dvyrf0cspfe9cXTF76zF/S50+QiVQ/MUmA4lsEZAudinQe4sCa5G6/OSF70SVUM
PTQ7rSz/8ipDHJnO1TPcgOgQME+F9HU290d9KB6EKmgtHO+uPG2fDs5FW7rwIgyzsdGC0W3/Fg0t
rF+TS1gVcWw+FP5GloukNdlyI6l60qlYmOJ+FAW80eOdPDhC/RXqg11daBUsVJ6+44SGZQ7IPJHr
dn9W66X/ob1kX6Y089ZexgJuLFPfH/4YIbPqxg2E8CrbFpUX4lf53ZpiIUwfvpkQcN7a9zFs6SAq
IXELSagPkHch1tS4LL61SKGt+5/4fPsEKiQohaGe8hdJLpIpqI6O2naUDBr6PNIvtRUHCB4+YJyX
+i8h+t3SuQvddyK0+H1/r9ggfxiCDzPZulg/WR9jaeachtvZGyI8sOphmtxynRlfxXYZQmRXc//i
YLu4oebZAoDKdbk3gKzOTSAIuTnemsHBY2ixTUU60Rwd4snQlEtx8MGruTONC+LqF5I0CFWK9faR
sP6Lvug7FOWKtkuC7A9XV6CiCbsh0ugGIToWIdpDPctBvP66Mml8ik4PT/3K3pe/Ij3wV1VIyLmi
JYCB/75jGVyPP7LhGjUtVIleul7Txd1+u4aEnoglAB38hun0kGPUBHk6taC2qQuPHSS0nYBSX8Uu
LRXHsw7XpniBrZWYG3kHLlbQDeqB2dEqGozr+86EH5RZblsZsFxlYe0/8PJdT+CKMWeRu2x6ngDz
yvO284kmavSQPgiCs2cD7V4aBUy8JNtvAk9L1qGfl/PJH8ISlQqbAdpCC+ZcJdaBmQQDek4OPZSr
UNAkEt4CmNMythPMBwGmXjgxNLlU2oLj7TI+he8AHQAOjfQs6aDUvEG4xkx0/OYDQgI6EvnbMb2s
XzudAkNUi0h2aq1EdsestEvmL683RATYEhy9QMt/Lq79UfVFi9zsY53nK/+G7Eospo9zbcQWyiOD
MXSXfzguzhjGp/W+KxWjduCb00iWHD5cJjunb+w4dwURVVVcH5hppcQtKDnkqlE1+Tv4XkIafElM
n5GsJwKkkYgY4TvnyEMrHfk7N3iUEpB2T7FvNRtbjeJEF71RPmJ6OI0aw1lKxnDNFkOUPxPREIf3
Dc9WxuiJzFmDYC61ABGxvbPoZVBY/q+T9uKtwYR4iJDX/jC2BHq3QhREQ8KlKEQfBoIhfAE30yTR
jbpFmDCeftf1DiIcRs8NRcB+Bfriaetqhr6m0osiRWDo2l9KjcukR/BA7z69FvSg3ESe3pZOaz/w
l6CtIA8k/m3FcLlSMBA4GGO4d+5xH/lgh3CGXd3jAgZBDFCu3hFbWjssBdlZDIPIdn1RlXq5whoN
NXN+6BunVq+Ast13m9xX5h2/aq0jalVfyohXOJ6xLn3NGxoubHKv8WYd4Zz1rQUPGhgVB+vb0uCZ
UhFmuXzJoSo88vCwws58eXAPQp6cf1IlTS9gREnDlxH6ByPXATeyPXTUZI788MRjFs2BV9Us4ZwP
asr6X24RVf3SwuOZDBIuqR35UbbU01ZxtxSDATceHRQbEgp2W2AwBkN0bThKCjOg5RjN8v5JGcft
/jvswNbFtiIZp0TR9HfE9vy+SRycbUrKzTMbfmowVSQKwAjO7hWLkwM9aAC1HigU4NSS1JTWw0LW
6OrEM2kbq4kIWg86HuVkmlWrCRuFmtSqZECZm1ZdLTpBRpz9MZT1DFIITAxiwPKbQbThVG5eZ3M6
c/K2n5zv0GEfVUMKz8LwMv5PK0O3BUB+J2mTRK4mAwhdFOnXRQUbY1v5LCeLS0Ecu/AoY2cGmd7f
J/ywk5B9lsHUVNIsmUd2heTfxz4gaLCAZTP+tYl6M3/gkSPqjrHMxCTuLh7rLoB7GcPyjMjZARGa
ZEQHl5ckc9BPY/WxoFWoDNALtcJVKzBgZjWyBZ0n9cxuPTYfRo+S00EcsmETIDMTr8mcVbo8EiIL
oW+wpeEew8ZHP+dSuSWQl2wU4BY5aHXI1m6wQiGY/Przxbxhak35Hy2yzxelXDArqzINtEBef77M
qWYdvcCuGjkPgQKFnxAA0SzqdgAJx4sihwfO3q1yfyzeeTsf6KX6bIGC21FbMW7L82DpKi+xvvh+
eH3bYtOSo+w+gOTrECkoXygGDStyRwNDMrgIYJhYZhD9UXJV/HYy1S/1O/GM4CuPDBUz22XeI3Qc
SPuu/XS/xmKsQKY7nqnnLoXHSn20IEAHzZxATGN3QaSSQ5/Gl0DYYZWNVxWkCDlRy6yOPommXd3+
iaOOjO6Jzm7K9HkHyUuz8uobKCi+dmvaiYCz7I9k1Ah/UzlOUE5eHR0fsNEeVuJm5W/jgQ/kZ35u
DjhnO+iXs1sI/F7SM2NOwXOh3VJ+aNEZtZruCax945947BFCzJI+9qNBqz4mQGGsu2QpWJYej841
shKX/VI0nbOQY3dgkGigBzZWuMiq8beVWNaVnGzOzcSQAiqKJqhPtQqvGd+153JKgNBcAA6Az1eD
CQH0U9hyCObkpW8SSry+vpA2BoVgXparFyOJk0FAH6qm5wsMRaec8B3ydVCIU0o8KxEnfSKtta1p
RvikvpZxz8gUqAuM242eJ5LVfeytnb6i1lKiy9q9eFJoteox1umL7rfqAWoVbtrhz1VFY7AsVoEX
F8lX/YPV98IUlWOMiZf+Nvt+K3yolkmmlcYETol+si/NL8RnpP4iBaxyyVx91Gfa9UWqA9Dd0HH/
aFh3b2fhxEOi4y2rNVGgvvnqDgpaWbhKq332xeVKtAA0Js1UPSN2tLlfVh/1g0unE2dHWIcepky2
LrqW+2GYNZzxm9WWb8XaUC6iCQhcrI6fFWhV9NKtVolHpWRZfVKxmR2rV2lEUnxzrh4I3EmUJSWd
i8w2pBoHaVm8fj1LRaTnBx0X4M/RjtUpyoZiXbFja/POECpEAIgfs3xyXav043hvaOJZ1tr1FHFY
yEuF6aDHUcaBrbTb+ZJzyHWDe8eanWHhAO5ZcsaZ/+QXL8sCL5dKzmXamsKM33s1ra4YIoEsGHk5
aDuS23m5zN+CBdqaB+bl24BVuEPGPRSsWnuv6XqQgvUJsXx51bKlK32X3UisosZzOc82ugl9a7/s
k/rPA2iwv7CJO9VLDF2LSqvX9i489dBOHv/Oh8CVp/kPT+q3GDwLhzPTgJHHDpjSrxslAfPWi6Db
ucInK6BvdKmAPDxoIPbV/PCmIvYFMq1JUnYB3rvvpU6bk5/9MmCUTDZGurF2QuD6Jo/QHFbQfRax
CxgkMxe2Zjp7Y81HZL0Nn0Ajm/vpwxNCvDMr53ZlcbH/4Nn9tLoQj8lYTTLQ2poSIl+OGlyEe3cT
7sJkfZ317AUeeYg4up/2d0DH/WKV7NgeQxrO6Hx4JORmFF9UWew5OAftN8muABd6ttSKrbR0ANIA
QGGIuo6XFsGbNHag8LaEiuyzdzWuUF6uQgDmk3hQo8AZfw7JViokfuQ1n6tF4QjkZo4b6GEsXNlK
fpkJrSFE7OU+m2HdYELgt3sZskDhFhnBasZBf4bvwkWXsnqhsHHFoLXzrB1oWYA8pT7eiOJ3jjmK
exzgIx4rVmBsvfHNNioBr+ZW04W1yTZ+9kfv/RaRCBRWZAIBA9fW4gnHutR/d6n3b2K6fl35pLC9
0B2L4Lot3t46O3H+6JbaRzahQB7H58T0fQfYDQgvNhX40WuyNcOJ+oq2mtKsgVH1QDCNpRAixONA
t6W/wyzNNNK9hIqONkZMHkAVwnBPoIbkgtc9ngcPIbRfiXsX9qulDb/dbS68za1+c2QyrQcNfHYM
YSGmtt1U5dfG8qJIF+saJnd0YWzg1mnppLCcAPH5LcxrgvygU+LVYItZ9+qwpSTqFB+lm2ztnnBk
bbW9UK2cb37hSUf2Kc4K5ZWT8EkbUvZpujAZpftcOAUZg/29hXi71ViB5go5p19jiFbdr9mwaQWn
6uqvo28voo3EgO1SBH5T1nU7AjYX9lz5tHVOxc95sRQ/mRn56s1jMWOctscRs2024z/538yHu2Oo
C7bm0ZoD/Oj1peUyo4JW6ZSKOmYKGN4ppC4oshqOSEIe98MakNGQMu9d0ej6KIBufA8gbKU6WqON
XH0cMBxgKeRfKHHpspuGUGe47jk0pr3yN75FRvPq8WOmDrklGnOHl2lfF/ApK7MnePUj5Erwoqzj
GUxGgJYLlWyYrXOnFFofGb82M5X8YXYfInR+c8+N0M+1WF4LZNd8r4DyU/30I8QSZxMc0mK4F674
KmhRfoDPqzf9qxpFhl0qnuhxKjfLrMOLMZZWNfG7gS6VM5b0765gbctVV8ILtepfcXYo4dEFcpVC
xPWTl0I+WgzNMLMVAQ4tRiwo53WRDS7OsIhSCLdVzcIrg/dITGbQBLnVmq+/IDrCdEswKND9bPdZ
kwlaq1E07wbllCwc9oN47wPhNpGkUjhfK5NyfhykY5OZryn89iVqB2wGz0xQAkGQR7/6vdSqt7NJ
3T8I6g1o+K2GHKOokbL5+lUWjxepftzMr3FBEMrxAT3HEWCgq0x12kJGyKg3Wpc+8tzOjB1U1jt7
PzfROSbcB6uVwOoiAGXoSjXSP7U37oh8swvxJA8G/lveOpRS0FOpIg40VSW1saSIb8Bcmo+of/bN
DIS/jiMH5TG8WdRrieLb1CZMhpRKlI5l2xPbmCgSPYmrFa4KY+8H89Sb8F9cgplaOH5IRlqxoZZs
p0PPS74/K3XZ/HLuGD07S8WyuQI9r4tgaGg70clNxK6sAlltqWdCiy5zA0D3OYal4Ea7YPS8w69K
bEmaA9h8iZiAQ4bPkcTJj8LrDNrTCnxH2a+9KZ0GREkMF3i6zjbzhKPk7w2pj56slWpNRxQ4i+A8
+7Pl8inzwAK6aXqef7EwMG3NiWSlTmquWOhVJyKWDDqryZuq83rzccVy3fQbMvwd+b6pYCPhdYLw
vF6sekrI/ovNLy+RfPIkg2dHB896x9SLta66rLxiLeavdXSeqWvx09dXkoSHJkyQYHQnB6cd0CyE
3y2Z0uOs9e8B699ZABkNuuA2u57USjxzAOlDUiJA6v/cfGa3vAH2oMQ730wQ0i6cG12JC1qfEqaC
ZFTEchCERhxGl/HIR8huSDekXzeSEWk1MAbrW9jxfgidepwiHQP5UwK3+OdF9kmGxASErKp+RVkx
hEMO3a/aMTt4a0uLMOvQ2K3w/9M45E4LEGc0wIKGQaq0AIsY3Eh5ym+6VLkqZD8hdDrCIZPnAHx6
TYNYKQw5vuI5urV5nqtv6gTAtfqRp9Of8JGd4pZfxbSs4jQvIjKrt7s7tx7uv1+8xy26pZ4hCxb1
nje3zd8Bly3qQDHRpXYz2y44kZiPh5zvTrOfOG6PdL2RoGyBkLBKYUA0gvyIkgsteWXkxJI4NFLW
6EW/AghbJHV1bgfKcY8YirwGYYsPG/Fbfi+ZFXKjh0xKbNpeH4LrpvPvJ/eTGElqePH9OHW8NkGq
wGP4FilVLg5gj4n5SHh7iNDf73OO9V1om7bL6/rBWCSTQNEL83aKvvk39bWir61h80SAcDAJmFE+
qHIyzk3llubncDCeLv9zAEc+oGpN/UpVi91uZLdzLPzss9HuMK/uHL+tfPGqYUIn/hMnKO0POzEZ
L+JYkqCIT/4/qScqpMHfEjqzQyfCuw1KvilVHICOJsuMlEsLwS9P7fpioSQ+HHM16WbQFSS0dFBm
FN7Eu8Y2RGV52Ypxhm4aO+bo8oKsX4MznGF+QlgZmWnbZd9RFWJdfATq6iEkMGwBaQL8+A2rOMqP
YhCGw9HLyhFOiqdXeNkJ+LLTnq/30SoUjvHDf+3g7ehn9RXppsZW/3ghOroiU6/DVmzBjZibjPZo
dKWnSW6KL5EUGXpAkeHJp6U6dxrXM0JHpXaGLyCulE8iHz7+k4dd0gWWcFkUHc3JtgJ/RSF/mZ0i
HtumeO/uXE6cbYBDR+xhsgxcGfhhmcPSbj5SnqR9006z4xjrYTmPOsCNgJbfEyUy9KMZqjKFwZyp
BwtSy+e09ZcFzCObMNyFGwvHrd4aLB/Qia31vOvpHzGYJ2l/5dXq9OtuBEnya91xDfiAUI6RTi6k
8y1gjlN11xL42xzBD7Qpm/IGaCzCeSHgdbdbEJZheYDhZ7x1bLga0MbyOV8nXV9rFC0Kt5opqglG
4/OgoRumDO3+KMsn+SVeSyfpicO71YQrDzn5b9ro2PtV90S1nmBPoVEdtdvUoOZzcTeFK3JroHHN
bz8ilqd2noOGC6lYV2UDeaMJxtp7vDIoEziamU/ZTG5wneGiAQsCF5FvH5YTxZj8padxYiTNyD8C
BHtP56fAZ8lKCn1n3fH7mIju3dHq9j/H8d+Tx+rxWichCXTGBX1YY5BNEU+6MqR4fC5npqcGtmHf
bLTWVPnfBFZMG6oS3VqC8G5t3OaOjPnDNrfj9t/TF1UMydNQv/qwDZ5X+CKlWQGCackUg8RfoLkm
wLbah83FYzuX7tdCWCgtynw1PRoXWzso2rayLhTSR2h9RF07QpIcpE/cf3iPYmrHilOIGHRgHk6M
AwdJfrycUKNPP1+svJs2LPqTQXQFvYBgYxPMX4Habg4VRwsnmQjhDOUH0TtgBzPv1XbjU/1a2pgb
DywrNMY7t+bXS3BGP0mBE687P1W1mNzsDUuYAO87OVQhy0U2ZWSul8XzaJEem+arRgTtFoFpwGAx
Tnxy26oozvxTSLSrkNOoiIP/ctvjdZCLtFrkScUSC5TqunRmz4wLuSf3IdEVO2B+zluRLTmjg2N6
AciAvh9HFm1ftQQVLyb6BMpUITgiU13EHaxDT6n4PYhcMjmPrspmteGEKGKfbJvBLyYrt0TjsPuV
F+pmjioWo9ZlizZs9m/3khQH5/YZyZp3Yefr9/lnQ9XyEpSejfPw0XJ6WpVAwdTFjynSFQchP5N/
lV/0QL+i0rNoWXA9Y4+268ikU8SpOB3mVgCoWJnqMOWG6p+1kHSdPwVigwaY62TVa4aIwaExY/qP
68M17j1tkg2lK9mbqlI/JDFjZC4Cc2wV/5H9t9NFtF9nMtc6rmdt4khGb4CBK1kFMN+kvxgwOFKw
TfxpvJCTNWey7orqIlfspnrOKUQrTQUE3KVWR4ywMtdqxFUIT2AWMlZN1QO/IpBq7jWD4oTR61n6
QNz5g7aESVeSreF168Ra/X6QTSLk9xjLqrZLk0N2gpiugIn9WoVroDuxspkQSW3CsO6Pny4SqCmT
1Jm7f9CD2yobXXtuImXrgaaGhLwL5gcwoGboX3OTEBCzJ/ltBm6ByMi4VomIPHtVXBDobV9mBMdo
GJUevpfFCd7NI3WDWzluRS6MEvu4pdSus1X2piX+8fHbTa5J2vK1db/dkAHGrn/I399sd8QKNbRZ
ls7hFVLcLIWRa/H0dIkn5r2jKy72YBXHAOrJLQ2KE4mpQd2P55FQat7MWEJQENCsjN4d1/se5QYo
QHWUM1Q4wSGxAeQlUo2ROkbt0qXPhyoZzby9lNzhjx6xh8itHs+OcxnJgd0XH7FvO5kImYWCeeYe
S4H8AZ2ED8DHGh8azxqUp0wq30opvSQWeqi/fZ8wClOzjPRyTBxPgu+JOQfvsVKGFOaxuozvV1Sg
3QHm8Xn6dXaWAsSDO3VRGkva/JeL1w18EOR4kc+WT/47ieg+kE81e2MySAjB7Uhq6I3aQ7Yqi8xQ
bYroidD2oYHXBLMLEjCzx33SuU46wmgY4VEgvhaTYFLHgaUpEzUmerB9isZG+X7U+HagJbkXeoEQ
QD92YTWzgn7oz9rjS5GBeodMf5rJa3CPlirXtlDDDatVTFgNyJ08ntHP/k8ThQTmfnWDGGQO1YUQ
vrNQE5eW3MRVQF3NbdzYE2Qv2E1bBQr2DXA2K4ucwUZ1VJEXcLHiJGw0ug7JfNS+KCnGMNA9N9Z1
wxzXd/junHH2JbV/aILRysmERWzTR/GrrOcNPIG0ZdcuLB3+B15NJO26usDdRel2sQVpUCyX8Be/
+V3Rgdi5l+V0eeoKx8Dlk2laSLlh9oZe/NG57dztWlMur/FUVUW5D46oNh+jP8TZxBYo/HOwgwcg
TS1ypIy9TbbG65n6fviKDAOwM+QluamVtjekFsTvtuJQgsN31dBFgu+9wRmzA3jcqtV8tXauyITk
D9cF2lZopvvIDOina4eg5E0m6xNTotnHvPXhjk7hUXSLGoGGYAvlmNoLJlhIcukeDjWhcxK56TdT
Wv2AerloT6hemARaMGdKVYSSnjC5q3Tju7eauP1B0dCnsyGSEYWAAtvL73vmk+kaS6DiaOZ7Xwh+
e9XnWL3PE6OWsDO/NF+EdRegYF15lDK5D0iEDBD3ThEG4SBxBje/n6cDczt3tYyNDXwwKqhmxFp+
N0Dwk7REPeBa2aT6aLT9zFxPUxP9pXMYhh1kUgGSNp3CgjYxWPV/zAgbyabKW/P39eY28XOxiC1U
4pnSrScu0b4G9NzklulA+q+L/sKsoZLeDo1mHziXfNyEAv5ZxzatO77mRNLMgj4Pp+UNeMQzV5kq
DYPDK1DN31b6447ZhD33vgD4Ypw+SGBa8FDVRHDBs7juc3Ex6MghNra91+g70I5x9mApAIghJweI
CGYQiQt5LqNXNwY4G1MWfksbErwwfQX+IjCp/8dkauOf33ncJqH3bhk0FArweGzpFDw2DGCJgkao
cxhBibvdwWncmmc73e91ZZoPuaMMbtsokufOzqGbHKsN8ynJYT+1ona4CFhip94K4DLHflAExP3P
cHhx2pMgjWhxgEyatZ/TLN7bLWxQ+IKwbzOTJiyUpCAPyIprXuZCqjBnO7ztPUdt7Lf0v8/AVSEB
IDILWlYk0jre3sPARdSk1keJuhtqahO2Rsc3kbuVNa4BwrYxDUt4Xdy9xZbaCaxEyahYHmefEteR
j7vmJ78UxBkAzbjh8KS40+fwxMqA4Eab9CpUAcsSE6gDOmljL23J+vEb3WT2fAXKaLULtzLOAcco
vn/CztAxFWuVPlYen95VXMijbkD29nz2sSkxXNKl+a/UGHuF5zHbIpVM8zgxK1VLjwJdn8zGbRws
yqFtU4vzSP4pS2CCXdfnwIROu6Vv8RJ/hNrSSJrBmNiVbgs7PWES3yroDa7iX2zmA/+f0MUctu6A
KHVxdRxY9tZv6ha1RZQ7obn+Y8N0CiG69dQfr2mnxwLAznRSyimGTwp+hTfd7YqxfHfGiThGK8B0
72sRQoGmcaeFy7LrUpvCGr20dfvJJYfXPxtkXJffh8rpOv4y9YJfbO0UyXIuJ9FZZtsJH7wToqLb
xXhnApr9vpqQNpgG/OAFcRuI+TRXzkf87rrwqz3QQlCF2zxRq0472IA4Zwut78ZAKNfK71c5AF4I
CezEDSITFaNDKwEm4k/ktqVShi50lEHldm51fCx/nK7NfhMXeWAZ6hFxioyEN9VgkMF+PA+HMyWT
mmHNlOS6mBkbgv5AZ8trOUTAuKDo2c6VtkLrL/cslPOtAO9k/NTXmOvUT07yDTJEp2i8nxOw4Kd9
D+YqcUR1+7HDu3YL0eMYqKXo8JYkjwHw3uL3/OmDTOTANsekuZc7jJLGLNpunr+Rf3xMlTlQGi7N
VXfOImGvvN15dU/oX7lqHLtDSPQSTM0oAvT2ku/CibaJ+fCGK5o5Pu3ioz0h5DNOj+lIeUWUiWM0
0+NYWBg+G6FYhvd6dcmyzW7jXMVRtb+p9iONo/bmv8j7LHKW2XxJJeL15SEY00GPPmYObnu3Ybbs
kaJ3EIhfqTzen7Q2TNh7U2cYpSKT+QW4sK+b3jiBXb/qZeRWd6EhAC9CtIfnwHi9gcS4oQ96uiOR
PkmJmsox1dUr2azvC08A//ZbhKxlQvi+cpkOqQmN1zPp3UmhQBTKNbto3d9oy2WnXGFfSz+LqXkV
H74v7xyXG/fKQnoFQUwE4DQhr1Lq8hqYJ5DPCofbSdhYlBTr2Hebcsw+5lho/o1QOK95WXWf2XVW
PB7O5uCGfqqVnQkUTXGFIdZt2QkAFM1tpQwORm05SBFdcXyTeMbhPCn3JpQhJ9CTLtOexF5GEFFf
1ApKufPM728qnBFFURs4DF+E3nYMJxyJe6KnDdJ+IHvzTN6JUA0nZJ8IJW4+WuSDrMMrqDJuv9d9
hNcHFQogsdbLL11BcsD4mAK3v9jt5si+k3KdwOH0tzn3wrvb91R8dMKHY7Ly/AfHh5css/pjyi3E
3Lt2gGshYNyf5FyeIgB/ClewqtDeUX6ByyYZt+XIRU2yS5Qt9ucxGlTGQnegJlieBbIvy8gjc85m
FSLhSLa3ApA/pbSlt7JPr5KB9vOgsdJzt0QRBarq9/n8IHRLNf3vnmEr8cfQQQ+1IeEmnX92jfzx
nxFC9tJzwuYvs5rtgn61ZtGYsHoKBdUlKnKAjXVROQxfDCUqigxW/Kvn5IVbwrTYtr1m3A0zaHbZ
myQthIiybWGpwvWhde8IzG1B6172AiVrEn+68FvriWH6hqDtKsGUVmCXXTXwDwAXTidM/RNpfVLr
3lyIonzXWQTw6WSJtZROGqMwQSomJxDGxAnit/Y/7DDAiFK7ddh2I3RSzy98zFpN/rfNrOrh+LTk
q36VeqvHdHyFp+ja3R0oJQwyxgGdegCeBvewxQF5IGFBFdvXNQiDFVUA9r+WhwJt3ivVRrp5h54x
ynbdRDBwKmi3Yg/J5thrGOSkKlW/QJBYfURM+Jcyh8xj6Go9tUcBYGLs15HAe/rLIKmPvx1pX4ME
B/yVHpVTPNW1DrhikqnYmNGQ5LOQVKzjBDOsowwOB4iS+IsyhwCHIZ4LcLKEzJxgjYtTjE5zNTWM
LVOHAEAUmBXVXDB5QWR9qJFfjSSNOkCTBFla3LOaNx0zqq9DkMEQFKgxe36jDDBliqfClHvgqxS1
Ble0px0wUQYKMs+sZEC/sX7Hyu1oWaUGMMpzk/nC3qCvIxPBpiQ7L55fn8uVsXxcwBYF4qCJPInh
Gnen53LuxsWfFnZCJEfM3TR+ERr6Jjap+gKx1My0Qu6bUycocNU7yGYUSuXdIUJnBFkS+UhBOcIq
3QuSUTcFjoF6A3H3lve69kzfdtvODflR1DUSmUlvHuFFn3pEI15j+8srMT53GeZovQA8lJecLwGy
W3QtWmzgeQyyZXeo+17WS09IGn1uOMn4+2jufr2qv20FyYAJ5ZaGbGosMxukDjAfr9TbMdmEcXoF
uhNQEOO3FKdG90uzDl5xTXkLdCFo+RW7xkUDSg5eKKpMxDgjrNe+OPrd3bBhJ+xjlcjdgu2U3+x5
AMqE+bv59HG0gAMB9bPn3IbKvfhg/KM1+lXenwE9R8mM7raXNoTcZ1lr6fwNw1TRfiJUhZAVE+fy
nFnhdaXtoHVjufiCGkRT1ZxJuQpl7d8KRLVix+oIrbRqBCEJe3IXqgJaJjbb8fdyvua/Kp+5tdVO
N5Vs1fALjcR/04S+xjvHeEl1qOXL928m54iC/GNeBDE/fZYaROulPOJIME7+l+v+o2eJgGlhCdgB
b0jh83K7WVA3CB2AH0koQJ/3kxqYG1NeIFkT4+rLIueYScmLPeod0kBBuHYMDxMfvY++5wwBnnpj
vJ0X67sGfbTJfRI9sBvsutqhjL6RNUwoVHCP0C/3bBdST/l2dNfVo6QtH54OMVJyNKtc22Amwl91
PeyNm+1onSjtPnhu9rN2o8pnZFEsiUlx8RDLJfonC8I8Tvl2wIj1x+PsBeASX5Ll7taM4RKqbkMg
v15nmV6JtwHazQwmpLVOSswubYtZPjP56Vb6Hh2ZLaIe58dgrOC9g4+XPoUNX+P7LRsEZNpvIiUM
e5tDFa7NlpM0TuyKHH6n7EsR4xVeZfUsD4lmhqC6I5DJVgOmZ/TBqv5jXsGb1em4rT7Mu7SFVpKr
Jlhban/u0F6v4qip/2iX6VRgkAdr/9Sz/JGEJYrsKbEFx5iAdWuMQnw1bOuyCgHn88P0XmTHkU91
afk/94d07XpPhaVvqi6K9q/arjoLgNwHkERwnZwDr6+1iZrfcnXX8tKSQzLBH7jT10CyvU1K2Gwj
7KLg+CykmVH+F8rzC8hwY/zYejSx8oRuJf6F3rjGZvgJYvkDQAExdiuD25x5ftBzbnrAEBucgf0I
1gw0yKZLDLPHoB4BJlZR6fQ7M28FSqcwFJFK9MPQPmUUDadNaQEveXdCjsEX83lzAdpGSlSN9kY0
F4yKr6x5fnTTOFVpq43k5GXF1ujYH/1Lro9X5dvNz1INBe0Z1pxrUSFPUUY3WinkfwMU4D9lCFH8
WecQy3LBpGCY5IN+ARzSpKx4j0cSiIvpbnh8cOCSn2MzMgvZQsjIdP4wvgNQ+CUBmKF8ZNjLJqpf
47wRcM2oelrxo6A7l8i0eTjMfqlmwdYM7YrOUFre8cmpvm7VWjAA/oyXTYKASkEnx18BQLwKNIZT
bQ1ukY6Xz8Y6QQOGpzy+1zGr7p7XSskIUvfWxIJU7nCwojpgSO0uZmmkp6Qben1LKDZITHZUYotV
46f8jROHgGZaD9UYcLBlCufzjLggmZRwqMPJKQlM+vPWmDGrUjRal/k/O6paKsjJ9SAMSGJPE5j+
tRrzlDffA46eNSjEEdJOruVQyMsIylEeGNCVBSZJtzEkGilg1dA2scJUgMylDJ66FNNj2r+fqGEh
NxUGfGDkozjUUSXn0JyICcAytK+gHx2bmkeMsDdCXgedcWeLoixawsKHrf6cLN2gQdKHX6NWsIH8
AAdBA5IQM9DdcJ+kNvHJIchNUUy4yosEvFu50GkyRzkI0YWuWT20wsv8xeZd5EnS+izpj4ZCd/dF
ctQAgou64uHkx2InrC4g+YrAkbjtn+FOQNdb7EQAJBphKyf+UwL4+3+PyINcdzTC0wepVTw+wbws
rR6ddGB9rrZ4fiARRlCC9ESNob/w75wHkIwzYxTl7LZXivKIcaAKhLBrSaC//0frWXn16qsJdKRC
Z2BFVjlKBUEALboWOKEH8+Guc2VAdcFjjGE9to1G+N2zhfDo/F4w5big0ADfsfp8A7RBlx6VeO2v
SAgRGZSo+jIY8YsAa0P9p9eZAkB5PjZXK/fC63PX/UBalOmj/9rz4ROLqaTxOXVr/DEqyJAexBR6
t3j+bJzrdllUrJm4goRoEJxDUyGUQAgofdE7BuNrfzJ86CXur90b7Fer9mexETZFL8a0kcvWVmIC
rw28pM+8Y51qReB96fmNOypzg8N0VKrQ05H5kWvwAhIJkN0EzbdwtMYnF1DWcZmfqXE2gESJvSat
oLfA5yeb8wNZ7ss6eFA5M5Efmu9OIroK3rOc5kSZ/YHdlxXCh12xhHOytzsILxXOjiDdj6s/XwUT
OGwNOiZAYfj3k4LXgTOQau2LjRKlLif+RfDcx8UpBIUfNZdvsvjHSw31GeuNb/nHb6czb+e9KyLm
yIBtTg1+i8TanLE16BUmTL2Mydd3Ytql2xTQsJwM5XBiSKPGcLyeORpLc8UkC5Y36vDwx+zn7He7
26w/ZVG2qEPXPAd8T7ZTb8fRVs3AQefwMxSHRgIyD3CjHXldKG4asrytROy+SfWgWIvOVJnen3kN
3dcICyVU9jGIhjd7EgKsDPH1OrW91uuyYEb0JnOdhdGTgeIxFRPM2tBrY2LZTGYIp+j12mGF8Jtr
owoIrNhduVYr2D+8ntF1N+dJieDf8mlqLM68bxS+hLc1kiNmPd7qCtRCK0eeDbQQUKF6Av6OlVfj
bhZhDfYvVzzOe911hIQUrKtiXqTPauYVR9SFo6BmwJ78GVXoBrqxYp1AKSc+jaWorb3ciOYn2MN7
ZRrREklU5QygVgcqRKNwCAioeFq1uylkVw0fNRejUlgCbFN+0lomq8NCxW0QrHWOph2sRw8ERR3Z
w4oxFJLYMokdNBsiPzn9Iv8KFsBd+ew0uBSpK3MxqCb38CJ2pGx7P0slvrdB3BpPhWKYxJOHKZsq
cte+hjzkxg7Td8+ruBtMJ7R/gqOnYy32x9j3GEM+Jbr3mwsNvpLVwy97uqKwrOB8XcAznqwM5Tzd
VnMfg+LCFwinfPQFpEGsyB1gfJLQ6CpAFc3ORUZuO6u6Fq2sNnvEwEVnTH+binWhJU0xksIUD8rq
eh+AzOIxHYkzmTN5vhFtcT2IwtgfTpWuDjHgTx4UbQ1LIZSRr8dXXh5uN5L+Si4rb0zjzPD1ocJz
8kvfn4iMzPvbj9ZPJvQsn7hU8OkHuBYuDIr9xshmXumcFL4tdeLXYUEvMImPltD1OUn+2ubhDiXW
QW4YIAo6HngaO9krzI5z7dDRnmi4vtgBfHarBz/8gpE/ZcxR6fgz+eVnVi1RaXjzszlaHA8tNoZz
CMfRq5sDQ0sp51AgqkJpLmat2w+0m8fIIi4TykTyE5j0TaJ+5xb8EfpGsjOcgNATICOt01u/NgBb
c4oBmS27Ahm/VfE5WjK6UD2wqu7Kdat1xWFzSKQHOtexdcOXL2wuYHcB1pRUmzOa/NXh8DAPQSzF
3Lyqwzdf7k9Y96W/b4U76QUayA+Z3o7a4k3N9wpu0TkEJjqChW0cQX0JW/U8pQ1BjfTc3ifZ67Xk
tZeWPVB91E7bUUxzzz3Ocvz5EsjGLbwPXP4ojEY3lwEH/+MBq05X8hjuaN2DBsbpdoWKvzauYfh+
7Wl/g/U8IDFwjbuzhGdglXJYf9fIpSkpRiet7fkW00lKOzknYRmzQY2VwerDJVOewjsBiyoIoksa
nkBM5BH58qwQNg1YeAE10CNzfVCYP2pow0Sz+FCJMn4F2s+DFD2C8ePeGZ+om00j22UiUcdfkbZ7
/OuonizImKZMktKeZ/CVixG7ke8cOhohXdxy1chUrGxLfpVI1xVyyrZVp6BKAM/V8b+e6zGuJaQu
1ep3PlXJAbGzPOfCpkq/VwXXZBgXFQLsk24a3wk8qIzHPxEOTTbOjkrF+FCNOvCi4XoMNbr8+Obm
9c0zyYCZxzT3XGkGXTsVjrqguLK3C/emdvXVSK4CLL2ZMwX5odsY7raNhv1hm/Gshw2CeO7MA4d1
dSuxCmfteu2XSmDKKdL2oQuJg9zvhvyfO5OpR7p+ZiOil0zn27aLySkDDo2EGZJRsqVeTMqxybQK
ztJNAjO731//xFg+nc7UvA7DAIB8CnONv2ImmdWFJpon/79yqbQc8jRfdyaEqVWMNZN+XvoFbzgI
8x6v3zuktLGeGQ+Y/UXNJxalrS8TU7bJUN7subCQJpt5KFAj9mQg0gZXg0MZqjFD2ZKOSMqtiYcO
4jJhj04iQQOCcATuB+058dCV4COZIZH6hBeL6eFWlBCw/L/+L98fnqqaEkjjRUBlWDFhbe+5H735
tI4yRYt+FdJUNZL2BotoaV5LYbaaKYg34DWMV9CcbqGTABu4robepO5z79NYNKq907pqG66iKRcX
5GpPT5TcISozaMBMj9nCOhcHDKOaA32ySKva0dDE3/vseDtMch/6Dwk4itjGDTjX3Q1BURLCqrDc
a+9Cf0VdTQ9fpzf27NSE2JOkGvmSabopbvKGDoIw6EWM1NNibZ0zelViJ1OsPiHqGJArlgJP+ud+
8DP16pIw2CQUXXNMYntxmocaBIIwcXuaLpwtZM538J6NwvhmfhvE68Z6p280iUsj7L++pHqFRJi+
f8Y0HLwzn9VezEdSWGrdou93NvC7gZgXxG2DDi5wNurXYdyUHFUdECfcITf+7ASdU2HVTNlafL+M
p6Q3+Gi5+auLv+zA/zLqkWXdWoyGB+xs1rVxLWnTNrc7LHNdovK1asiGPUd8zCZ7TsJ17rAX52lv
sAZPjih7m1CqwplFBx9P9MJRokoLB+iqcQoaTBoItnWwd96GtN/xiOprLYekuqgwOnIXYgk48fqF
qBM49nykcHCWlaTpsIpZfvfl5dBQ/QhzBBdwH60HyMpi79z+PBqEruhteCebYWpUNKoKG3lNhrbX
GM7ffFsrA0MRFHr1SL049zP6DNxEmg5ZZKoDffNx8nmCvfWLZ+i7PB2d8CvvSGhir64lVw+mVgw3
Eq3F3cnB979mHgy1TO8nwPKDHCmoyj5SVLIvXB+z3Z61HohLvcaBopaqA4drz9ObHw0vL8L3HymR
s3XCPGaGgmVwnRBnRTNWxESgAhYNmqNOeczSPEhCSKkh9ZaVwxXGJ7rYxS/Sr0MD/YVTk/Q9m7In
VOeDh0qwqoP5e74fJg+BSX8oGxMFYiTVNzCPYYdzqpFNBtvlG3wqL4Kica+gTHbvO0WBA6aMajnY
yXdytyqGklybZai790abSEzdaphsvvE7kEMS8+y+efr095bXZNwZGOGfv2YBggDPtN77CqWVb5Zd
8EZHrtWoBIVt+0mdGNPo7+iR3Ohs+qnlXosxBvOVT6ucvz9w1YCCKIJUoN8tHmmXCh/X+ZSkt7yr
4XfmwgYDbj5c8Q9y74ud8AUvOy+uDXyAno92kXLFl+B5TvXjWL9pMQ8fhULewgkgTfyhp2xha5Kw
u4Pre1LkPEIgzeI887s+aFyzxkyzVwmjyDLJK0NvZ7kaNBXsKcL5y21WEFPz8AFZhjsbKzV+0QO+
/vbVwwMqsabrxDnBZDuj/GLAaXyo9j+Us8mAuG5/LziMLoJI4US1PE+t+4p3AuBxIEfBvy4zdwqG
pQgvyb3XxMKs9VuUeCPsoP/pG6YpGKGdcHzhR+Snmop0RNI6ZXmzs3IbZUvx8YFmVnFgcj1g71oV
rKuyfN0/llc25HBYaCzcyiDELfQdgv/Be/+8o7Gz6PwPYcwZC1h624Ea4iluKbI/kFy0y4uopKto
n8PgWMxWgu9YK093y2TTVQbhlky32M18KysX8xiClx7e1nfuPw1QpPX5Qn+XO/lwtqKSAn2wn3Bn
LMK1afAHDhXwlLp4vfhKFV0ms43B7thxvhBT9RhfUAgp9zt+aVbz+8EyTAiDH3Vyhnvq3ZDXjKq/
MR4nR725ucnI1Tb4uoRrI6cK0muVMWhPhEHUoDSJU2c/0d51Y2ez9w+/fGZ6Pf9kmomtMFuIn4Zl
VfuqwFkm68UhsH2kNoZIQhMDml7q+0Nz9YBUVsTI4hKCl+O7NBXIDNtZ3faHuCl8HODmljMnuHnx
c364eYNbA4UJptY7v/rYvb7/v+KMU3vnsx8jRPeZuhNzsEOX5bnJligCVNjkWpnBQk2SEBFowmtE
nKwvRGpGd940M2G+LiQe2tXFLxFHai1jFtPIWyodFag+tCVlPG0DUmb5IVpCXC37IheXG78Jzg6d
Ht7RbU+jkCfJaRKSXLdlRg8RrStFL/jtSKbWz1DLO1mahy1LjRgI69qNWzj/4W1XSUM7Ehya3Oel
lR7u3a+q6YMQB3ORiMyyrBKl+TW5dRFKnx/nBxQ0nCDD9B57YfgUX4SJrjbIzMGUfoNPDByowN2b
fdJBY3mWFuZP16WJA0AWwhxvYjtN2PmzzFhJ2CNvtxQG/z5yL6G4sLrfGV4vxhy8bunMjey0zmMg
APfkkb7k36eRJrySb99mAH1vTLjifob0Nm8Ocshp0IsT2A3+6NCW0IA6p0hmuXIOb3Mte1JhHeRA
/8KSDDpGAc4gHogskNx+Y7GBaucZOmMx7ygHWT7j59GV+VPkbPzbkHRzZDnvgoi6JFLBZA1FYA57
sp4qMrtQM0ijdeP6R7dYi2OdIwCHHHPavy2pXhYAqEv7JLPQxuAAyOc6KYcXPsTl0p5FeJwNr2EY
+GpDWHo+bz6wFd+dSqUkZQ+oG2iyahbsqBd7DQQAKi1zdZvgI8PAqc9cubZeCjDW8AnPF2bX2fj0
rr4vcFGXQW8iUF7Q2XpgvlvMuZhvuKFGS03hTI3tOlwAZkLlNQUFCmnhn35mzYXeCsh5ty9Bsqyx
nuHrEmKYuaNbBkQhhRYeKcY1VNLWd7FF9JlflQaT5y1yamb6VCC6oXDFZPdeC85rj1JC+Jqmm9KJ
r42+XGDtV5icvvPvkDfLZ+URBip6ozeFbAwM0t9txOqEfLSV7V3X3YKfdM0owwpv+nSoCL9B9yxd
WAdyAzHL3sw+9oT5nXjdkXoFgnHciwy6lot27UG78enC+B/QVkzEmRMFSpuXfn5xWH3MZVVZYjyx
xcEUW/ISIvJfmksWw6Yd8NnU9dnA7QQMeMYo0dGeRAX6a30bUFWXHsHNRiIhNoiHb/XNh1Q4w0RL
OuDgh252uly10OchQvUBInDdnew1bseL9dXR0OFnXA5waj/j1xBR/tQscMiHDriYuVnsSQ7y3RB6
ScQNf/dxJvyfsOwwDrHg+q+s3Jtt8UpWfHt0pacYXe7SHHo9lb499WLrIr13R1jIUkTI1U+CAwAf
41OM4bgLJ2b5q4txd2AkPegV1aDUO64cozXWbKySZcODaQVabAnusQ0o/Y3p0Ml3xx07U2iC9lBh
gAxfHrsaFsgTBRhjHVj2izx36p2qnnioJXNV95WNnJSwMTGwVsVwGFvwik3MAINaHFPamiJsyRyP
zGG/8zS1aXJjhcAjOChqsYxw3f6IngerPyyNCT0RR/dstCVl04lbY3qBulJ1talRZO8rLeasTa8M
9FP5HlYy9mu0iHA36qYWFTWKoFaBJKLnamFrEZOjP5864RbD9KTy6TPE0d+Qc+gqHzKKRYUC3gzU
ok66LgkgIfBugkJVzmsDpEx2HbcrIYnIOfVykrDVYn+thAvUGI/iNNJFN2AqXw8QQdJqz+UZ0DlU
X8J5tY9cxo5qyyS/bEaVk045Ra85sWEF4AB2wWpEyAtEfCf07MZXmRyg233ke9NVyPPdPuJDejD0
nXsv4OA/qzV0TOeFe+INv+Kisx4RuELI2guDa3rhTUlENpz7xdpGZn8mg6bAeeh+Rp0ovvORcNok
l+U0FEcIpFwufWudSwdSNiJuYbfKj2s13ZdNncKnmR2TgUIG4vuqh6t3GvMCxzARvMog2PnUkVa1
djEl8TB+1++YBf8XHPDupkMr3eNMBp5jE3KP6yGyoNQK71XCZbpPrJZKdIikGFPnP6nJRly2D7HG
RdLCykojrMqF9LGkNJbq+mZjfHjv+2+PwxinPO3tIsQTAfCsghHARPCNm9e4alLzPZJfAY3FjRIU
uwY3kFYoOy6uGyRaHzRotwvgzNNiUyaphT4cgrjRKWd+fyVJFop/4SJ7h+I08NIVqs+qah6iuamk
CJNDYFSZu60Sd2DKG7Q1qJyw2lEvUY0k7Uq/ru/vC1zBDfmsrn1JDp4D0AB9QSLYtxAFkxSrBPd6
ZY0M4jkVD49Jp8lfZnnKQbMe5YkEg4iMhyXOW0iyn5XK7m1Sis5NfnwxQ2Nt/RMzTvtTqbyL8V8X
1YOkVSbUlOlb5jOezH2XP5TtIc6XjmvlzpBQTU5o/n9QH3WGiNjCKO41xU8BEqKzpeA7vcIcV+QW
eK6fTPennphTd/HiMxN9t51oxjNnVP/dFinQDPK1Bl3bjNoXZIq5BtGRMgzpS8PLntpKMuT/M9kf
geh5xZE5RwL1ZJ2qOzF3UM8EcpaYnSoaT1+1ocr5cu2W8Ay8ny4x5Wqf0APIV5xk+Qu1Lb4OWrtD
0iMUqfZjV7SGlKpkeVuULl5s/Td9fRZVWRcXPuurwuNATPpZr1XYvRIKA1ffIsGQemE5AP6s7bXx
48caGZId/chmiBH9OgR0O63GB7Xh89p2IJF4hTdA1JeKpm7WxxcavAOqqznR7mUlLUw010DiDmZa
xU1853PQAmmY+iQjuBPHj2y36/KBaYVYfFr0PkEjE22p3YQ6dvszcmeInpf0kiXDsbWMpyAl3NLw
gUx7wKLqlXBu+YvETrUe90gP+xgRVBhcGNweF9Oe/o4oRX94Xqlu/kVey0dkr6ZY8Xb/7u5o7aAc
Ft7wUFatBx9EHbRp749Vsj9PcilRGm/ULR6IjEohBQq5I+vrarAaoHmEdvoK2akMF55yZvUiWN6U
NiAjHfCyiriz167bPOqYVpx41CTr2Wvx7ND8zsM2RhqE+ZxQuq9iffrClsxIwWqLAeb7nC05Lt0b
TvgufpMkcsbzxOHvkNrVkRY2eJIL6WuM8n+2KRGTGFcKJOvxrGsHdnAV0yWq4SMfvEhxSj2Py3MF
QlzYd0B0KQ+Q/pvdjdJ1XvJkoEegk9XK3+6CxbeyZW3f2jcq5MNLihTLu47VwuTg6YoojotfMn/3
nVEJhv9qVlJnis8/n3UU78RKoWS7yd+bBm771kntcEjNWzVZVKP7oGAdjg+jpKmIUdy94QsBcYwz
1rjVmgEnleH0ds/aiHDyz6NI4AhtYXZynj8wwT/gHVNRHpTXmYdglUQDGIJvo4ii45KRoigDkDYK
kvx1RumwwxgESoQXnGTb7DLQxmm6yKl1K871MXvglfAvEXvx0qOSvJT5VEPYgdwJMjbrULATyCjZ
VLES3oGRH7tV8A4rg2G3GzJq5u3U50+pKz2Zkb3ynpGKZP39rgChhuzMF67HE1a+MczYvO0uXArP
JQ/T4eXi2fCAo0ogiTs0VDtkdz1FRwpzIp053UMXByAP8cOYtPBgNzM5Aq5TeAHgE4Q+b50toEAK
+xy7r43LKJG9BDPE3lDfZ3VWibd0h560jVZMFHQ0IKBozVAAWdkK2FtBrLPOwRE18mq/v5pl5IkF
MyK3e3qYb75iPWzSSuy/A/var2NiN04x38eUchz4gLTV6M7VDSpLrl7IUPdlfKy19lTr/4ljQq21
z9m3/C/QEIUg7t3q5BQXwAQQSXIY+SzeKNFQKkTlVprvd3UDnsEY4Dc5ZjcvbZQCIHudwqFVxjW1
Unay4pgjHFjsvl39zrnlD8ozARG7vlU8CwBBXE5GPunj+jZKgS1dbW5qBquIR/zb8Q3JLecUyjeu
3KuJw6ekjK611y1dVwy/XbL+HpHSn7Gpzwoe1+XjyqCAoP4myp6s23yYzCYRuWlEmI9aE2Mx1Ya6
87hyNHukETWLlg7cvOxrrhpvFlVzJ59zjo59q+BG7yHrk7XezVpSLpkl+68b8AsWidxcFZ5oXiRE
3OYkRwGfqbQzl5diFIWKCZbjXs3klV+4w3QHp30pnCzeVwpRw347cfiHNK9Y/ogzAOtdwhhyakXm
6BGNwUEyRTKxrPod47sD32+E/7YTSXzaqpICKLkkPbabp4y4TSubOD6hS1tAEmxpGQZOHcnAmcne
Z/73YQLrjo7QldSe3/ahy3mUWXBFElYxR4A8CuL77/mFThQE8OW/84v3TxQ8zRxT9Cj6aCskqKlH
a1B/VD6ybQ6kvbSEJJc9xlR8k1EqshwBzO9xzpWp6tn4wPc6OCRzJ9AyjS60HkEJEDu8/XUIlnqF
bX4QnOBB1oO0iXpJR6XQEaJuo79TsqYNcwDW07X5HVbAtySUdrt9be8tC+4Qchn84YmJwzsTa7si
xRQrwXVS23w2vjjef3zNycbns1Xpf4oHMCqeBmD0/udfMirhEyU1zTp6SLa+VjHp+ZUm8M6nEGVz
cegkno1GIkfZRFF4nvmdhPUegvpKJfvntSNcW4Y41SS+LI5IBgFucJ5ZNdYXWiPrzFhHZBNGDk4c
GPZOabUoCbqqNNTHqAcR6VLJsqoWMV57lKnqQvAgGViStCDDAfmCA4lDnaVEZfRL09BSaRPrLV0Z
dT1SuoybSY0ZX0i1Mu9Y9md1HAPGdjQ4utDI6gByfMX5a0Tpjmor14OLKcMKPdkwNkCRIYaE3Vpz
xAFfpawznx2vr26pSS35jdnCHFg7ZSowk0+kg7jjmPXBM9XwEx2g+MgBY0Wk6Nqkr0tAEugxwphi
8o2ygz3Q/h0wd0ui7bV2Ke7bMf+SQo8Ief13jzXGEfBTaJ26A/FBCvd4RvSatU4Ob0To9sE6NV1D
BUtyomUfg7GaP9WP1c5DTq8C9mb+n742LR0J+D2tZFDsXceGOfqobVm3PkPUb2qMhW6cG1Tk4urf
9kvvVQoWNRQl+L17myLIsKudXh8WvCtytjH0GcPWDtVLwmRTpLmLJMHhR0AiRj/BOBaJ9XUWcFe7
7DNoeYv6Ki75eTvSr8iEa+vC0Otf7zQNdG4e72QEFr2AofjWC4TNGPCp0SPdb9css1H3fXlBQDVW
zyIRFYUarL1eZ5b+xG7NnZcuatSWykUYWJXw/3pFAZnXWBVJGAa8QhFOZf8Ts5UrEMsV8UIMaar1
UfmDPkI3UlGALMqZ5oGJOqyhkPfKn3fACeac17OYGFe7q+GdCjDZNi0tZet5TLfU3ivH37ywmWep
BAt+b/Hr4bz6gvqBYMl8dCZRHDO4mAw9Fsyug0/SHTYRyi+3qrgx6tQe3QvTF4JjKvrpMxyLNm5T
a9HkqwkKlFLGrDgNWjzXKvZ288nm7VCy/bop3TPXLRJJV6qfPljRkrbVYCFolNEmS1qOO2WbZlMC
ZgFoYbgJ2vwb68lLd5EdkEfKjKPaOVVMJus65gS0HjlprxZJnQURnXJRlKSUvz39Lv1OX0y4yueY
h0BCUqhiuFDlx3I4rYaIIWvY7Ykvi8ChDXu4R6C/4ISJ6eUxxg3bPkZmNRz/NBlo+f0vsFsE+r58
RHjNACbS1AxpO518o4oX5cej897WHclLjo842IzKHrY6j9E89FRo7Q8eVTG8YFsnHW9aU+AV1l/D
pJEYI1pgNzvFm3pnionm72o2Emr4J+Mj08fr4A7Vx0zjxk6k35jGK8XQ1UUiiJsEQEga9wxq45Bx
kDlFcMoLmEEoI1T+1v8pn+1EDlYgyoxhHrS6Gp+NdnCtS5sSS5fwwrki0aWUFnUXwedrmP6tGgbj
wjs7joTSysEygF+MziyeI/Azkmr12TWThux6fqVnHyVHW5E94TEYpYNaG7wx1o/W+y/dTXsQqPa9
nqVnwV1VcKffmTaKyVNTjheC9HEAsjOeSsqMytuR5tHgIyUKAxbILR9FCp2ez486KDwGQ1d+rh8i
2lqDQCj17G4RAmfgvXoTMs32hKTByhhdLtQr+gONzIT2jYful0pQXjeprpWv/cs/NNh3dL3bF8WH
G770z50OGoryhGcthn0UUKahmFJ9UAHcq3Z5ClRUgYoW/CQeurGFmjU7e9y9oJmgxXuenV+gsXsM
KjeWZlPC+7RImzzp0oNPCEho5JMEDSuBMRlm7r6xA+M6Uure7dSzn/VKj6CrkfHy36+k5NIak7dA
7C/JQXEgc7ae+odXdnP5T77CIpEr8yH5KX4zhOXyHxvGB5iSYsinaHjd9WBaztRKBNAZRrpIYNXk
kNvuQ8I+4tP1h7P/yadciyoB7+m/L7ule8X6yE6svdJaNlt7L4JMk2wCe+sNhOnHoG4HfDKvgIiV
pqu+z+coJN+38iXCnAC4qzoN1LTj9dEXs2Q4m421kT+K2IoL7u7hYNtNPMBBpbgaL2YhoY/vJITH
hR9uFddYCoBMKvRZ1aoVagOTsUV7paqegT0w3vVUHow6FGN8qXw3sOfz1Dl5wyvGP40kpf4aME7g
Nktmm7odjeF0/jw2porNjkaRpbzcE5kwtmckkBLULN04xWUIvLAak8/6mAG6jePyrHBzzMJF2HUn
JHjlobjU9jQCsGYEIjcisWD0dCqRIvHWLRWphXKav16Ch5Zcbg3NOoWCNdDKnszSuXActgjdcF8R
0MvEf3780neQoSvItJGfTzOmIW4KAwO6mxCZoFUR8G7+RDxOcg1wauXuA/5tuJHhX6rMVgiSmS8R
DmrNxpfOpUEJnYhQKleG36pefc7+NwlBiImlSANad/B5hNEQBzjILPxQ1JFML8jXCKlByn9IYABt
Soj9UZokpJgpF2BJWofbnaq3RM4JS04ktHAAXGmypwUi//NKxvYPG6r9sz/XfjevBgX+btqfhYc8
HobgI2mRzwkKkAcToJG5GNdmHpPh2/1Nz5smHw4uyC38iSLDbLzGcxfdS+L13AmUhPZV8xyHvwQI
Xs0r0scCLjcI9HkcLHaDP26o7JM30+ovwRc3c7PlNGHbfu8UKE9qkcmoIpRF31kcq3Yyo6lQo8IX
0v//rq+O6LE2kYTBfLlDTPQlZ89zMAQES5eNhug4nypo7uLqJYX94mFjKHqoeDpp93xGUYYNxnAl
8sL2QMCVoe9N60zQrM7HElT9TyiMlX6h7IqmArxAcLoZ1ziSNd0aTfFo+geVolfPgZmtfL7HAtcM
lJ4lOerfOvzd3JtH5tdLO9V26E3J28LKxwWe86vPVotW1i2LCs6DcDa88PE3dNU702SK7ohft1zh
vZxZjwRj6qmgmzYCxoeQAqqDbAF39hFt7vkIzyfXjyO4DI1rbf11Es3sL32lW5nBipvtOsKZHZfs
xG0+EWMXDE3D0SeVpFP1U4FiuZCpELQGZGG6okY01E83Vm6fJsnJJfKNiTBZJVJkgote6T3FSRtD
CGRHMxU6cPnBF0dMpBA0FNLUD0eBF5b4jKODmhcif6XLyK05yunHtsMs1qUDHD1PK6xWrSu9C8Eb
TtzDBn43vaWWI7xUXGsLx08aC0PaMhsp1qg2ptvOlTBR1usbtYehEx52vkPu5V/ZAeeGdQ7Q2rBG
LDff/dp7DPCyOVNpp8AEfcdwSoFkffqc54ENNsFu2incBTnn3vpsBltqRCJsMSP0hMVQVOukVVfk
yf0GnAJOCo3CxwfePZNbNx84bq7IKymdo3xQOo7jpBKbWjjyW7z3yeOAB1WPB12mICn4Bb2nBSSF
HxrFU8rvO08Z8ovKbEHJJ056XOrHmL4M0sn3hwYixjOedKD8GcbsEiVQGxh7KzY8AVVAMqMkjiY/
klWCEt1DGGlbrfo0kiYUF/l9PMFy9O6lIRqH6xcLvljw1EsIpvfhqHK/uE1b9TPZqmOkdTk8NZxI
VGcaCRdR1hH0GstzDOfPFVnbIY9UFVqrWT5ocpw2guWN/3Z5kGlO5PmTA0MqARlzOTM/1plnjmLA
pHjk7YBM2I7yRDqdibhgeN0Btq0WQtZec2tSuAI6dd9Op5bPuAbV70DrcTsu9azDDoQh52kVoI/E
Lano664bBDXrpNPPjeiDni4KtRdITt0oIRJIhaXofOUq0/kN0xVhHRsKek+vpqlWIIUdD1TnYweg
zkOZCnoLmOmpAzp8yz5DR1ic62IQZ0/nrFld1bCXrQJeIYRYvEKZiuc7jcistQT2fMKnAk5DC75L
hzf+c+CkR8vF+Iu/BdRWdQzA4T3cu0S3GNJ5SXmiHxQgzOGTlSYyyyY8Cbi9wc/ML1gHtJ+sjOaO
y4avErYWZNw0E2x3DY4k+buS4YXnL80jUOlfXUSS1O8MU01x8Phn7RJTbzOxt/E2Sr+MRRqe57Mi
Qh4y9d0mo5d7USNA+aqgtnNpGdTF6Pf/6D+MYdlvKBcXdxm15UtMesq69aHCcXkdY7A8LLcjcOBW
cEdYxzhzK+ht/I4v904tx16hRdWKky0eeeBKtmd5anF9rPF1+CiDozDdwhDa/50neR8fDdysL4vj
JnfnqiG9zvuwrjU2Uxh6jnWrtWmzK7VE9iIjAGQNWVecu1S3fHEWXBfv3wZm5PRuiJycZlAzFWfy
MelUlGBDu1MlV5xA1Ex5aDPd4zq49zizY/Wxmxrb0RCiP64qktxakVguM70z2EMI+HEWfNCVFsyK
SGPWiqdIAbL34ca3sU4FweDQYbuUwVCmBDUhAbfO7MW/G2lfdodSXCqH3LhbB1ZqBUpLaOxQJsAg
KfmG/++JdJnJTclZEubFuYCA/uCIJevxt+WMQp5KpzpHmlI/Ffjma8DwOrYVYjN6LOTvnbuAVb/d
vIqZaq1pW6HqaIY6iqNSb9W4Bg9xrpMqZ0OgYs90pLKg1mthenouMGdAx1wKo3Txi5oLqx9aLud7
BvoS5G7ZdIsPYTqjq6g9mIfjzfJtDkZYwWXAS6KlP+3oYLSCXUxt0M/4iR1TqJ+AtFbN5HkULR4N
CI6TeZ9q06Z1ipuZ/xhDpVFq3gkvAjT83Ng2CQXY2vuzSDbcw7fCbrLUGzzQHosDygizXLBFHxfv
HZ895W5BtkU7KjfeGQShJe3JxiVs0g+kjHO7yKUBw4+zQ1P4dGXA5pDkSKJkvfGlDtlA6UkK/m6h
q0NcjehhRoL6BkOZ5MysIAFr3aW4+yHfJ2Tn9wdskWsWj0i6nST+nmnbjs6C86+BMkwOY2ceaBj1
HWMMyfeY9Sw70LcuONifZhOMuGEyTwz+fBNhirYVUbxOlnYG9d7eG+OZldFzwLGkSP0fFh1aBcb2
BtZ1sz5qwk5q10yeoaM0PCJhi4M1cdhN0oKBtSNQQ6wWb4+K6USU23jhuTd3hWy8bpgCgTWFbUb4
SqbrTzTTfOE7TYA7Idx2hJH4djP+7I/KMwCklHEtFZJlZeVbndpJqk89Mop06jg2Ve/natXJFIZm
bA5berZPGnV+3YRcdoVUbRxNOIgbmcc0uN/WzbYWItGx2cNIh69vXrzFUI99GBc+XaGV8GsdrOfX
8Hv/i+K8zvImpwJnn9vWGyIaFumpiyYNcuhWr7Ca4OeYIanggCm4ZFreXkiMVAw66B14n8OQc/tV
NN/xfRUXqo92fdwIF2TlgBDAtky/a59rSj7epQXKUeRQT1oGzQ4y7fiRZ8h7vQamTVXqczENaUJv
Ruzkivmmg/RuTbUR8ILOzkBP44s7ynvYZHs3/yUWa1W08vZBRfHUak1EJSsFh1OMlSXW2FCo752f
0ujG3EAAWrMbXYKlo9uS7bVNo+hCqK0Y7ee1wOrQBnu3b2QkiZfmErEI1B6UQ4GrrCsMPjVOS51k
D5Ws0E7pqbayoA1v9VNFw766C3G0kMShIJmMj+cleZeEVVp4dtvBdhvM+sa6RWXPoj2rzRdAD8Dz
TOhERa48lQFjtZkMxXUSoGrnIHho0oTc0ZibI36umtiuC1Bsbc+VbCRXBcLWSCxm7KQ4xiRIx/Gx
03WxI5MbvNFq6l7a6prGv2N6GYEHhhQbv5ZV4KyzhvZqDorkqBvo8U+odZSnYwCTMNqF2vux5dEW
cZK2R5d8c8R8X4aSVhnI3yntY9s14vq0KlwQaoE8TppY+ySnCM7H5a+G80oQYgQscQD4stCzWD0E
FmxinYZ7SDq59/2NsmqKUlJigSDnKF7G9ow8AJEuAdW1LA/7pYkK5m0xMvMtJx82va7WQ3fpDtAS
CuwlyC2iiH2i/o+qnKemk5YHhqYT9P5Zd0vKNRF3eQy02slqH6tavekQ+Pd9JOak1EsOj6wkLrJh
Rndr5cPQMoBoRUI9U8jqI6yu5edO93YTnr8aNGP6lW9xERvmx1ZaaW32QocBroiw5oN2GwZKHrvU
RcjheKgzNYvV07NaMrFNuYdyKY4EMmQ0qWFpIgQYQpAYadGM+aVoVri3d9rm3tuLteicMaQET+wK
ERy3H1zAWQ2a8w19+A/qtFv5aC9vs2dds2+BQ8wOiBz10pbAhCoXOdcxuN0frE9r6ZkI14iNDavl
ZpzHQF2tDKOJD0SlsWuTQ/mMh4VCTcSmRuJi6OwdXc35xZm5gG5eUoWP+HODPtWb/pfmB0BPp3sM
Akh2CtYSi9c+rZnNymqqg0jdOMJJzaMfWjxxb8F/ODLwRbRt9HCGS3+3m/JtGobNSh0LB6Z0aOs+
ClwRf1ZebYotu4xiRgmVrx2OtImyR0OqoeJH/3cKmmrLiG8WMTxT9b9mWmaqaZ5i/tNFAoLt4aSr
0PZs2D8Ps1zdxn4XT7ZIbbpdhG3XWKiXh7c7VW7ePlG+Bun4xSzkDVqC1jhh7T1CgNuT7GwiiAdx
qcy6ODAQAxOJUalsOLhH+fLnd6+Vwrz/951oBlQZzkKPSEq3Grez9KpHfGc4v9+E1+nw+OK5y9gC
00RAarnxAO7/+CBsCMxY/P4ZDpsgZLf89gjzjrtOJy80o5bhtODqixsYN4BpJsMa43C5+qs8AHUC
w1158IqP1JFEQ9uT+bl82Bo0XJ3OxeOGEFT76VtCTzsD4H5zQ/nTDUeBk3nuxmepO4xsXUJCzI5L
a7lhS4wG7+6WFiyf8PjxEEbc+WuPbdH+L9ZxcYE5GI2p6qBggOWhEU3guKSh8dfTEBjS+Mhbkw7L
2lwl5kiboKH4Zh1Z98iHhZ18Emano8KrNMbzIdTyuuhJMWoxBjZi9fI84RYV/For3dENxbAu0FuY
yPYfXc9LzIe7awxIaCp+5raiJyY+/ffASoec2hVoTnL6Eqp4w2JUj6TlRtcZTIq7mtdsUcm0TUdp
rpQMnOh0ysS4dWTAoR8pK4+vWGNCh2ld4UZeTdkRKvSMzmILPlwmiQhvT3YQfMy7/xPg6syCSe4S
zLK9dj43tJqE7t13GjJUIe5A1fLN0+iRmjVxZMz/9hqXiaksHiwI+x+k1E2KaCJP+Dq2MUArf6p0
MDjF0vqS5ksw0NepdK5PEN7DOWI6x4qVv6nf/cI3c3Fp0j1diU1yH6N1hO+YlRa1ekDBmzduLUN9
NDYlUghV+9EPIplqAG+LPErsjwuW7AdLQrdcGjGytVuj8wgVIL/rynvzsQFg80PMTmhQYQB0Ia0x
1sogvlCMnrxC56cNx2428XwnPw4HfwNQ3Gir9XzgT956PojA9gPkZEUvr+shs6WssJmeE7cRXlly
IydKqHg8pjh2p9vtEL9H6oIFg7BsKwBbNK6+4ih7ZClMAwTSJ3Wa+gUubiA/TGQPxJ+d3hekSu6e
C9Dr6ltTDN/Kk5uwzzw5mXzLfxMJ6QVN1Iv8+vIZq2BCFybBrroPtjAPg0Zbhu+rTo2aSFxaaykz
fFnvf2dkmvVyiuqkvVponhjx7DkucybA4OnaEwLQuIw1LvEjl4mXfXPW34I8bvH1P4NxefEUKtuy
9oh9hrY5bBR7YdXyQ80KsuD7AXyDXICwlZScF8YGOr0LX6f+Km8UWwf7vdD10lXxPfGhjc705MAL
PCVv8Zhdm8D+8IvNu0PCXpWETMmjxsknn5ftjsOCDS9BEqeZ8zarappyrkOfgTvN0jsck9J86jyB
c2Yfw+DWD+LqMv1pV/yK8Caldol0nKpl/DmRTbYiDGx+5jWk0Dpcoh5mIa6Or+7hIULlXUDMtE/8
XW4OsAm3vZDmgzX8YjofHyol/mX/bwnTVMvhpiv5kOzjF5SLhbWtn2JMzacQ9ghElqlcXGSgzlPb
DOwvRduK5csXF+ZakXmHigREIFpwmHa1BdlxT7lKTYAL3R4UvqjI7ywvRYBSCrRZK/txWCLBBNd7
rcLhF7U3reA/2lEQWW7+01aCEIBCY/EK9p39pMWzllzbkd7Yj+RDUAWH+OgBqHNanYancoWUevwx
NTvvfdNxYcxhRMHZEkdBid5tKsTAbSyLA3o5JPie3uLAoTT4R3Dm9FfPBN8RphMktT9P8QooPM+R
eJZJzWH2KytvPrmhBOkonRDoBOt2hxxWSBp0rYdsOpaPjCd3yhacMCxEPw3E3+OSpqf1VsSxmtCV
gVaZ6as0WhIah270ivOkxIXNGcWe1c5bLXWH6pxbr7bhwMcdVFnN/4sTSPHq3pKvja6nI3a6QIt3
IljG8En8lXkrKEbTzhI+Jl9KBKJX/SXAauePPgVzf4bVUgqSpeZVov92nziC4tQRB9OykZSHu7rn
dNRIkp1ClUaNWQx/5bDam8DIPg3FzZFeMLZrc5fvrPaYafM1alwjz8L8zcT39ruL3RCS5pVVXzB7
N+od5MgMr/ShV9PyhoIhyTxm8X6qDmSXjIyEy941nYoJq54t6hpGG2PDr3B8dgoD0YbAYUqUZnEl
iBscn81co2+f8Oiy1UZ5LiDuvSCZtR6zs5rWtq75FlJy4CU/cUMym8XiIar5mo4UOmlnfVlPT6uI
xP+dfeMFQXM3tmm33RcTbG9Xuq3juS7B9A+ZLwIGMLRn3j6twDl5PgCmG0lW53IBPFRC7S2frCQP
VGZzyxcYDPsuybnX1+9cygmxR+RI210mc507j7HDLJbdmDYMfhxhZus/fJnhLyHsPbUWXoXWmhY2
gPLzBEUJIo5ZNP02eaKqsfOHE0hh8gK9E50WaPxUKwaJg3IJwXGOzZE4xm1qyWQABG9GdRN4g0j0
DR/5RqFnC66AGQ6Trl6a2e5eTAJHy9zGXgAV39k4447tYo4ELiU1vfULa4VY6hD/E3bqO+qEV+SN
V7rlD9qyz4J+FZoVNGNdBDix7nE8OdL+9d2I1nnwiHBboL6hrMwHuTBtkxeav3Q/4NXoqN56oKuL
+FbQ8i176SxchX12qkl+awPwgaalaC1EFIdwwrdiWQmsU5HSx9PtRiaZ1oQs6B//F9rSxKRZUU6P
h6dOSTVUl4JxmR8tRhGAjf7FCXJjmGeCn/ODX54rOAcHsgeODpnFhbGJUdfYwyIzrqkeda7R2eZf
8DcqhdlIw6jA2IgbG2LRMqUMpNUtnn3+WxK4mLiSe8BTKcWVSgc3+MJ/yFOdNFgAdSBs2TOEAbHj
dwMIqGKEvD/fyzsfvvRRRnVfGd6KsWJ5dc+TCEdoZoA5iDutFZfllOwzj9x7C0PO+8nMD12rezWW
Hi4Mkyg0u93KvCAbvhaNKyH9zfPJ48UVL1s6v+d1YjsORSg0Duwyirn3sqMMp4YBmwj7kbkDv4t+
kOHkH3GHorWEnoC3/UNDlDGT59X5GqpyVBAMfPT/d8CbvxvfQcp0Z2Zv5Rs37/IdJpdOO8PFwAzq
XbpoyVHYacisyamL/LY8jUilSuifaEJIhCTypvkdo+NYSI1m6xhb2eTWFy9WtlJsl1UFr7FL62fq
spUeIw1DxK8weE9GgR8qJGYNqlbt1ynMsh3fv7/1dlKDcG5Cwqzfi/0iarAMryTvwfK7M8NEQptN
RlSozgQd7ClI1Qkmxn/a1lPit453aiUXoFT0WtHUYpHv8AbvpdlfTL6kTQN+0NxJIRkxIprj5cYE
xRTCTuXb1dmTJfkWzAHwGEONG7u+zUVQjvnoPbpqqs8wcSz6qON3dwtrljpWMiX5+lADqqvOChQc
8zI+39CEtcrbrUB9t8HaIzFy98s3i4WdGqKhww/3umoXghFXAfstmOhg5qdclFz0fh+FdV6cw15y
AvnjW8hxyrqlAkQnWIdVp3uQ8/THiylsey4L/q9OntQMnwTYz7/PJSxzXUyJUc5I6v5wyMKOI/t1
NYpmpvj7di8KlQdQrLnzv58q2ZAh2wZHDpfzIuI9/DBbEVoKa5Ap27CPWmmkMXWswzkFpP5m/Rp6
45/wWhaL4X3FVUq9crZCi1aNiRwMtw8KaM55eEnrjJg1L4j34ZsSZwJ2hlwqC2bajU0w3iJSb/pt
F3w7s0lelbn9nPO8ru1ZXjl08bx0hSVXwnsk8BNL5cjlh5Qw5iYw90/oMHi/IelBTQQm5TMHBWSw
5q2hXeyapwNl/Z5raYDPSijgdNvnSZ6FkXzGA/xMDaYwEtio2pJ0R20oKNQlsMMHDqw/Fc7QHf25
VMs2Oi8tJiPScsVJO+ZlROMNFMpI+wc+JrgFrZGcntcwqGBzsalR22ne3yJTyl6O7UbByc3gUuRG
BfhU6hK53kjCUgS3JfImIAr9PlpLKBYL68RQh931ilsfx9ubZw3UXFds+bgEMQ9eheqrR+MvuzCD
LHvp4kIm8PLjeEimIzMyIkNwCV9/hqxoT7DNN9A2cMncjToq5DOtl0EWDvBXjUo3nJFJTaSnXSLW
krDxO/ywVZ/1aY0mFPbZBZGS7iRB117G5V1VwUV/11iH0JQpJEh2LPDD2OuGohPZj/tcDteuK7ha
vflHGY9EO1vH5KfIfcR/DKmhkYm7tOPVnIIvj21zacffFwkashZ8f8pq/3g+FGSYehLdhsgOcqCr
gEIkyc1+TzjRmLYdBQzKw3K5vNLMItg27X8qpEABYHarcNQMrpf9bHr6+JyVlBm6YDaTTUnRuon7
9DCagFbY698SDH8pACZbdMXScA1Hpcjo8rVgH/jTInRugYTLgs1KIjqdpdY3lQ/DOTCPClPnAIPT
d1WvdDaX/kA5Qq/NuibJFlDliZB9Ccy71W3ANCIpeUzgm9+MkdRFYS6f2D6IfBhtDDbMBWJeSd/k
rVIP4WwSFjdnmQn2e6Zcm23/HqSvwu+hAnVGaJ9M81BAVB3zXaT9kRHlJSOzYYklsxREUOSGSnnK
8zEjD1aegIzJOAzzHufHadcCvd1dVAK9qWBlF3ZOiRyFz8dZc+cfM55Aw04y49LiJEuR8LmYtut8
h03/9RGWHGTa3ppXgeyJeWhZleWi0b6B7/y9NIgExESwQg7m81GFNmSfXVi4ZwZ85OP/Pu7BN1r9
t3RMKMVmIQTvMaTHHINxEuF2qlRv3mDkaR2hLwP4tN4DIIWK+d5JILI1FHd3lmBf0tDkFlto+/zA
5uWmkkbYSPpazu2TEIpgnkwNVg2C3NwBKfCoktDQWo0zMyRtaPi06iuXqvP8gqQVuWWkCPBKmigM
EiEHbbzlEGvjUfNWal+zvGWI5RRH8jqWbrGIZZv6k5Y/G6i8pHUg0Upot63wtzTYTCIMiU0hKp+O
MseYjwET/VwhGqtzM4XWAO1blqkxS1si2JHXs5G601rtsTW6FvhTCFIubiJpWONIKP3Dp6TFMyP0
dHEIIhU0rNH5OyNKTak4IagLek8eirLzZCic7cNghy2O7qyrplYGIkz64THYAzvS0Lme9YThbGtK
GIEjJYBrnynD7z4UMfLKhHGrlw6hcaTBtvDNRJTQhHajm2q9Ncfr6YelDLUmICoZJdBqp9OvITyd
+j08AlerA3kMCwUdliRmzoGUuexTK7e8w9PR5TEE4oVfPMLWjT9p6gXNort8aFydHaJe9ny/zaAw
wvTQbRW/tCL9eEg1PSCUiKUeYfXzVxI4F3hlKzyComS3xlKEqkwg+IyYVkSPO1XEmjXXyy7FBQIR
DeqfUoYI5QLIk/XAEHTbPXDbE7gkvGv4uYdbeaxrEpLdcGbDAjWERd+oCxqzk4JJ7U9/PAY2CrgF
tw9J9yFlqIrs6vSDPaca2LHoDiU3qLGLqUbx1G3iIRcNjbEose1gcr8Fx+DO8Ces6Jc68kVUlEeE
rNsPUS/H7wfT6Sd9yc0KAHFwXm7cdMAxZTg1FxaUAo/UYVSeLmLVHez/0v49aE2e05lm8f4xO1Eb
DKViiM7Tf4zJQGly3X26ecEw8JMyWB5EC9RgnUf7vscQi54O8qQc+bH7NR+PFA9zaoEwpOTRtJjC
C6j4NRfTMaOrESpc17hu3FgpE75I01BR37UhjkpopxvRwkZGYuV9Da4L9hSM/qYwtPrYZAkqmeBn
HFRrIp2oS+6PiYSCiWF+tLdAXKPV62rboRa3QMHbecpv7WanVF32V4K0HS14dbTo+GKa8pSERjWH
GccmHgyABd7FW6N33tT4f5W1fCQu2lRzAE20ffz93vP+UGqY+cXvqgAOpJMRaUSR6gRHZk4Sc6Ep
3PIDMAG8VW7MUGxGKGvaVysM+QBpypOZK3UuMx2210Yjr5471cCYRHK3zfG28/hFbwvAw07Ax7U3
OUs96VU1Vgiu2/SJOqdxdSOjT9UME1iy8cTfvUUqQIkzYzELXzk62iK4r++UnPy8yiLuEP6x/HzH
jkNqJfa7NhwUONSKrR2E81soIOS3uH9L3OllPs3C9NoT07bndtXom9scMZi+EnSWfoFjSHfp9JC+
qn7RXMSGJWG8CqlGW80HmfVlIRkXtHex5RdpbaSRloAgz8SugbndxC1yAmLKxYKkx6Yndy+gSD7m
tDZZYsv8tGOfVQIlcOrHr9OlaGBsKN3P//EgpKD0mco00/WUnxtRqZnpfx7xI64RL5tfWCvc2kGU
Yaj5qXCSzM4K4pTxqlh/35mYaOllOxQPXubqZ5JgzZT27e4bO7HBiaAvcQd9JlmywsUdDyEbpXmb
ULQ7VypG/Cyz9x/eyRxoBKU5ryQk/qXVZJDqAZjKqq2vk9/2xjfyJTt4K6+KT5sdKMufCfq9zOFc
ny/H37l1/WDSj0tNFYXhn6R9IgPkoUNdAKO7q469yqjc54lfQB4FlwZKMD3ZGJi9RF7427vRrCky
aM/hPPROdLGchLL9ZdmrU3/b4WGIe2YsBtYhssWZsuqfC4Gl93K9OWdDCCqHfqzOZobT0q7vyth3
z3kM+vVY3IHycXWiROB/gLvFzyFospqptYNmKGzz87GVGgOqyoFTxENkWc7gRRswp25dVwYo4BEY
+LvqBKaxtPKDf2PyRw8Gn2KB4EsKPCLXWioCv68kGpgA7j9+uHbPdzRQZI5RUogid0dxNg4F46ou
CNU5UBjFP2GCsXLdTRjKLDf4nR64ikFbk6fLVGZLnRC0FeYh5YrbxXgK4hWSeRhTdqyzHZ1xHmUC
poHexyoO0KUXYZm8Bi442tcHfpWjC3s69ojF98ZeD/JECYz6DDUc/nde4SR9NCCm/ymBzkml6p0j
m7shH46s3lWHAWMRVAaaMmWcqulXgO9AAvKAYMqXlEBCM16lnJHEpHa40oieF1sFvlo0CHdQC0Yl
hktjFj6lHWWuO7pbZ78Wvr0EV/NZf4sEHFA0KlwCj3oWgooAWUAKE0H4LZQo17e+lR4OWa3QjIcI
ZCG3tU09T1bgrkXa3p8yQpXkAyx3W/tFH6PygEEm/XAvfzJ5CJHMOXHG5jaE/HcjK/nRKLwKOrtG
NB6fejg+6mjcIMi2HbLw4BdOciE6WukAZBnGPi9HsvMbzKUdPie+EWr3fjxg020wtUiyXlAT3Yi1
CVkNyvYQqubpXESOFAPG7I1iTbOVKi1DeBsdehUitzscO8qfN/TNXNurEY/2C2pdo2BqF3skbnu3
87jVFQAegFnJS8lq//rTEtoctUvhjV+YcQzEFHI7Ir1JtCAv7Bw9MXVNecsNxvvHc91hyRSJEaVF
cMwjEHhey1kdqhZdIffgmw4mylY8BIvB37CJ6SjV8kYkL5fOMc21K/Y1xV7FhwUYnR8hbAjwAXrS
b0NjoKbegcTi5Xl89JBhmRwU+ByhKvutM/l1Z8kED6AjnTH3oZ1VxlBJTHVaRZEYSSCOnrsv9wqD
XO2iqu+y6oTYQ+kkIxu5Xko++uFoO9VFA+4K2QNddCweEymBNtX5OSGXD9xR8OtDjT/Rpe2nNYQc
f2H/d52Yx9hAufj9Webb4uVJopVqufEIerLdiTSw1vWfdcoZhtcAsGtMU/woQ9yUp+3683esbMmk
5vH4lvCihfc0/1fvgpaHGSNskymGsbW5z2VpvgymhefJt78uQ60wP1rrANfAXLlJQBmjj+TMQjok
+hpLY9AmtCHmM1cyaK/+TM0/8lFmZtkEMr6aNZW4Yphp1/OaX+2XS2BCX/E6DFpbzRZX0ANSKpSa
4A9qOTqPJ24pdgWRrx9PexckJ2mopglzuMmN0L/EX7NAmR3ALuuTuA4KKOZdzDZWm3NYbpflkLek
c4Yqj7m7bO4brkfxJM7vVM4WXJ4OeceUFLIi79YP2pAP7E9mmIe4NAuCY9Hp1oOkMM9S0CcxGHo9
1LjLLEhkPxu5yZHxBmMur8/u5dy30Myw6fm/WKyJw+DISDZ0Mp2OTcr2qs6Ssmqbo+X9cOaGr0L3
RyJVSNMuZSvnnesUR7mcbD/Kbb9AaeBGWFSvcTBr0v3DbC8lVvUueXQoket/po7DNFHTJQMJvpm5
O59JOhO/NjITbq1RH8r1xDnQke1Oc3mV+J7U0X7JGixcIBMy+HDT1yc2MPwXysFTTu8lHA8YHuwx
8gmCPQhmW4ahUY/2e/yrxJMy7HJN+4wLvgRxBnrzGeEpQWafNqkaqQioNOLI5CabUEu6e2tEjV1j
a291dSAl79OK2a/Gwlck9zT1aauJ7GIwimQbQ0aL01b21k8VCWPWu6hxtJz7Xt53Hwi3p6wwWcWf
Axx/henPRc4zTtbFCZVjmQDkgM5/9BqTuq8288qQw9ku/yfh3acUPRL0srZN+rLzQTefEa6RE1Oa
8QpwBWaDvFNVPfn08J4TvsCi90JJa69nqLWJcPAXjwoqLpCa/jTsofR80v3IVqlX2qnp/rd27vo6
/cAC8fEQp0CIGk9h1ppwFX61EuDflqB5aoaVWnaPTdk+rIB9FdGrTw/n1x2ZgOqRpDHf3bMKKUeA
wvxOdjdDd92BD1d8LgShS/7t9+jRl863RDpuMUcK/vDLcb7IwyGvncTidJdCEk9akvOBR6F98+vN
vtxB7SSqCWTeuBDTB24jxwn/ufCJQUs5Ac+sOmS2Ao82sEoGiYOms4SYT20K+Tsm1e0yG+WNGZIF
XutUgNA4UDAYjTCExYJ/eC7sz+Muw8UrIZFsuv8ZYlfUHgh36Tbc00gNr4Hh7u98uoqRjgpwUWeO
nniVvqAxeoMtcRF3ZqcALgaCT1B2NMg/10k4uFP37wjhyJRQTazIyjFlZ/t7+IiUUa6K4ldsz5wu
Kg8GO/UZ424yyVu1fTghMY8BlPoMYtl09hXxKcr9ZwdihM5xNDNo/Gh4DthXvR1kkaJl7TTyLUGw
RCpF96NjIAQKdszgbSf5sgLnoJY5PoQ5RTyqC+Y3ml0nwatbMPi0x/uzqrimPD2057xhr2oc4rqY
ZyMmkeqTdFquMcc/4rjs44uxkES0EZdXk3tJ0A865pMOLe5jjyLKdRuyKLjqw6DXd4N0VoKSBlRi
rMiGF/g2fAuXqfeqCfiFZrOyG/UGpbJYJk67zsRg2PkYsnVVqc0LohwV59tktBkAdDgsvw8ZuXLx
KsvBinKRgs8vYx/Sc5x0yeEKkFtJJQu6jbHPnVrYLcWNFANAim7WRvj/0/sdTMGSE0Vt+pbEYeJG
HcDby5rhRRb/4ruJhc7sDVFEbfBYwyg+xh2nk8l6KvS5ZVisq+0vrM+g+39bii/JMez9cLBMVgK9
d0uOZcHO6i1tkoWtGczD6pkJC6++GWQQkAsSito36293aECTjNOwR4sBv7Xb/xH99dNmcgnf8IYm
HiaI3FtU9iOP673CGXNPYAI1a7ZOg/hFH5sNuWmACSNcXeqCCGt9lyyytwrmbnS8ue6QqBXmEjOr
PQcnSSwzfFvp8PjWnaspWxKEKy2fZbihrwgTR3RyeqYYaDZtdfUcIXa1UyNs87YN5kBPeCVLGxwy
EyBx7J9BImMr8+uIabO/D+L+B5DUZMFBDHiIiIczL93XodAtdIsmUduKH+kBSerwNCol6R/F18ZZ
Suq8lR9MNW13kZ72L48ALUhNdBAMIs1snweDh+/Xna4tSfzuizSDM7LWB4vpV7O3K8KTYhQqqG7u
WnvWYVuLn5RwsT552c+mdI0ktELvBAXDoOubnQfQGAYgh9qwCMvPiSQr37D0/tY+vVg+pbnH7xKx
d7GiF75KkJbzPueFVEYziu2bzcpTdNmcXoIsKcUZ3vLgsTxW6/Jw2Q+uArchk0RtDhyKdrumI3I8
kl6hB5ZfgkITBWSt1VF8lI9l8WuupaUrOGxOUBy/tpbpUV/wcRnM6fO+2Pky/C0edpsOzw46Wn2T
wshC9Sabp/y7enw9WSl65XrRjlBi/s03KEfLMFSBlDJQgfFo5M6rIm4FjxRfivoc3NsqOqkr+zlF
zXC11FutL/Ggmq8udmiByV7SguM27PuNT9kBRgfhHL5N8fM5Gzx9tdY4F+VHPuS7tRxUTWM+bg7/
v8fG3YnDcphtHPRsp213WqsM8KRo8EDEtZRzu0uD5Ge9yiBO/pfh/t7EKM+HnKY3pS8U+fcgWTqS
LsWsP/0Wn05laOTCBtaFcoCLEQJyVNKhBcUiJsOnV56qzsPiPd0oxhZ/Uxfl3H3KJwTKsDCVCCwv
/jRnpYOprOwDlKd22qA4fmkpFvhoV1zzBIxVMJk0byZ6w1h6hXLyYnNCwLWUgeR/kkXE+ns2l7dj
Iplvq5y4HDXf6ISxiKsU9g+zzd/DqoRmnnWyg08yyf5aTsFtzJrAu6HYtOK9vJEYTGIm0CqavzlL
uy9UrmOtpqyu80My4Jdy6xmPqo1p539/GnvK2fOENM0H8Zg9zPJje8zXbDTAcNgmmPA2LIrhBkca
j8MOcg37mKM7eTUbHe/f71oKC3z9MJQvu3IREnTfaXh+st/vSCOpNGq5ihZqyeGGQG+HoRTZhMb1
CjQl+XOTBt6UaCtgzeFXHQrfkBCaLcV5nXLnqnDEGKVIjtQCQ52Ay9455w9+k0HiFirsdIh7MYsL
lw5O/vq8i3AjEQ72FlXh9vCRTgcgMiULZ6w0hO1O/HAeOPn3DBL1aKJh87VJNh97WiJYg5NUZDY7
NX6VI0aeVhdzX9s1afzMgvOubnSk08hzwKlzQt52lLl2GaZFlqZy8eAMwirHjUeaYXZlkVfESr89
PRmRFzWnsO1LiburOoIquVsEKJx+kvA5vpJQFneZBsabayMgMGLw9bb8Kok7yhEetqFZo5N30OdB
NdYX/4aWZnRlU0WDZj12Wt4LjCgy/NK1d3E/dNZnSYeQ23zRhcfbgiGaHhqaD0fgi4PJXd4NAdTI
+RV9gqWws/exz2s3Sd+4OWikJ/xrXEDJrKFs2Rll8OBTyCuSC0QdOuS4agtp4ObivSIOxdVlVxXb
+Ssrv/gDk/YiN7iBnH/u1oNwrxvf//3HBYGSMGo7jnPuawH3TxOQ2l2o31UrwrbBPNrUhE6vLwBU
f84QIkPWgzvV4NaBDOcKe0ojR4kqB2fJQ/8JAW0zitiZHGHZq8WZKWQ72GQ1ERJYla9gjPrnxnIH
CUdrkf8Hn7Zja1pkg97wyt7TEFF1hI9f+ZbDEmwBmOJvyN93F6x11dISksqAmmPbLutXe0fpehgx
EP4l8FhulGd8fwgRHDY87vBk3SqrhWI92gh9p2bZDzH0wXWY7StMQvos/3VzUQiElFrFeftEUypG
OFordLrXw7Zhiiui1u70mfQrk6QUY+psDXTerib9SlSARL+giwL17A/4/1psHga2PRbFxCwyZJtb
v0eDaXU5fjeuUxyaCl+G1MtuyUcpvMzJ9vWR759cIxxgliibBSqT2evyRAEwQXNL7GVmlgE9j0qu
vvaSOi9UpV6CU9+IiUW64C4DgniSsVkIvkXBTUfUsyPHPempoBcTJJV0xuJ9ItP/Goh1ieJjKw4N
2aUO9wpiNLbKclmFCpcKEaw5z/+5w2GnCuNHf5db8Fn6zGDRciVrFDbXS+VvJNYl170gRZ+WKl1G
Z985NSMEekG5h7PPK298+CK5Bz5XxKbZ+aKp11jFGKFDZr7NI3t8f9ml82Tv2JfI2Ad7uOoGk+ww
w1nINlE+JnWvK7rZeMONZ1qWTZ2blf+K8lu13nLf3ggWVAqUYVuIlmNFjwRhmLz2tZujAMIm8K5D
cS6Z2krChyQz3hpIqDOysf8yHTHx7bKMWLx/xOkycGJ/Ek5Z/eGO9k2KYDb2cLvj17/X7B/bfTw5
WvO/rrgBLpKhjsG+dOJEz61VuWZDUnWi1/NA/+vAmTMAQtjHXIWXjkVMq1RoFDtZTDVQAFKADaDB
axj35rebnoztjaIwrAbBaD4Dof23g9Ak1rEXCSIX/B7nd/B/U9bFi6nUlWnl64LHLnUt+AyblGVS
D4AgR/eTssl7g8DQuOBYpC2OSvg4xRNaO52pLce4HNI5t227oDMu4VYHWCvWrePzt16StcByRcsT
imfYns65S31Bqlm6U00Pl8yjL7CsKwalCMRvO2s1/NAzniDlxbn7kHtB5f0Pu7Gpwt9QG9creCta
K46Si0Os856YL7tCl1n8VnhvO08cQBrcuWitO235z5iVPBPksBRT0s+pG6CsSPl4XwtOzg7OL7dt
pRF9EnE+ddE436ZxJgPl6hThbRrJNN/XzQBs11wCNsTM07whYQMR0BM0eGuYTlMLXNEG7FsRWmTI
+WYhJIY/SkbGbEStjb5W/XgOFBY3wi5qAoFdsgdkk1plxPjXj1my42XoWSD0Tj93kUEkofqzG+Aa
H6b8FHaUTh87vvT8EY6UiuTRatQG6f3K/aX+XGIz9MuwM8bs1qwya59A6aOfsh2rrOm2r+nHMB61
NjVTsbnP5nU+kgrSIY2m1PqEFSrD1DZnFSgePlnkmMwVpIeWIUaoEHBObKUfvJ2qCrMBTz+Y5RlP
jfaiJ6+2J0qCrnSDu8Sf7CrejdUna471W/c0X1khtqE1314RloXL7CuHWJp/K+Iu5Rzlmo+nTxqv
FFeKgWAnjTtrsS4e8zfJ0vMK54ZaEs9X9fqRXFHAkhRCFqyyHwNcx3tZwwR/4lrJPrB85ZFJXMne
6mpHPHHWidb5aKcjVFJ70c3TuVsEPkGPq5Hd5GPEgMyytPRs+ut+kZsDpm97CNCL+MY38gg0gc69
U14qhTAhtfsMFKM6faWXcdzYSDLTYfXTypFeRrigQiUASmftThfYY7Y88kXrI4ZRhMyXCin9Fuge
h58yoqYsA3B+QVGHvc0JmoLB51NMPOSkdn87FId0lA/LLVPufyIRh87ObHQMhTVrpLaISVIRevko
XYXSQW8ApqaEwYOYj3K6KzRZwX4DuQjKH6AArQQopYPLtVP4b4xnmzjFqmiUHYmjfPMUD33Z4seN
QWKRJbovHgGCDJD5a+3Dw3BaxyfU3eTQFg2apQf9bjYLTCqmPGFI87hrYW2sUssezC/Oz1v6g+Ol
MjsJIEx4LnoT8DkdaDr09zc2yJIzGBasrymEGxfibxElI8pX+SyfqVHCtlRCpQ/5y7ypKKr/RTVM
v/vNIzGYZhaTWVzEfEd6AiAyfWSl75Q4KherQ2t2zCUz033CzYiL/UONg1OUd8Gea4ZQCHP1Z+KD
ZvJgN1z0xU/pmGq+PBnhzTUVF7/qt4xjvR5uc+dDzMuHkVYcOP0Ym5B6o2KryI9sioPXuPNUS4//
ssjkG17L64ruGwtFMXGxRXNnyOwU0IoPglDy3rVmqbBZc3DPhd3vjcNIY98ORZSothZ/d+odCPDp
h7fOnVWZQdJMgRCrqbgyOIcbIOxY1BUAWFP9KIVoaTP7/ZFx57e2VcCKMQaD/4hdxm/S0vSVcOBy
tJfvIvw1vxtI3QaPk0w/1GjvG7ZE8Q1ofOnU7c8Pzxu/JllUaJ4DQJY8UTMjmedm86yfsaaiJEwj
tPUs0bXEj1ydgqm7Vu2O8bXZSOq8rRnSkliugAuXfIO7HQmedxVJHMB4CZp2NE8ortHdGngGlQZq
tmkXimp97JOUa80W3+MrMW6vy5uGhUfmMCW4PqRJosRZk/jhQoavbnVZ2z0duBb8gdBn04IqHX33
jmDy8FwBJ/Z498EQvte+fznTDniMydZcXuqia27Se6DZpcgp5OWooIKRfyqwEK7Xbblinr8p+yzV
RQX1oNCE8DGH7o4SbEatrvFQ68m/3Hr6d+7BKoqpcYJzYV+ZDC55j13H2CMe+lYaHSpPrjxdBarc
Qdxuts+tGvDmYnlO+5K1LgWLF/q9XpquLsLVtfTUSomVOEMaTd+Uucd0bxcQ5ihkT5sWQI3iTBEV
DWH79sobGJSXynCSCJcTjd2fjiZGrP8wAqsjyt0B5wBXGRhWPTeHdtCXZx/63n5cxX56vsJIzCv5
heEyLV/QR69iznnNtiw9Lvyl9pKm1THmvAiEYnR6MEm+tk52GjgcVociSjLIBewuxFEpEPC2V8H3
78ISa6Ag3pItyeMmWAtZjCptmQQhGCRAVJ9VLXnvWvo//pP8cJ5ozMENlvMo0Kn9bjneCXzKkAXM
h5krpKbwKRW2AoC8tBaPZX+f9NTvmdGXD63m8U87Shf03mMPznUblzF/7km46uss2mzFc4O+2sRc
5URZu4id4/AmbIHsdV8SnvjNF/OEmmQh6K2EdNRpRxVSnKhcN9ORb5rye8mc4EGGXsbqLBX8RHof
56hHX/1QKwBPPTOULAQ8XiKfzRZXx7g3EwWlgOz4q5/sUwA42yMi4dragitFy7zWzxVO/p/czzoQ
M5C1Ji/OHAsNjFbKWpkQlDx+jTwAOC9zo1tut3L51KHSZxLx7Xv6g6Lf4GfG9kFfV3gqTkHLi7vQ
tAWgSFK9EfkGp/QD2gTOKeOc+GyDsUpwdLsnHH7Y8b5fhKMSmyY1R541Lfpha9K74DGihe5Gmmyp
UtF4sB4/kl/sMRXvWxU6H3WSfG6pHHsBblQwRSK1W3Bxm7VBVIN1F5xsCDIV93XDQgY3DBlHxCw8
MrJpmziSl3zlbBPKMDn+fqU2YIrpe81hX9uZ70F2HVXpcqYRFKUOHE8wo3uhXpgIi/lVPxURFVuf
1XYecQIJQOXLVwComOPaWew3GjF7kALvtv8lXgdzMBK07z/sdPuT3iTmQRF7dTDf7VACMHP1z4Vl
8uyk386F+9Pwmb5UixoTN9bfpu+X1purKbk8IY9N4gJqd9Jeif2gu6+Jy7wSnDgynMLXzHlrHyeQ
0IvGcBkuXxMfapV5fRszxNu85QNnJToUS79J+Eoc/qvplS67KQ/vXt2bMPRxqo6mV9MSFW27UYfQ
CldZMlW0DHMYlA/0qB+mv4GLrohpQl9RWHT2Tc9yq/t57Osp8TJ3o5aY4Kg0vbhIHeGthYku/OFU
EPBCi1VlnKvNbcw3HNV9cMeTLFXLrRAX47RC3nf5ZxzL7XygaF7GCWqPcBsw04SMyLn+WfaajB1z
YBTnMwrzdMSmG7R1u1lXMVxAv9m3rWJlN1Lo1xZzy4ul39wwbxFVZLNdq/XrPEeP+3Kbpb534s31
B3h+ubt1lyg0jqqqxBdMIY+rYVohx/3Fe5yJAnoaogi9VBazpxwHXxL0foapIHMQVBpbkH6tO5cx
5b/QkurtV6fAMH74Dhykap0AgzAZVe9Ac3mFkJPFSv94tgcJZPI+sTiM6kQxVEGOV3kZHXYMYE/l
EkxPU3FxXGbeBMyplgxlKmAk22ITtC1DyKT5h3CTFCYjTS53PHSgLA3aOzdwtfpRR+8pckMRhTev
1DYuCOyL1qEPoSb7bYXExLaEjE5sZNV0obfsfrcoeaE7YHQRuSPYRIhjDXxztmV+3t3HzhpzzIOr
MvXsa/KegnaZRAQfrJ2aIaWgTpwHTPWttebiIynu9tyi4EJQSaNTt6nHbbRDMDU8aQws7AqS9ovm
8eD1Eo3U59nxXhq+cLg1rIX7/hQ3Okf/uDJ0No0+ouNGhxdrX90aS4Bj/Fbl+2qPIiJPhKaUAgxG
wmNrJejyYjJSbXETPp8ZseT5TTrcpveeRG9KNQ3RWbq1xX0mx7BMScKRPtm8qC4qLkXEahowbUu1
8hPnnY1I9oIggGT5IKUonVS3SaeyduW7HBGqUMMdQ45m8qyL+TMsomDD0dsz299/gWfY47iuUKu6
jih2ygR9stEEZRbhccIEiLEZT3wz2ZUkl60TohBHyeYj0KghkUb88AkILSO8SFoCVy37g5p9usRL
+ISRkeDmCjLS8gBSI/E/9DKMhm2YCrDFzdUy57UqbbAO7gvuk2Ipk45KMr5/8KSgr+f2CxXKbx8I
WIJRZDoQ0y1dx9XZgTWretFKfqpO6iwrfNkg+Rv6J3ByAXlfiV/SbOKL7zhEE9bZ+mhfY9zgGGGK
QybjMcr3Rk6ZvIR0Fp2wEaqemhjTYzTHMD6wu7kywKtVjINXK2STwCwN99Accht+Jky2T+CVoz8V
rL0HC/uw31kg8UcYFUYWizNUaYb9D7r1jN5jRZ+bODdAfefPxGQgGPMwGANKwqlqCw8Rj2ko9aTR
WpK9DvTHf/lWIWK3PODG5Cc7uaSSfRBS0TqoWwxpI0Yki+oyDfbXTOGaDUShVIRR19Cbdp2nmMrk
iEn1NLfXXbQWwIWaeWi+LUJ1KEjbhRnLNVkbbsM9ZoQIHpAUWC+fQCPfWYiDLyUbn76+kXRm5/Gg
dJ59OQux28KCc2bD1SJ26+xCJm0jjSp6Af5DnlSV5zoH6l5tWF8MXBOwSCxguaFwXP3agYZvCmlf
hSPaKpalLaSePhnhbfTjrQnGw/CgZ5Kp1FsMhCxdnDje4jK79bYwwXV/emwmR8GXpOv4aRTWWD1q
wk5vuXrszgrVTtvnO5gacvJJJeDmJdfONl+nOgD6MAuNgAZ0QkL4KDkGCyGT3PjGdiwEuhb4xd9c
ZDMtcPM9Y9c5Kvbt0nMUd/J2IYpSCsVw5rQO7ZOJHuhv92JEWNKypqU1rxoTfIPA//z6CJV9uW7X
hLnskEX5PMDj+QgNwttmB/CnRc0oldZo4ljBx3N989xC/1QgOdACYEJWvvrZOFkDH5CiZCNEXL5y
cAy4s4dabLDrRVK2IVQ5JIy/weIW/OCymI9iGhWlB+43+PBk809LvMR3ooiAZliX8kv9oVqEbA3a
gKtHWYOKGjdLalFkfIsHJTHdpYMG9PqaJmogM5GgO4oRmPa5kADWDkxyCAJ8v+r6CKwPWKz1wN3P
e25dDGszRcbLM+JBDaLN+0JCgM5OQmSqCwUScSNrhU/n6WXfmoMXmNL4G4bHjThaO1hM+VI71tBP
qfP3lbMS6u3BsRwhM54rI0WrR+6wkridJ4DuiRTpOWDiFqnPqzN1WXjzsTnScN3cMOJa0ybvmJqv
Yqa5dQEsWU/jZS96mvhtHEL8PA/DNxFuLTjXJMxtYmZNyaHU3XXPc8cNW6Wy91LQiv51GVACSy6l
PmFiBSO/lu2/phHlMtuDDU+D53U+y8UduTAbBZRJ9XjZ/xSICLcRDVE7s9BxwI1fREmid9PsgNTx
DpwN1HtqRI12fvio3PsfkNhUg6vzmmWNxCNbQ13Q1J//KxrXwkKDqZQSPu/3TkixeJd36qoVoGGC
HHh87G573arsU40rV4bEgMAGgztN0pC1xalUOt02SC3myDqjLiBOEkqC3zfrmQn44rN15Qqmc25u
JLZfYuViP/ehsFrn1+hoCYegPHMoy7Eot0nyjqW3aC6+cdwE5XyaAT8sv/8cxNb29ZVb8MktYzD0
fgG+ej/cdxbHXqYIbLXsoeFvpUFqooyZOPupAA2OE21Jn/ZFgXB6BU1rO9RwWDYlmlvG3Zlw8kRE
lNAM4I97XYJQ6PZ3YyR8rAUXrUsEistM3XclLB9sOuT/CrAmYjbAkjgTkSMbfQiT8usx99WMZCn+
drHLoCveET6n+XDIQt3AGMGzoWCZlfzw0x6dXTo13YBdhu6svRNm7bGAxT4Qi5l0iR4CRUC9W2Yg
HZ/eNqQmWTC/8MzmpriiV11KjN6vIWHFymoM6Pi75LS9Q2AoFg/mEk+T5mzPzXGuquZgEz32JQ9r
f2OOIbWIlAsJxSLPEdl2Tw4jABKXW/t3e8IVd7t1JBQ+C7GFeZeyTpXOaEjKHsRxQNH82XxH31fK
r89xO0Lv6ndw39fyDLoRwID4mIxyY0vwo69s42LAKCsEAZyFmyd8PrB/LVhKN1biCggID4dbT7jv
cKef65lw5/VvCNVFbBIgJt9qq+nXDFZUQrA44NC3Ww4WyXlQZys7Hwl34jIRKHv7O+7ZdH5wI39c
a5crzuPW/om47MSRg9RVazXwl3p0dkQScado321atXANTPXHSErhNmn325UyEerauzqyisDG1BZJ
L6WiCtTbEoHtTUM4xkjxR2k0un+eLknhoynEh7kAIpRtMKZRU7He7hXvr7eQ8Wk1YuTO/hDqbrXf
eeuPYDG0zYXyyUKvvvm/EVm91VlJgRjzLwGZSYgnMBZ32p8nDxXDsLUWtZr5GykjYHRNuL0qrT/0
4wi7FuVdiSLufn1B5NWAaeDoyMt0x0dZPFNsGlh2SznFQofyH0C71sp/lNDQDsZJnP4HfVp15LM+
JGyiNiY+YvWPr8NfGABr8wSJEJuHzyOtU0MgYkfp+rwXp9dloq9Oo5nBQg+TGMMTMfxsTRd9bgJV
SqVYwP74J/N8ZhdkQQLANJaobOlnWEBSh+m8RBijTeaHBKhs73019xQSShxnLfVDJVfsuJsxhh6h
ukZ7DIJ46VEgF9+IUsFWh8sqawqOPNcsL1hWxAq/t/kgs/z3rB23yaY5T6K2nue1Cu7Di5tnEHO6
IbGRHu7A/KqZiQrk0b2ucJNsekcJZNgsM6oQyFEim1kdzexIRhiJMgOmWkigfdvLfWZtCPI/YFsf
PnUBWVHvD9K/63oO7dfh02cpECRkDFdvlPHufPT8om6iagGWmwv95PK3x/zQmMzU/5FHVEpmDf7k
LzPB+6JDjbftAN/8TRTCR87+heQfdLQ8VmodYZraN0IBFZGgphkTjU42z4il/z/p2VMTfgeUpcqN
5FvIr+HF31uKBiEqXvowIJNXA5vEYb2GaX/t/QOKP0iG0RLG+PV8mRredN+zknrQrC7/QMC/Qrpu
dgu0NL9nDGOPNxaJxCTHcdpmuiVeSI8FBy6zo21UF2PhidD0mDzL4cAso4a6/Ii8xt58/YAi0zWD
Pl76G81y5d71C0oBCDlvT/MDvAwyQTbJoPuIIWzsCObxneo0zKGgFe0w5sxBru9kG0LkgWNApmFd
AZjuUXM+XrTRnmO65amFSIr6UnEbCbG+kckcGejRYhx9oNindFdH2EC/JNVoCSAeGNrafmavUXPU
DI5f8UoG/QC8l3s9nc86cKiuXGrFwYNDjN0Si6WcgKaw2c4KrmvqQCwaAA9E1rQxucc6EwlACbtv
soecmmUOhotDOIADU8AY0baCo+a7ZSUhYkNCivb6Pw52/A8qjrXmV+jEi+4C6TzJfR7aF3oQ5dh0
qHGXO42XvYfPXqGv8NHS9mmDQIPf5Z1kaHzfvpbaC6sDjQXt3uc7dBQ9nOhHvzRX/z14BAcLTe4S
GmUwGlu2DOrfJkL2mudXjHCUu5mswbfVQlTxHk6oclikXoNLGym7r0gCzogf4SweRzBgNyayeI92
Gd9eRIlNhNTvA5XLPAnh3MatsNDwz/dIyIRRs8rlkEu3yUf6+jIH71FOF+X+aYnifoLR9VUH2kR5
NnCB/YECeW6mSvEtVJC5w1LfX3Cncvl8z9Mgg15bYle2hlJSd4LuZkUsBo6OIE2KzCRf7HKgqfjN
PUSd18pH5Wsrisd3sKpqJrvLafDN8HiL2h8AYD/TBrMY/Gdmr6KHAAJWjbgf3dNRgWviF7qhkgac
KY0p2y4pR5WgJfzt/USMj4Ss0z9bV7eBFbl9CH+PPe5+t3CEOiLYE/qPMU5ObxiofKxn+AetMPUu
D3OXjRLuymQMLAKiDEGm1BaJHDBMZxkzM4xn4tXihmUA9eAPnZzqU+AJaXdzwbHDzKrkPfVPX6X9
05vJqvVqyj4w5uBLU3ltHpNY1At6dVOCKLncCNRika1BK9ToVVo00w9iUG9vEb89KceDqM4gzmjd
GAw35m1coLVMgqf1s5PG6GCOfTn9E7OgR6q13bmdq54Gqv7Vupnc/g+14POq4P+Fw8qfVpaB17Tw
clPtnhWmUmH/xDgnKbljdPrRUQ4LAwa+BCk48BgmcOs/oFZgSkxmI1dmTIsVzlf9HIC7QnRRqyWg
p2pWIRTA/2XP4HszXO7xXzb4UvlUOI4geF7+4p7A/Tf5cSFYQ+MJT6ZMG9Dqku4Al1CRqZM7LHx6
+7A+MdLZR/etkPCAZELi1wdCUFF7jjxl4SGsqdH8HDcxtRm6ooO3O8yOs0p5m+l4eZRHFaDkAGhH
cup+Khnq7lW6d54OcIgPIwah7WjVVpKXZxDuzj8je6m8T8d38uHjH2gV477WTOn3+S+yb34N+VL+
8BzQ2y8pLBuZPGF1o51Xao6OoP0XgLxzI5MryEfVizVpBXkd5sw/9vNQJ7oLkSVrxuuTjheTcxU8
EdbjRVnna8+W2ugypxySijSv6/mucD8x9IRoKraVNSWkYU4bNchrRCJ+zFCAP42RbeC58OFBv0gi
1U2/2fIhM/DFhAZYoGuZXVGB9/1dSPxtRBI/jSn37mDWwcqw20Kpul6SGesAvp+L3YP1cHW7mWVM
V8Wp+zp9K3XkvVBM6wydI0/W/3iV611Yh3xalAaZ0hSnp0HBgqdaF0g6V0eWWSRfA7s2/kK/ltJJ
EbPXC1yEPg/bWZ4/k4WVo9Bu8LHL21sFboNCisQNjsotI/OpK3RqfPLZX99hh07jSrz2onL0JxZI
oO+sXq9LTVC/yfAefMNs3QKrcSwn0NYqru1h00HibAIPOjJF/Bcu/pyaH/q9KpILHoX9TloAdmNl
f7uPDxFExubs2OgafzSIxE+111lX2eyHEvRuTQzYacFV3KuWVksFhiEf/r6eOmGQpsBFF+oO+14x
ANqx7INSgpPNWPaCQaKP6xYDqqt2dklWDS0u82Sx6aMDz7raXvSVJ8N7NvLrhm13TREgT5OE1ZQo
xCWIYyrBM2MhY3PTgYCk643kS0Sk2myOfhZ6AP84AnvYtePnxdPnslMLr2p5ntdGA1MN+PF8XsnX
gJfiYTLPfLwDtYhOLQ68p+kd+naqT9sDiyGibzE4a1S514XcRl+JVAhlxvgXpBecelOdTYqDBzi2
UoibvfVUFW+y9iVH1WLvEpQCAu1dwsG9SVyDEZgW0dJwG+vGGPvsg48+do6GeWWmcRq6bKHYYpkv
w3ARy0z58hHnrwI8VsI+F4IP25LpK3FTAuXl9/wcq9+elTr0DLZm6f4XjH9/CVFngUcIWlWLfZlh
gLtmCn6/+jyfzznatyOFkDXS9zS+Jl0xX222Ou7AMBwa6afqUSDiDe5eGLqHbx/kULIm9eCj97zR
IzSUO6MbiZF/UL9m1Hnxsf509PV2IOj2arWRHqiugOMdPz/m/+4NzigviTz8Wm897g7tV0aGKyam
y3lugmcakXuLVLvVdeNqTJTN4mpl0nF7kS4KydscybQBxjLaASjVmtZ3AA/WlX+Uycm4wcdrd8Hv
3dQWLJ/TuOJb/TaeUYPt7RZWcu4F9hjw7VRYQIf0Zbe5HNgvuAQ1LbBAIEC+c88vOiSWJpreMKOa
gqKAd5fU4+z5Xe+nLzTPoC3ucg4N5Tbvj7Eg2P8SJxnf/zyCPzEmxywVnaIt0XRVeLgumVpKIXOu
FzwZ0jLXuRapnVgrS8ZGqbmtF4opneoMv63cVJ0gJ6vMXhpM1R4qJy+OZMoA1GI2/PWSAJMPJ2GW
0NP774yXnZQ2TyusN60b1zBbUn/cuDZG9ThO8L+StOBFA+h1Nv4V1mtuOaonpXUz3tNou/nV6B7u
8c67vD+AHsDZHn+aUlA/z61dlfyOraIaEqLwLdQcIsRZHhmwmkzOFfemlVvt9YoI/ts+/q+mz4Oz
byZODo1gQyEuYEuNoqvUnZ8JdiWzfejMEiyWtpAIarsSa/CL7JOV23HceVUh9hqnvHWhTobXs+Ke
eRlo3+4dcPUBXDxDIR/xd458B8Ir+aBptLTnsqCHf7SB1t6/TbctHOYu08HjZt0L2ZUGpsyZfGFc
2WPs0t3+Dzm2qBDdCOC5NGClqL0gVpZhKXBElJf4WuC0IKf1X6AYYw51JzpFOYxC/Cv6VeVvqxhN
vXmn1AZ94z0PAL4wwdcv+WcWs1eWlYCAyzVzLb+cQFxSZ6HytbttBJzqv2IE/ezrU/oie/4RVMX6
s0sIVbDidWwpXvpHf3JsmbUjBqn4GnfKu7FuFmRDAq7dphxZIztD+cuUlfy6dvLlbjol9+ThUwxX
LcUAj9SInap3JR0yd2zCAGF4ngEq9ue83IPDoA/ZCa3kb6irXUbhjlsaqr8SluDaETW6jPCtIJcP
4I2/V6+E5mMWLz82dhCjkX6euRDIZlesnRnXUtjm7PutPnc/qARPpJZt5iB+GPysZS4W08MrwINC
6KbstJBLbtJjYfTCMT+13fiPSqkjYrcZSX4/WvOetKDYBDjmTeArWuu3NzU81FlJifg1cTuyTvpW
LZyjh1XVL8T2xhh0y9KabuPyKQ8I2RTQ1sYz6rU0jav/yuEG7jhoRRRnB3xwUoWNpLNA1VC5ocgA
LWz+oIqPF5nbWyJLnoHtc3CeK8w7O1hY00sCkszf5VwopUmTpZBb+5wRO9rbDlls6MEWRIftc2Ud
6/LBosMyW+leUPA1JEXss8BDR3cdfJbOyr++146Qx/ff4M9/Kdh3cLmydd7eiD7PZGH3C8wzpK+6
1dK4tDoNZIXlDyb6HOB0Zug70/0jxyDTjb+Vuq74sSPxCctBl/NwP/9A3+lqaaZH6hZwtUifdZgg
5fGFSCoG6GmQZp5gHC+giwzR8vY+tn5wPHO6RUXpkOdzraN0HtURgS+FjyPtIs0XD24htBPssgY9
SbgV6A2pYy6bXdi9fAySirT+o/YtuHWWZsXyE0BLJG9VXgayJe2ANqeFO0cUX2oeSmUTDDg/Ujmq
qZYj/BcPM+t+H5X8YcMm3Hh53VC+cGwHxT8TnCIoPp8BMfiuPo7FqVYG9L28JlBZjL/Me0l/8KA2
nXyxvgWGWUaDCzcBOFns1o1rA3TjvGZBCxeK8hgTnFaEqA9sOKC45nosq2gDJoDlR/xZywqjPl4N
SWSI2h6hpwFvVmHiW2SIr05OQzyfC6QpxFSPSfsqz3OxfXjqNiMWymUQmQDUiAQDj0osS3Wrt9rY
G005Rg0Wiu+sCjfbxRxb0nqOtoO1VSRgI1j5upWw0tFrDdXwbV3UiBCsSTJCyus/tSPB7vJtuIom
7lWi8KgUagyR5cdOm4Px8FJ6yTtUHUfLu5wB5eWZiOyTW1m8SUAUFKFSnu0hqmM5t/isiP9SIIcW
A6cWbWfH7BGG0gfpbx0KLe3vTMuCTKmuBexTP6J16eFT5cbdxpAYBF0IRDsM0PIqS4u+5KocjkzW
TjHlJ6cFsVC6/bBvzK8SnCZgqmNAtHmEDKgfiIXfrcBaNxYreSQA3ICwWRd7MF7XusaMrbW1cTU6
bwpKQ76alP2qFMZTK3S6S8V5h5rgCyozwMcgiatoMexOjRW/onc/sE7YQiKYyNGgWOgJBDJVwN4u
At5+tFEo6E7fXvRUzjtedjvJJYlmVf/n+klmYdrVQcQlg+hee9xEwLPNCGJK8GyvpAHSa/bk4VqD
hTT72IPfVETv3GMhm7qvcQfWEYPzVVUJaoTa+gF+O6HZV4vSnXSoNexMpS2Ryt90H5k5CudzoTyT
p7XY6jVVgB85QsynZXg/jERC1MQOKAxzQB8E6CgHeu3SHDaN9Fk5dG7t24g1qu44p1SOM8ACvDc+
If2T+LIc7ytL5IBEimio2G/kcPlJqUheicL65xR8XxLrxUvVW3jLvDWFx+6Yt9sq7Nt2evUN6gR3
ZIuVtRPoTFL8wUxz9/5T248ovLwTgzxk3VT0ZBep8+Fo0x+bGzm+BVTd89OEv8dZU2V/uwGVrNzI
VPZd+VhDmX84dz1njfSJAeYC1HLehwb16VcTXOMNnj8l5Cl7Y3zfmilghYdC7Hb0uiaDPeFCJ/aA
nNH9UJ71DCurAoxGYygCtc2HclHqeVGNOqx0UTp6HO5jOvNKm5IfRR2TW2ezLtemwYx1Jik7K2fn
Lb4jUnERxH8vPVyPNHe/lPhJNEThgS2x1GBYfGXUC8255RE6oDYxTjhEg798379tcr/bl4J2WKRk
Oxp/pW+rXOtIa2jrqu46UB+Cl+csuNGZB/ZsFK3qnpZC2m7i7R9199OXnnUUOZWdQY1JvBaLPQQL
XXFGXzNOQI4v5D1vN6reX8MtiimWmZH8kHzccTFcXl66fTdEkG2qq/1R23TfUNqXDJSkTO+1KPes
D9YaqVHcYpmMnNPteaoqCBLNI32g8hNHNFAcC1xI3S1XS5ofiu5iINuHARSniFHE9WRm+VyAtSXO
C37XlSjPywFpl9UCNzJbawqaBa2xLyOxT73UzzpssFBYrFYiNrj2xv2pi09Ipd3DQM0VBo4qE58C
+4x/JFRFbbssG+pvDqkbswRpQ8K4VtLJV3LKTiTOQtnKd27GJOT3rerAsmtLqyT/BTCEK4uxnnDQ
4XuhT/JIRIoeNiZUY4mRWvOgSfYSRQbMVCIlWMbCpTuJlorlPmK6j7sGTMA8mjUDyfv1gGmbtEyd
vITAUtEj+tw2wJYsZUaXGeu4rSmI26yUcbhSHIG9FmqRuH2mNz1qiE1N5KOQdpt0iZMw+ofMKuCA
EVsN0pIPGBjO3Oc5FNfAL2xrdER+ReFQw7wWvIVFDOWVDZnkvrP+reb9XGB4kfBVyyvk7DPdSCKC
A56cqF0d4WbifYFQKUjgfg3A49sY3hsg5uRjonxEgnemdXBgUFJzGMLvfRnMLQP9Zyu+Wywa1QsO
rj85xlbeeUpd0oiBNxFc+EqZw1u8YzhxQ5nC8j1USEeeGZu5akaT/+vZtAaqeKHDI94J+ogxnQxe
CwbsTJk0w5+Z+v/GtvEpAsmScmN6iWGi3V7PEeB4l+VvizpfZmfBtoomy4zWgSCkwlSFyhFxWZZo
LyanWPGlbhZ1cChcKBm7lQ+6LvCeZrizP0VmaNsN3rTEF6pQcV8CGPw4eSxlH38lM32DLpu7velh
zqta51sfIvIp8uQJH9xRild3TEbc0fYFfoMIeK3/T9cwkrCegGWWtERhmpH90C+b0BFI1etPEJ8A
PN+HKTGLX3uj7uEw/JBfFuJPJsA4JyfwvlNABp54dTX58zeKXgrQ98coByihVnXo7zCicxoYqWkE
xLeW61rV4doXE3KV5POuIzWtTUkjkN6YiykB+qbFTDiIc6/+P15zvnJMklQs4hi3mZTQOpnX+2Nn
OqOqBK1GIpdjkvxruXrm1XuIuBBuE0NQ3zWdH2P8LL4FvpX1QIUCcGqVd3wBn6eoiL0NcMV0KfNx
hcEbdWIgI/WF3/J7TGL+iKiO46kV/6CNAcKLS3lr6G4hiqLYP8lp4tW9lLKjpt+u0NYKeY3oqjhP
EGm+YeQFrRRXejoz9TiaKvyfHYMkKLygfC4Ce1u3ZekV+tkeM9pt8BnRfkDdeZOgVwXRXWdPxN6L
HmNL1ptkUJA87a3u0Z9hCKfscw3ewL0ciutXB0bjP2ieCBwK7vGzMb6fZ7PpAlgDkUrd+cVlg/Jp
eaJSqQuc90VcTOcitbI3FIq+/aweH1F1Y9RA4Y87rJJ5a+7N5nU66SniE3xHe4LgU1ktC+9f+gIS
+TGbnAhJDgW5NWXg2NcE/6ANrZVjLnqAT09yS8PemzPiB56FhYUbCXqAb9ykXvrXcmT/1pz71Kb6
OsMzxOxav2sDT9RHzyHxkBljthKSUkgpQhoXUeQHamr3OPMEa1ND44SSk1O4vNyn+jz5ZyohZGvK
KHULljWwlLOfXToqxlo1CjDcg0Ootqmn6jK3YRlBsoL7HaI2ODHdc3EpPdNlfNa15oCD6046cufe
M9zhhnGMdH2dMFjQpO0Ti+EzFeN/Fc0yQPC93pjV+mhvlIwwaY0oACcoBa0FaeUcab2xBx4b6q0a
gKvyom0aH72a/52wfywwHhkU6EY+WDgwrbSf2C1aUnfTEU7AljMv2M/QWsSidsYFitBVkDsXyhdj
vLsQ0CKZ2AinvHS0IW7541eWcJFWvbVQmWlVE2SEocqJjxAla6JZrqsyn1OCzuXar7Z+cIjAakEx
Pnxm7Erh4kNEqdsX4JeMx8eCGU+Z7c+YlP21/IOWLq2HQWz0X3gYtm2L/e2QD74iVMWDWEXO29Gr
BqdToqTtlw1vnjaCqTJW+jDCP73zOYOYxdO4SgZVRxU/WBGE+5T8IwJymSxFJhM8W/AmxI7iyunO
3tRchHiOMZwX0Rk5jRZWrT48bnU3ate/qDlFoHtuc0dLc0CvCSaYArV+a6TPjNVMGECJu3+nlEQQ
JOKCoakVaQx3nf/OPsg4clG9aniqOb2JBtAYLOySygbPu7OgkQTC88v8G3aW/+wF8PxFgLiihuSa
+0N8fz9d0gkBjiRKxk5Ug46C6P1rHmM3VKFMAF2rVaoUi/pKKZGxpFY6blb1FvYIZgiRjAbNdXTB
sXFLTQ5VKJg/z+z3YsiVVoHgBuxGdLjcf3MOP7GpVxtaAjPOLfxCBOGUIGpBffqDMF0ziNnQ/IyV
ehwWO0IxARSAtcU156I/dLZJy5DN7TVhpBnsgp9SMafyIRg5VjSP2u+Wj9dOJ7Z2idcna4O46Guf
adSg+Svv4mqfCNeHAAor0quf8vE+08QvV38yOXHlC5w8p9Ccp2+8wl/DqpHHh0FlCl+nG7GZ3aJK
zwiGfFUUX1DiWjFbtffarxuZe0NRFrPfHgbQbExmkXnp0H1/lkP/STuRM8kf7WOapxVjrLx/ZtCi
n5TA4H4GvBfS6gcrY+rvE5NZV3TZ8P+368vCBIlh2RcvsIB+84vWwdyKpZhnx+YpNjkdbPK7/Ego
OlNMYg7WdTQmn2FfSUS8KxrawCe8gdnRN7mAjilSQU3Tk+Pfw3uHFdp2iEQwVwyi6rgH1kAFSLrk
nWaxeVQR0P0keKJC5s1Lhb9myQWOAbwxEgd3UuIa7AR0A7trr0xrOHJ5MZQpNocokeLuruQ6rfJ+
OtqHTevJXVAJWaAisadETNKgPi02d4XviOFd5xhhpt3SmnCaGrkv7UdzPx1S+bS8LPNOHCv+lsIg
bBVimz5HMa119s6mvKxZpQpbuidxEll/yckXWKbOwb1nI+cd0MiOWOIhQbFBWl1ezLRiGxcC0RS3
FdkHN1oOKqGkasp0ZEFraMj37hlcDuw58LZGulth6yEgF5pxN7tadf7hTnqDQY9bqm6xrac9CaRx
L3pNRqg81L3rgm32YaIKD7Ur5JFcH/t01DEkq4qw0d8tvkl6eby7E76gdk6w3avjhXLkJ2gIqejd
2HNFBow2PTCQ0jEggzI/8Xrb9b5iH9TEFkWAXVluP859IJKbXXnt2KaI/b1j3OA8ushnY31AwDGo
uKQKvcqpoFeCb2yBmmmvaK3qh22O2dEaiFe/1BBQ9mA+cZHZHiiHI+jOSie/wft0kFIe0zI3wXt1
UNaQTjNlYL6xkBTju5aZkyX3KbwRy5pbH3zoPfKxGUUV0+FOMGImN46/IvYy+a5grc3PZ4E5rrUE
H4gSNz+Cc0eDnQK85rfS+Yqx4krT932Cc9NNdgsNI5vwKapjisWYx+l2gEjyzoskd+V6/ABVUYhe
bVbRpiftFmiZkFIXoxcrVMQCDvhnpwaaxk0BucdzCSOJRbQx0bgvMJv/ZbbyOgZW29wFzNz9EfcK
TCQVMBq7PhLn/oXZ0Qv53AnLccUILdgev6hnvm3Us/9wiWMfIORW2JUmHLyon8QkyOImTs0N42cs
5sirv7QDtN0Sq6d5UMBbtheVX5dYSAbLU3w95xIviF7Df1hDmNP8bvbMgFnYVXC/yPynn11HCQN5
zFSIVTE4aZCnab61w8yLzjViMQUs+mA9PsindHBdKGEZuHhPGW/WYu4X1SJ1YpiU4KUVQhZRputz
3FVTuMbSPOoYLYYR3vxy2FXwAWkIeKGA9R2gFvOGQIVRceNlM/0mMbO2Z84s1h7EAbEcxjAoFaHN
ZstCkFrQjVSQOHvCDZvJFaJNTWbtz2mp73oo9RmfpDCvJEivh33qVFyzKZx/ZAHf1ZY32I88CQui
15jHcwWa42yJ0pFm4UpyXN2sJ7li+8/oSRpnisnX06O/txz8qMDaftsMubl3o/xrf7wCfBYkF64u
5LsglFcKa7CZ1H0OC4zN89kXS4+gJfZz+ACInEBGSJ85jZSIbcpWGyB7suaTnYw5E+bGHGONXQhq
r2CrzFYd8H0n2IacnF/LaoRckHGqJKEsYqTk5JEzJz33TLSaK3LrpgAFkvhZ4juFL7SyhqOa0F6F
DwSIQxzTDf14mnbQGEDbNSM43ws2OaXeF69LU6Rkoj3dBP2G3XxKMIMjZ5ABhjpnovWGnt66OkuD
3oJCD8kWJfkqZ4RBUVTq0e4uG7zU8F/sIOW4HHcsR1mZbYkFRxVwOI2GK82cL14jPadyTWhAGAi7
X69DGp3DUQfnteoh8Ww7G4Hki1EQ3KRvxFP5s9FiDppmO5xl00bu4JSGa1dv+DVVtr5hfQJK7oV4
JGCuLxM0fEovNMK8T58QB0DDAK4Xzy3B1iZMbcdUTXn92pZ7VQ8C1inztskKt/D6p4+9kG8sH6xb
87CGbanBp/uUk8fojd2LauwltstkTpfNjpPl4oFS7nSAekfgCyXOptlJiUYNvqGvtSJClDeS1YZa
c+aCDhooXglNycv/9teubcZD5v1a4eHqi36mHEaCxByyAJApT9QU3nlxOwk+VrdbDyScKh/TDsiz
4KQs0jRQPqR9y4xMqOseffr5BEOETtmXEvwHuhnUdrW5OSmRa0E0TYEUdaRLkRQhSp61fwolu1Xt
ZjnqHtiYjJbeFtxqsHpfmlFC+TLZBe1hPm9DgH9VLq0M9iF97bbSdGFKh88co3AZ9avRLeqpGdap
y9ORRnmoQU14yi4o7bvGp9TTtxrvBbITjbczBpGYgqaN6BFUHizoJZT6PtQiLFga93m4tOIMekVs
ib7mTxnnmjRXuwsVcE+cNR4+VspmcGZ1gVA5Tplm3zyQqsSDBy+0iqvAljzpseJ5ceQtsIwjQlXc
hH0vO7vajlCC8apc66cAdKdoojo/ZrKNQwwxCecbqZ1kkYyKLl87OqqWLZscRVmWJwwtF7tm9vZU
5n47JicxzAZQo6AN6vUDNeIzzncPFY4QJF1VVCPUScnwz76hDJ9Qt9buRTUsljvgyliJv58KUYe9
9lQZQbY87DsgH947hh7FNm+D3ppwxFSNC6gSM1UKURpPXo71cB/BXUlTDGaMDmbDpCDQFc5hWeE4
oAoGoTwk/aDR7zLKNWp1lAyNuHzfO9++nd+a8jzKmffLUy55HpoZTx/bIAM7qvM/F/R3DVEtpmbE
pLoB3iCLBXf4h1346c/mPNBupN0W14mzaKnWRn5HB0TdU4R7SQ31NuCvgX8GgqlM+nH67+1/0VJ1
sctx5N0YposkklG4AtiDQkD4R3WXJ3lzhpOZul/iF0rWTRT5czUmMO0JzprElQEs3qEfnY97js6y
BadahsVN6Mm2Am3fs9AxHVGtezdKpOuIxK9KPlb5Hi9WgIxG+xbScY8cpjHzyIAzUZN6KK2B/7A8
MuI5XPXO0z1xkiqTo1mmxYk97Bn0pm3HPi/7rDjUoiY5zm5BI8XjvwMY1i64TaF1HgJNeZIbglQw
cpJocSYAO3HfyGnlDTd6yMFLZ9/4cAqqaAZaSGwLIvcFS4cNmJCufLkemkPpCZnVs3MJlJNe/wOO
yWbc/diKfYHp+ZC36TLS6N9XGfQ308Lk8me0MaRsT64f+uFQJOwnWfQ7c8hoVvlfhcpWThoC48CL
hxsoNP581OJR5lDbZIcjsmjNEwv0hFOdj4m+8lKDEjr6WdF8WiFkcfzn/GuSHzy6CL4v+1noh+hR
mVU5a+3iZqaFPtTsh0JZ/tqCa/rJu/1OiErJL0JpuP3ScvnOs8KUVZNRdit9YlWbPVdcACaIlXTJ
OUigpiqyHqAnvJIy6bufoMnqNwkh7yqK7RSS03ool2gKiqKRdQJPJS0JxOEA0e6VKLpk723Vyv93
dqD5LIFy++O3Y7OVLiopkzgUCAbUpxLOPG/FUbc/6tm8ckEojmzRa1zy8qiiyc+ftyOAWpBTNUP3
WBL+VYpW//bgdUB+NuU1LF89Rs8zVVsSQJAhYyKJiPR47RZx3B/wbfD3BN02Y16zoX84kyodeyB2
HpEuxKn8UWFIfuQ7oRBRzolcnTagWFrCycqGgPjqcFWvXhBhqCiv5v1XFcv2VA7n62VqHchGg+gA
3m08mw9pso1Tuly1jCsel55GfoV/HuH5tEDvBlr0MHt18mJAJg5hWlZUxp4mWqDTwisn/vVB7j9z
M4j29zrVjeGVrz9Sy2qkGukcdonX7+sIOfcE8tb5136jPs+vG2ysQ42BC1KcDj1llizMqF1j6RQd
D2UgW9FO2IvjB4/nDa25xxtboAtnre3WlSiy96h3mpFraG0F62ceSPy7LxSYKzhZnWIr+moY2bK5
2uoAepzWi/+aoZ3RTM5L+vtsZ326nw/1tgfgvh7Qyi6lzkha00pXRSBKDQcJ0zFqXW9kMzZQ38FK
QtRTvw4oirEIsQheQGY/2J4y4BCm0mkIf7EbYHSWfpC9JcuxHsiNNJQNk5l+Yb7Icu5+//sJR0ZU
rjHiZ+jeK73glMTIPal5YfvKMBdDIN/JqQeOlR0fj50noNkqB0+w/6tMGMEVdHZevpuf7xa/A2SA
BCZaiy3Ar+8+Ni1jB4DRzXH83AK30hGmFQjxe8Vp9jjEIHOGk9rCtRiJGiKRSoK1XR0jZrZI+oBv
afUuKi6DNu+hyj0RhMBXfbb0V7jpu/d3MKJaqjfh2DXwfbKtidUruRO/Z1vsEzT86BgvqaE4buS7
OmlWlfYEEh60rKz/CpVFnlrGCXpgzRhban7Qsi8Cs4cXR8en/+NXeMb5Wwjl2R+GREDpKn18/nR8
8hNhfDsUInchHHjbw6oSGwSfQnEIXcAu6HjL33kIue1GaBmTD5QAyxRxSp+VQArFpH1q91jmP9K6
/3pCDy/R++DG7UWFiyUjpHoDqD7n2BXdgqYVfYq4EVlUa2NQ3evBk5STc9NQita8vZ+gEy5h5vrE
6IeunzoEeO7j2zUYsqmy9c8Ju436QsKeNc6/fC/Z3ZSDKEaagiolOJUwChgCI1zFzn7PbmkoOPHA
uhFvBL7dOZbhoH5rAqmZ+fleQp8Fr187nSuOCU62SCjDxdsELy1qXgl+mfQVmq4xnwcP5B5UJ4Z4
H1dhgrg4Oo/g4k0Q00nNrKR+8TjAueas8l6nYQJLxE9WjPFZmr1DSluqsrB4AbAX63UugUOZoSav
/EZFzwLQ1c5IECXSWU6Uu9zaUMeoXG/9ZyD5kjvwp6no88CNJauzlWCZre6muUmgVr82KlK+/tQ8
CQYXsfuWDzYW+5EIFZFtuDCwW3ifeaaahGN3HM6jtIHY9+4yYWkReEBaNWGXmXu8bbAGcveykuzS
ExlZaZvFvCDVew3+yixrttvvHG5PTZEx/sRlynq/oeO5d9ZKD5uvmHyYGD3tLcsmN4b/7xGbNqBq
iJ1ZpjdYPgaKL7hRePqDgg+sig8yyC095MrtohaXDC4hACJddoZDZcRmwWNM7Z95UWjrssdY6zS4
jP+2W/3hxIbFPmOjE6xc+E7u9wHnjNnYsmfMoR9veeELFDa/R6wVxkrEL+1wjsHWlBCHiG7zVTxx
laL0TavdXXk1gIblG7bbXrHKhjLU5fLmsTQhYmCVUID7cT3/KQQEvdk2RhTHNjYyScso6LPV/Yqx
Ku6/7ORZByfmu77hbWNY5z3b0ei9jIJLQ0CAkOD4AU5eznBaevYyiHKp0pDA5u+0NL7IaA5wv8YQ
bnQzAqNyZt4+BqfV0Xw3Mjf9QQA1sPVUK2V+EDsPLbmBdeGueF0iD887pzOq0Xv03o5+nMcB36OH
he8F7AewfSVPhAYIs9JOSlmRDDcPNUbV0Z7o0MY48/TfhuT2JuGgeeB/dEyPUMLKqrsG/uu8h806
mo3/Z22HV1P8vRPp3+IwkQpss27nGUfUs0bJpWWlzdTx9wBdqJJyUUmhto/NhxliDhVjBxcLdzIr
wkrLUfj1kvjbmRWa/7mDvgUhhLfnLskPoNN+iV4PmgGbpEAPdpgRUrN3YOj0KMr7zF4lmV3dIjQj
T1G/4MIVQh3IaImhmxjMIaxF0I173ETrEWI1EwdzUaV8XarOpo2YonGxtc7rYSzJUkc/UOXibSnM
sAFNE+zMB1PcjzjHqChFt90Lx+7GSg0OS7xujrFYsO/LhQqrS8UNOMjMGy9JbrNAbhW9vZ4VuVl3
/oobEwDThG6CVAvW9K3cYWnzhxMcRAUIoqZgTojAZ9yd4euHKANpAFviADG2r1Nu07tUF96lKZY3
hq/gmh600XZqILxoRP4EmRgqJtE9HVAXx/Ny/W3KSsC8A9B4b2FFxFn9L+8jYbgW9gT1/+Qj6K3M
w5AQKfetidquZYdlBXkBXVZ7YeRkg6XimDlPmnm0MEyKRcPl0ZkK+4Cz936byxpv9euNl3QaXG19
Aw5IGSirefVUz3Ya7BeEe4OVbQWeZ8X0cMFomSVJaVjx3mL8zYvfsy4Kz71kbFSH1OftcswTL074
UNXWAc90oz4IF6H+XJJz+UPAylSWHpEtRO9hOw+1sbAH1Lqolhi6didTlL6Eor07qcH6TBcwFhpy
/kPekTQ3Z4u9Tb2cRaS7+aXtkumEgaBSNCl4b++MzcKTkJmc75zmVH5BCraGISU4uX1fsC3rfHbF
TXCabM2pwDqsSDn6plhnKNi+l1Wneagd0Lp2OQUcqYrej34HAe9vKb2L+IGSYc6WKmRh6euaZrq1
fEEzXP5DrVuvneHF6Am4tOlcHWLN6gJrNnc4XkVDelkZHLUeerbKdVZqWwU8QHaFqqWpUf3yPlBH
0mS5i/nhITPA/MP3WShk39FEy2Es9KsuT/TZjNslelzuMQHdq0J6Y9UGUTWzLzySfc5sjJ1G4hZp
uOpPPe5wMelDQ8PARj+yu6nDSqjjrr2KAn77Ra8qh2LUDctcqMjHAhgi3fO/ZsGpSIXezIjmRgCi
oBp9pK2/hi/yj26PkH0xPBgmk5namlHIf7dFi4RZTxZr05cwRz0w1NV+g6JopMUB4zw/vQsYSv1I
VKa8EfASOHVnqwCSbK/bFj9lajGDsjLYroia5C7vVGBJIOKZd62U8ohxNSO7whOka4QtPDOq/3FJ
duAP8xWGeDHge5RcYIOcL1UtPfBRuEK9ZeMW9lRRt6/VGApTGIBJN60QDOEGLvJWossElYb9nimD
QOYWxIdrrj0SgA28mCUOgzOcfpzv9RLYE4Hio2eboslv3ZaoKktlX+wI1pQMauG6qOc1mX7OHnY3
4sUP1pPR1Qofp40L9/nMhLG+N5BKe0jeV8pvbeV35c2t65or+PPPFeTrR0ILluSnHk6GQkbPcigK
nR0baiez9xyd+Z/FQxIF6smGT/SSqVwMg/PrdOvhNr/IOSRJbdrg8RaeTQhpSt3+KXIBVRRknhb0
fC1w6svb35iTiHFuj4agwm9AgTM/dxlHFs07PS6BBE6m0hlkxMGQgscI2o9mZjEv1j75l3nL4Atq
oJL3cgRRo26Q6MUwaSJnNo6eAMzFXgV9z/bSfXblo7qU30RxZr6o/ExNKNwvJhlU49GO4gWSYyKc
olnOaEZbrKtPVeL9N5niH1D8zziazh//ekr/vmH2K+/1B6OLf825tnw+zCZ6d8L6k243LeY+Oi4w
cAIHtP5wyGNnlun+j0DJfYYl+1tJ9aVaFL9SqvmMJnYMU0OHmtBzrc/2qadWgkNwqgMFSvcZ/tEC
RlQB/B5ZNyMuqA40A3+Rw01152QJH+z8PJ2VlO1I9TXhoxn9a3kxNqyHEqzbmK2u96TVku0egY10
+221WCuj3H7QCOQVuuZQZ6G7Y8q94DXZHqq7ndXotz+5/QaFk7Uw9Wy/fEyWOHIhWpbwMwh0NaU+
aTpwJ51wnMVxDQGVSQ6Wq008m1lCzxqmNsjcBWcdZiibZUnkWyUD0QfsSDhotlovvf3BVpdZpytS
/vpMBDkxYu6lyvihi2mG/8SpZMrI+GxVUtnvoAVc+v+YNYG+Rn5ZxKTFfADuy4bpJBdanu6INojN
yYqbFqGGiae8QvUE68GEeM5c/nmq33vmA4FJ1fijhrj7E8CbHduVbLaAs2yX+3fEruLjRtNGAnQ0
kq/ybNxfCUTcQLc3TWxs86p1G4qSWWTLyHFM9rVkU7PMBvEZ4sKMnPoRU9Z8BVs+tWRhX3g9uBxQ
SFxW+swrdyKlEbrJ9F7s2Qv/g57BBiMfANkziX91YZRmq7N3vZtrDsUBmEoV8Rgi4Z21Cozd1g8r
HzitXXAhUFo/BNfIrLcukSzlRZ9nu7t1Rr7lKY1PsWGevntdEZujX314rhHEUIXYPzLnqq3zaRJn
idif+6xSnFprMgQAMHpGTd1QZ+7Kf9ES03N9Tugk2uXXKh1GOLlxe7u1PRkVPBp4CJ5IfsOwYysL
FYcr72RRNMyBgkLd4Fu9o21POYiY2ZGkWb/yJ+FWFmns7T3zZSSXmefNBpkUT8PooFbEhWPOqpUw
wsup0ABW/YkTLV7mrWzZpX+V3gtpC9UWxn0gyZChrMn107DyYB6SC5k+jfSPXjJCpxSOdBoZ7X8Y
Brb4TRKPlGXx2rD/L1+EAD7qHp8sBryI6IvSbjqXL6x+cScVdbgMNMyn5n0NFt1WWN7VT0l1E11N
Zp0CKiL5lqe6HYU9knzA4w4/WETSxT/QjpfZSTOVAOxXrWgsumlfMsttlowRdwuL7flLOtxAmrWL
zY1auS63QG+SabKrByEizOHYF9IVxr/ywdhtvqNYwsF6GrVca79sjMBKZWzFFoAs9GmcRisH/dO8
YThFLSY722CgyJGNqhVaqh+1yVMzWcsefjtMLiJVuBJm5Y4qMxeYiu+C0L65q2ohpO8oPQ930FNZ
oGnIFRueAl0WnVaGUxws/bhJK4tJdtVpmjGtNRMH+43X4u1Aa72Ir2o6utsHBgayg8XyyFMzJqpb
DXcYEbSVwAnlmT4zYICgahPSuzuZdn0kskrt+Wl865xlAKmki/2tAx9wrkDIbt+hI+HihFPkgbZ5
adFrHcpGD2r1vzLbz5r494jYrCGXJEwiSAxrqlQqqhjc9U5YtX2gc11C+ido+WGDyD2tGe9iUdGz
vH7Nf8dfyd8H9rh1EZSx31B7whBnL4ETNxYgsSz8XFfoVyq1t4nT6D0PRNV82BN9fW7WPjqAMkAK
ni12u6OpUV37YAPzqtaX21oEWH+KqWB8Lqqt0/efQs74MdtfggYK23hVcnLTA8eoc16D5iS6RCRd
DNZTsrSSgp/UCw9lYSD3t2w0WsSuLtHpPf3ACb7FJpldB5/CjAPEh8AfbvdwoTlf5KgEveuYqnZA
rIhtni/6eTU/R6P6Rq3QeuL+7gfX+x9opCjxZs+w0U693Tpi8Gx/+mGmzUqCV5zQMa+i9X3tente
7YG944SICYhqN+0uxfuukloEIpblb5KpgfNSEHEBVXpIqQRrVNjVmFaCS6qrFpFTrRqMmApa5mNt
34/qmgc8l5xeqr05Od2CoRZJvHA3LNneDXCzc0NL3H3erMtQart0Y4Dp1Gz058JibZzo9vnNFra9
BCLWl1zWzaSTTR7JXcv/vY0aXmMkRLUzJx5Qsl9fcDGvIRxsu/h2sfdsxWNTJRDfAV8hJGoXVu8C
P1g9/SKgmDFyu4PS+neC44SoVf2Y3J+jKcWLjEG66xCkGedX0m1Qz0P1427OXp2uxoDj9OUYMsA9
8cDpGcJoCLNOEHryCaAXY4+HL5yFK3lXcHI0FHV1YZx30Jf16DkEwKNjvWVDSJ/ZgvRXzYH+TTH6
E5fO0+T7cVq2JQN/ylwLMIgFjQ7F3GBsTZAbujD6818/DJSrcjnSoDHEFuaPC/EzY6Kscoupl8kr
V2xil+GeLII5nVarYUADnNQ/MCgGftfPyR/NZIS+U10y4bDr4hh0IpOjaK2FnxlBdy+HRSp7KBbZ
dtB8xAGPAlYB7z3u1/lOUL1lXRkL6gHIYoge/CGe72KScwY2ii+Hy78/iMUJozuXw4N+mC3k6UeV
yRE6baRkf6Q3xMWi7lzi4Z00vV7cc7rWAOsHSUqbojPE8A8QGgRQVmorfE6dHg+VcNAV4Bm/AaAc
uTLmsGdO+z/99gVL7i0I01cf5XUeW4YjbArEec0eA8haSb3QSLaSioWyr515OZxNnNna/ITyRpsq
Iyg0oOlr+9AdSFaj53vOZODkhqZ+GPTeM9ifj57yyvfLvqVGfcFUCvyA/XOPnlGDfiRlwj+UPr/D
pBnrD7EKlDQu5BqbPc+aYry9vyICEie1YRVeDhdU4V3t6Q51yZjD/nVX1itQtANezpwz79058AUm
d3cPPpzvHDkeYoJAJ1CJZTkI07yMQIu34sXu2Ce7hnP2RbOdgdko7WsSuP7X9eCGTl+XZsLWcc+F
BpU+XozpsUUCZOAajafK4PvP8HPSlFJFtRowev+5tKFH2dQ7YuWMz8Bzq+Xyh+x4GgwAJj5vdQQS
JFtVAmgApw0ATgOZ1DVFLFDsM5GyhkmDxWtKYDcdngTm/jvFp+oSdRxPUYdpA/qdPM9GOwvyv6XN
c6R/qdg7FPjb8/iSiL25xX7Hq/z8RYZj0E/li849ses1PapHBFTJmQcr2rMb6xJOuHqiML7DvDD3
YSGwMZNotrcCFA6FQhV9ZWAWqk7OagidTHWG/3pfhCwLm2i21G2kEb1VPb54CS2HxOxHQbnJsGWW
4cSsBzk6TY8ZEAsS+eCPf54ThpnUDwfxpv9UEWnfAS9xu+D/fuhlz0eaCRqMDK4qdwGcIrh300CF
Bh/NljFr1RPL7dbzd1EX1P5OQiBFnlqDohkMEUpwEJuoekueIjC7FbvEY5JITpfCRO/FvjWk+d5R
CGhPO2n7F6XFYNobS+Z8v1GZwPNulOZyR5wbCmoKYAuyVCtI+3HLPiDuLS2NTtZWGrOUz2wx/6/A
C6Dbkik48Ue5GCviMmxoqo+6tXmHqYoKnnFe40hMWzXhxCW9lXern5A5QSkxXOc8va8XFS+A9WEs
SbHpzQRck7hA/1nb2JmlFh/RvOqOvisH9qgv9hnVjnm/m/N3rva2WwIWaVV2OiZal2tFdBOlzcZH
BJhmdIH9ixJ1GvpauXB8OG5ftwIGHeheRkIZdDchxLix/B3P7S0+1mqo1Tq5rf+10VwZgcs2om0m
53e4B5WCekgIOWfyJeptUtUYJfUBAQCgz9E/py12ZW7a+EtFVGrYkB9Mba1GM9AtMl73RUykxPuf
zMzIIOxJ7Z2ejLd0ql8VH0JfpFsZddiBu490wReNPq2vjLXXt+9eQ6lhiVX9iCG4/zeyZBFfQlm+
zzSjJkoMgIj8IabXkggABaI3939dNIU6dbwmApSi2radC9RCPeerzK8s7Oj9EtsoCgnY+Dh80J1V
ApXawBsE5NTq+N2EDCHfVyUhQwQyVYCzGDyzQq37998u1Jqw70IQN4PZbTMPDYbFT2vQTW5wZQeH
B+k3jcXlCEixoKBy3FNyQW7JmXpzcr3AbLfE05dHqwuZLPcmFpAakHCvfU3UKhTQPK9otZy6rCiU
EePXQhVfToo5rWtezRFs2uQTrBvtIQQ+ybQxXHvSjSJ/9uv62v7fYLKJXbsBm+22CpsSaHbkYID+
zhWD9p2S7QTylWzo89ArTG78/bGokvUqS3KmJegO108dg0zORYdbVG4RilFq1KqICAMaoOl2balf
tYhPgVu7NW790rLNSJkhw0BQs478MR54avcFaNyMe88qtkzLBroOhUD65W9uTmSqzo1MXFw4/NQC
wlxIDCGlEb2dYHEQ/TnyMonLmHoXQrQPX8Ev7Q1V1Bbl4B/lsv0N5M5O6KJ1ktAQZyfn1tB5Q/NG
Z1+lbw77uPMkyBjn5fdKAH4xiPTi4IJZf8TiwxBOrewDvcab3mdh359o8nIIceoI2KZbcwl/ZcJ7
K7x6j70IszozrFPTNbGG+c3ROKdjhL7gUKPL00r2kP2N7wb2jHOEZYOGndOMBAUD0JXbIBJqD1jj
N3yAehBec8an1ULO6kzqDuZk/KlD4quwz9qEh6lPxo6ggBcgSt98gs+VGjMyz9yxVgzEaA4nc7ZF
LbVG5oko6uDlMpwreF41o1GLla5mfw0X1c7cU6J1Z42/md99iFJq9WGIRDGXy3r0LwO9ScSLLtzD
f2wCsV5xCctdLM3onAa9dN33bJwJi68F4Il4yCt+5twwXXFmRuJlv9EDxS/ubyDYZKBs5z04eG3r
wzR1EI5Qd+cmX7CE68zBb6HLrR+ZfTOQckEnlDgXsW/I5QZnG8+69KYtm03ietswPszeFwmSVHvc
XOQth1Im8c4EAf9blelP2fQWMkTCpl6VxvwHr8A6xxwfUoldqaHiK3Oilbg9Akft4VjuokWyoK3P
k31dzFpvKFh35/GcOnjyUcGs1ZIy8JiyMInZ7BCtZXC8a98T2ILhbuu2z8fXDozIm3h5yUXGZ5K/
ftH8fgOSyPHJTuUalDph84A7ni/ecJF0StnWoE4JANNREtnzVvheGh86Y3ecnkxqGTZJIgUzPZt8
MyZNlJvd5Gd+SwFg6Q6afdPryYz0fVz3NiYw22HpUcOohjb5dgdIEBSahyZ4OQZJNJJhSt+s0vuK
gsXz2JsYx4nUZy0LJ3M5B4skkF4d0A1evzZprMukZE3G5WzvP7swpP2p/YgngrSPrt5Gsr4NuvKE
fF4+0w6r3wN/9hIhvnPJvYJkLnCRCpf1doBrO/TDLDePdAHnn2FWThil4RAfsNJnGhXjQwZTL4Br
xmJoOPr8g1wXUFYOxs7eGPR30o53MFVRQEXRQj45PynMjF6+l67pNM5zQpUq/ftTSqecsoRL1QxO
GHUt8M3yj6laj6brypR8x0nN4y97/3kkopSWhYE0m+hbmPKwaMekVRAeQia7S1NqohlwFsIzxsJy
c2L3zw7OZxCwe50E1iPK1slaU4fcBoFZwI0+e3kehYrBsvhRCgBvp/XNv5ka/yyXSLSXuVii7BiA
i+02V/s+qVi7qmsa9bir9UX8KmBQ4irSNLJe9bgnGBY7NxBftrAgs5mGHKmgDBjhnkhCobzNy8LV
6PlbmGrzkkgxn453LS1ma0auTSbPOeK6MGhv9/3zTZowqj5915yZz1+/XOlTHVu+iZb1AU8vSUhB
6oUBwIgWYEEsp4/PYGWHIZASCkwM34U02tp/T6J/eXQ47JxIo75YJ6rLL3bsIxTYLkL/nHZFQz4s
tC6vr9TIcQzG8gIiRP2B/FxTQf9U2MD2cn8+9g0jMay2T6RmzF3N9dIC7NT9WwMiZhJ7cszHjR9q
eVFj4+6DQkSMLIs+MZk2VsZRe38efa+4Bt15u7f2Mbsi61RpHlDrtzCrsUFncQRWo8s/zB46AWNI
9QAnVWx3Kx2ycZkT2u61BaO6XCI7xwOKYmhZMKHWV6py/v8Kv46NmaPlM5gb1M0K0D9JCCfdzX9g
2ja4n8yzEKmlt5y4eHiuqhGiCvXyZ8d/suqh4UD7HPfYD1L2MvOD1kQafqVqGmkXfmABMJGjhj4E
NyAtgnzV33aw6v6yoiQMXeYslO6o/SeTVQ1fy8NUNg/CpKAoLOQPu+kf3lb8yvPAxg8kYXNrPUfU
JQmpcBCrbePuljevQD0TOIZa67n7u0nMen8uOwbea56uLI6WjmG6ArnKnEKm9w5HACsKvPC2ehYi
qV89VgwkMWYN8KUi7EsxHPvxyQydoD+jsPVsbloroUhuyXo/QUNkrUs9QiigJumN2ZuczitmZhEU
rObf/ZmFQeDKGlJ+TS58OBqfNaUv/IOaAIlNoKYh//yf6YoNM3xZ4WQy5JGAfgmp83656qb05K8j
qCMGTcFGsWu7A8FRkG5uJ7HabXfRwIwcAqSGQxS2x8DyH4ZdwrOCKc3PDeaOsUQGMsAO362r0EfQ
1eHXEWBfRF2Mab81PBEgmFhCOMQ5Tcoq4zq3uocC2VHJmn0250UrQF070aNLXbYOCC3/rFYY6t9f
NZal/5GHVjRjnWlIUn3w5jw4n3QkWLGu5IdUhyEx9FH6xKsJ+x/iDH0HeA4LOZl7GRR9gL9LhPZ1
cSKzuCBHXxMZFEDHemc/SLuJHL1RknsIgt/2XPQCbVszv2udcbK5CeH2qfHkezU0W35wr+gwJJSK
QG30x7A5QIGjJ87bL56MI1Ap2lmaOAxtsnUIXS88/CCgPT/MB/732cej63J2F4igLXe0K1hmfT+M
MTQmUBi9u/q6jWnok0KsPQZnc220IpfFeDVxPDlu6tGIywggWf+z62Kw3RgdYkmtvRfvupCTJpN4
p/+RS13wYRITYNeZhpMN9lgtdJhObHp7CUNs+ryrC9hXqX7n4524HSJvxkevWtt79g9oWed2R3ez
6cY8Az/+ALJW4BLlV5G80eE27KLzUXFC8OFr68wFJF+Nfj9cD4cFgI+K/g657Pp6Fc/ijtH/Omze
ky1DG2bvDJlyPfMvZruZt+AOyMIdVUzKvvgV0wkqXi4Bjt63+KY6/9tOYB6e7K1R7MwLHZeQeZTO
YcfwOLJZGeu855KU9m3JIkibaZwoURA0YpXsujPWWZnCBxCz1HIG1cdxwAnMzVrD+V+VpQjMN2Cy
D2Akc5TBBu9+YxbxKZTrgkdLp2QQpZKZpk5aiT9H9NERsDxbU1t5KA6eB//AIfckSkTdFxFLvBlT
WiaC6WeYjU2T2ZJh+mestCyrvv9+0K5THi4Y8TfFSuc6NqDnctPtpIGN3L1J+zSM3KSl5ULRLR4c
ZoSAIWyouWap2plbf1KRrC2rSg3H9ajYUkjj31EfcvutX/pNyCDifu7/8W2j4yGqgZD44WsX3aui
UZde2xZyjdQ2Dy3BCK1kakasXhhfjh6o3yKdS8o5CUlO4dDkqmwsyH8Np3NOQSRNXxSiB8f7ajkn
+nbskfKPoUpgB1h+bdV+F4vhmkhAYFxQ8I9ZjTjwBopnGsfX8TpG5Z/yZhqANzZ0SOENZel1uTwd
qMagYVgiRliwmhgositX6eAZJdpOj9rbAkUecXYkA4vwOVzZr/bUwIyQ3ClVj6NUOQOkfroYb57j
jwp19s0XqjBaPxeEKY9tCq6v0uJizjlG8CNsKlUPKkydKhv8m2g6xM5drlT1PkAul9wqx8DUVKxZ
NLSByb9O2yXxLkFfgZ2VJK49iZxdln90iTHZ3iDylNjdIw+jwbXDdw1RA+jdV3GacwpkHBTxjOpD
/Rbfd7RYlQmKXQBe4+Rn4PoNtDIrojwX/U2cGR11muUKf0yVE3jDaD267eoFmsKWB7nk9kslz4Px
m46/ADs3swQNd1agswbSjjHr+/CS63SAfhwDJqqOLTenx/VBZJWug9eIDo/bxVfRmlyhiY7L5Cpy
Pqu/Mjca+b4A67f6ufO+8IPONTUGXtPsXgXy4EbpSOJ2JK7W0kbwCMHocri39k0uLVW/SrZsw/Rs
mPEXz+AC8qvGLNeuhgVqLH9MmxfICA4tXpMlks+W+NuijQkUwr3e/unLYgr3PkYwozibplTQAvD1
IGQaJ6WO7oA/SAVQjoHdtGL6zPVwWmxCV0j1WsJkDmyB99TAhYGJ7c5I45yWeQkZDF03z+SbpcMx
fIyLk4jkrEMZl4pWadAXjvsTeo0wfZBlFjYYHwmSmbxlhHe32RJZSjZEtUIatwAEhVM/5sDPGUMC
98gIXvvQGRAddGwAyf02wgJR69rA2FwQwUglip04BvV5CE9SNoFZnH55+jKnnG6diFlD6yfyX9rv
hUi/uWhmv6Evk+6y/442HLwRUkCEtkA2oh1Ko5yHxY/Js4ciKYo9x09Luaz3GgnB4LSaftAYWyc4
H3p8zYge6X9mmnGbyRVsSGPQhxidLfBzn5C4Ufl3r4bPMjewJSNBautFjJG4HVUppvguHeUXXlWv
okWypfSRLmOeWDw+VU5VQ3xlgP0a/3tMOHuWRuu7RVWrXVEzKHgUCRV/f7ynBpeZ//Zjp0Z05O8y
4gBgZLkjd12gvnlccK2+CpaNqq6NczD1FsPZSs1/rkalwvw39eUMylQbv7D7H7NgXYpmjvwcmJpl
FyQdwi0Ks6CTLuCJtCJQMMUh0RgJooLCHW8cox7RkCtEB5qje7PEwi/QFqHyjbYUQCqyr7ipohRq
UPKAsa/oNKZfXfE3kkIO3znnf3G80kO8oR1pDmTKYLT6YpW7kBZho8+YqA311gcqqKgUtEn8n2an
E76n3dmf3V6WI0T+ZX2LcxG4PR6UUfl6LsgP4Od6dDYeLfHi0dSCrUarzVx+zHttJqSEduw3wiEq
94a1b167DyYXnWnrsxeX+WYAmAZqfy3wRqVRV3KOXl/6iwk3Y8YNjxRBppOtmiMVNQnJATMdUhKF
Ym7K1iJQbrRE2m3HGg/Y/5IwVakDwXq3YReNJXv9eouBQjrk7m66s2X8M++Zgiw4RbSB2xdbCHIE
hzNX/e4GPhngpyEGDCusSaiTXG921fxEJQ0QFFz6SMUe1F7aSSHf2p489mqDQikef0+5rSZVwufe
SMtsU3aoIQ/LskG3oBuClCHUnc3OS8mMKZd5w0QvAWH0Uqxh49dUJ12m42xDpu4xZE68NED7YvE3
d5Atu+jjdtKpEZh7eyYYT0mTndt7XqOlKNNCWlMr38B/fc4QaNu7sVtKBc/X89MxfFOoekSs9Kk+
djkPSgx2Zx7/ZDF9T/D4zF+jbY2cum5tPlAAmOqAB1Zz/LcTSSi1EpC2qiy1eKP1hhr08YEAkz5z
8r4JEqFAlPROZcdc09bWsw4uSRyf+D5ejLVIm2R8QFS352lq/o8yLqGczt6O+UZGPIlAaCqsNLKN
+8kleMwUF1FhJmTVzAexx4ug6nbc5fcyLNJyP8LyCIYKy9nSAq0FAXXw/EzS6pTqhy+vKaFEV9Nw
jifWuHMc8gL9J3nnz/bzwnYj4ciwDm/67ELT3239vVB+iIU+j8nY3GjhMBps5Tfjjubwan1gQ2m3
BGIo9QRyVF77A6OtZhW7uWEAUWGIZ2prv8dlMeIfwi5DCcGywT4LtOlKO3biw2kk+Qx/7OFRbhHF
auTYrKLUGrKW3V+H5fhSvPWyx7XNAjgMWCmegSgNIjsg5/ckpCkOiWExX9TKcOIePaG+ORhWLouE
h1KIIysOW/5k/b3O4jS7d/tP/LXidyRwMnR3k3aAwlN2z//KdYEg/GZHeApLYA+UCsygV/9n5ekw
WGW7ORZ4BQfik/ztiqHgKIGLxSFDohcXHffUClgVJkBL8W3CIjpFJrLcAoRd3Hg6YtWCA+H511ZP
Zych71i4ALLQ5BTBuGlzgO7xbpxtT69+qihzQnX6FX2Dbma6ogD5uKLy2VIJD3PFJXsy0mQbiRJ8
IJhjZc+Nc7gRMoXXLr6jmh+k7Dmv1YemMOl6eXOF0+o2q3uE89eGJ5PJA9ltl0+iMsWhw3JVgc2z
mAby2st1yHalq4B3Urc6z3/tRWqi+vKqraZ/29TF8FvqCcGcB9MHUxX+6kxy8ONwkpDto8MZvqcM
9Jfe2BdHkVxO170HW8tfQi0Rm4wwmDHL0dp3qsAGCvhFRhvkcz+X8HU5UUGMjaWiaMwP6zuLMZbj
NnOz1NG0K1Y2Uocv3sA0RCwKxfaFUNYgCOrLXJKDawY8wS7i7Ckr5OC0YNFkZr7pk49PReSEexa8
W3OgZNX0+EU3iHTMOoQLrAvvq7UCqtVwU7WFtpVUA6ROciGHA+a427SAVR/QqD2pkVY2+++vkLDy
ZX/jt65ZIDaf5Y/SEJH15uvxp4nGUmhlUbj8R3v7mktKewXV1hFuNhvy2nkSQK7k5HvrlLrGr6sf
cXwINajiBbVdn7LNawo2E5WW2/W7megZtYTt7bOi4G8QPd492rpA0y6fOEZ0Razghlx96UuSl8+t
9AhyW6b6u0Hxt3aaw+wKmsIZ1c4xA/i6Xd7Bl1mJz3LTAWS6CSlnca5NGGjq7AZfxmbipA1SHae2
5w3nHJWmIhZlGpSgfY1SzZ4/MXQiIf2wtQlmhp3klPV1Eza9Xje/kI7Myt4pdPWWTFrPD4f3tMsJ
SRUwV6lLRRP0yYI+QgJH1oJ3zfcW+RWTahjAVdGZ25FRx/M3Xb6YMkMK2f3wsT6ZMnd8ix0Zpijm
acXiJ8x1RR5BT3crsYY0AxUM6QYeUS3uCjVR5eIvq010HxmlzJyA8kOqbH2b2DwT50AbCV2DVlT0
hX+Z47H4/9iZCiPyvUvF2LM7u4l7IA2pzWr5pzsHHHRe+rRUNeA1D24OwJskLGmlKBoH/zdGe6pC
IWi6Y9K1E06NEX9gX1HW51IwY+J9EEERxsCWnjPZwsqC3M64dx5urmJHNktUfD4Me8CqZewgUvTs
2IX2/U5CwBw54t+T2aukxwU/4Wi9FnIrZwK/yaRFpK+7TKsnq5ju/+hA00y6Yfjt48piJiOi7MmA
doRqsvcd0CfysfBRizqOJTUmtg3JmACReD05kBd/+Znt+T9g/HLcmSJabAiSGFMPDVEn+cIcr8HK
0fP0R4MYwSH8y27wljqp7HMl6NfeK2ccqyqpq8ymm6VqlbQNyKogfmT9i03oF5mKTp2TN8OC4c30
273aNB4Pur4gYeUz8gvIC8yVngLDF59uFFaAsa61E0rRYCH8Hai0+YAealG9gJFEMPHEjmyMH1Dv
8nOICIsZ3A3LcnIaU9GdSXlcfX5e6IPRoGpDhakM4NZi4HCfRT2huc4qMhlGjteRFHKJAOPfk9yv
90I1CASAASZjOl1KbrsG2qiJD2dFQyOnUxIQQj/qivAO8DgawZ/Z4ZCBQfmoSNgudQ7RBcEafUY5
qFUtqConk9ypWziQiryJzN/kROU/FqiE9NnF2g+QghVdfmprHp5RHs6mHq55G5vSEIKom7Gu7TuI
GVPhgjnVbcyqlCCLD1vGxSMdkk3irgcT9yf95fdx5QsRCVcY4oMPAkdeIdFl1Ai7mzSf0JPK3NaD
5jJ0PAZfWO+SjSIKjaRhQksJIreqvCQZ0WN973MP9k+tZpneNLN2ykl4MLXQVq1L7qqwy0DBvA2T
cLze8QwfJav7rkSUSxNvzj4XkQY9sXGgBa2p/NamonphW2Sm1cMzJNrgz2yBUchYj99iff9pW02Y
twNrfNeAyh5cylO4vP2RcWkNop53wddsdZ/YevlRnakVN1yUpeF5htXSNKwucHC4qfOjx0Gg/YA7
/JsqTlpxRppDJrunkDS/TC6qV+nfFYxQE5sH+IzQN5P/5JH+EtNKYrbSGULbVz9fFgnBvQxn7zMb
GmNzH6GMhH6coKYa6bPw/AmTM0TLwExPVFKUR/Epwfvh2SqLWJBOTXdcvWC/Kr96js11NSyjgSWq
Q3pS1Fph98YpqJ5cczi1JfXBpiQZ2Z/v6TzkB8AvztAbySYQ3Fgi+ZQ0VU+u8rduKJxYldE4Rq/q
yW+5hMZnQcvPkfq3lEmQluv9mQdnRrshi7rrJbX/YWdJqve5WdMdsEQ7VpRoxVpG8Bbl8pESRP7i
8vsBZh+/cXtIvBMDR2tLWSDY18q8BJgEi3F78q3P04wdjK7+OXZb9WrStPX4G9yqOAW1zPwEDq8Z
mytCYEYkVFz2zpFNdT4YfVaBYAX4o8Jwa7p1S6Yf7rkAS9vOnImp8nCvSHiYBMBCCnbWSSeKA6Lb
qfRDXZ9km5MSKaTzyNvBLUA1A/aqneJpFPh173NzVfrKS3+R6lkBj9RYMs6hfUr22rO1lKBBqOT/
jwIDLt3xQICus3nj0k3LnSahH8ABk3gmO6rxB6wAbWjCJs3wwFIKZO+9dn+UMVjQpkM4DADllVj+
0zXEENRt4V70gUvKsPB78ybreNnBBxJzIT5u4y7/HaPNu8oJkihM0YnKFBdtsmyTarEHqaWIaKuM
sM0KRLo0F9/WV0MHpTa1WmBzToIpyqZS5jnMLfgagNl7STRsx4fiBJZdvAwE5+S2lVLFsPPnss0I
WqZPGeeT1dfdSsNzZzPCFF/vlf+kcpuYfaRVEor0H3LKDoodN1QS0E+VGwQKZHSHtpbAIgk/qiLG
+V7gu65v+PaWHfkUSGJnT6LqNHsowU9ovPn5o6yFCGaeiIB8alynHBOZX7SPINqaOCOQXazy2o6L
Yz87Rt4vy4Jf6iAQSQ+2KOnKxtBrgpoEhr9Cz8GUjukGovwjKUPx7XTW3hgB32dIMQbLROcZx8kW
hrHj9/d/VFcYZWfkc/mhdA9qy0jOd9I9/G6YYCIRmMDs8+sNu2w8F9A2Mto06wTc8hTEYywUX2me
03kiuMsZmoU6WrQFFrpx+IqX0rXfppFWqkmW1Sf1Y6Vgxt63nI0bhnDeOeR4m0FKM0zt5eWkyu5f
8KaqIuvETyD3+b09Kn5CRcqBrqinxxR/PU7JxxKfZqjqeKShTpBDT1wOFcOE9vjDloCWOdGLXb9j
sImn986TG6vrog/JGnEkEyq+41CHbyBxMUh1+LPA+HtZJy2Dzw7f0BdRezmNi7s5/HzrfajKU2yS
8Y6hW5LMecqQYEKnHwsTVCmnjyxfTE9FxeytBSSYIH2qC0ZOlOk4cQmye9zxFtoZBJxTchkjWKb2
sflo/yWBBnqbAcdZxWg6eJfZnOcgiWfGqM4WrA5QaS/AIjnGYWPfRrVWsLZvk5PvC3XyueW1wAmZ
UQOXNT8/s2Yi1oOG9NGVZxS5BDDg9BPL/wf4mFlZ0eKd8ScJiavYsyjuZmXndlN+U8LwPu/m79Kq
Asu9dtqv/VI1Ss3K8R9SsCxXZJJwM6eEN7pAWkWGZhLjkgLY9vrnLIkUuYMV7m+3OSv8Fnz/uGw1
nVYrEMtQovBAz3iVgFWWmdmIxOYFPnJYHlodkjwdE8V12ZVm146E71lqxTcT+SjHN72j0j0lT3p6
RPp5xytpR+3d5VNsMmlk8c1qdekzIpA0TdUaCAWrMcA3mQebU2H7WBfwo/4m+tLl/4FsPknE1aOY
ocKKCszqUkI3NSfsV8Az0frcnw6fwCx1EKbIRPgMsj69s7u8oJ0NMxq0QxhjU6dDIT+U7vwNwoJa
x/51+sY9QGKeTlWf7zksTRKYVgRcZV5/2FBg1bsRdH3DDBMmkHc+v63dRSdAmWErmcR+4zaxD16H
arncsyJFbGkPWFgCic0iwHX9PVjaj02xDSvOOfzv5kT7JNLN8yXi4oXZdKYZiWlFjAm3zRHxTKUP
s42TeDAhZOqIj4Zz0RG8DM1e6lQY36QVDVeo9nPTswyskKyI/lf6VMUkQbSjWiBFTw/OQx3Zl1p2
qUK5AzDedv/9HLRCZY68tUReR+PszWSv58p4F6q8RnMzdHEVIPqTWWsPp8/Z0I66Enc69a7T4dZm
KQimsKNSp0ksfuqlPWpPEw4zXU30fZRCMftjmEMZVz9Dt8o16+pcTbky0ea9p0TPQqeXKFvaysbJ
0wL98VVcRRUD2aZ0YYxsgKgtLlNz8eSLkFWyTepjMviXfWjnZosUXoOPGKCWrQp341r0hiHALTU0
KySPzVP+ZqwJbrHwyu6Vf44I7ugPY1A6sKpoOk1sr1j5yDXCFWNpvyVd0NIWk76AypEjOHQItWO+
dK+5xBd3c19R1T7QFfsdiZDGbR3I9lJFDITW5R4vw/LBiux0O7giDoNYdJYTirN2HGwsO+49CPdF
AyXhSwAgBHf3cBre26k0YCkAadS3AmmYPAerUDuUnPy2wGsGVDr1EPmSnTtoU8O9MR8ENB4f0SUk
59E8ZodRalyhI0OcY+PUxaIomzmz44N3C7B1GcT85LUzMiL+ymd/eJmbEWYtp3IlxwfA8xk1m7lK
lRSfkTDHu1ny1IleT581U8eyJdiniNVxYkauy0q4zNxmJDqicZSeGDQ0X2VGlHabpb0I0L8F2LGn
GqxpDazk/nZzL5WjKqDPOKTQVioV1fM3+sBuD5ISz1V9UAp0dOzLBCjLDJFvITiRjtefP5py34g9
ZFe29qXHGx91vHbngaIhdh+ZYHCssbbG8+onhzuP6jlDCtrF70zK/NiJ3rX50o+rx34zVZSiSH2C
BhBvM9cOmQhB1EMeJ1aa9soQ+t+X09cUtmi5YqvCtkPpNXQDaGWdvUEHPekcSXUGmCAi2Y+8UOcG
aVnCoRvnDYRY0Pc+I7UALLhfWX3zKh07HU61lmH+7Vkg5PriXb/4REHTT0od47hAHANYytdYF/pK
Cf3k6+B5Z9IWZtlTwmJjxywecE6yPYJ3J/nvFt05THeXygWnFF39OcDc3XYoclr05mXxqIW3ObN3
kOisstnzYGvZs6+yxyiuHfvA5CLPJvIBNBOYIYu9FcEyIIIo+A6eJRgaIJSMSBm8jXgwlZv5y2p8
ob8iBxA1HS6oYPk8iyTBdHab4+DgppDcSDwk0UeZZ/UW0LWF7fo+d11O7Pmls3Z4UF6hwdFXpNFt
HC4kvlXI0yaGpQEDFjOIP/pMm5NfvStwAzdIKfiQIt0eM4ChO4rVjPV86VsnjIIpWAykJIVEal3f
sw13pp0epwo9eVvhXnV+MyaFAJ/e3vsjUcd7tTZQk1HUXBy/CJhna49+F23eKfCphscp9tc6Jqxi
MWf1dTRzD9pDuUOhIiBt+pDDvy5Uv9+kWBNFo1W2sUnpdax/9h4PJIVuClwKCAo8tO9LOLWZQ7+u
K11Cfi+nGGPO8tj9g4nSAZqfXt5u6FYXy3ckzekbQwoByIq5tV51F7Jw7qMxTxJUJnVDw4ipcEby
PpeKFhAeQoI73bkKlRNBTXTTmh5zXmchjjWVc4fY9uaqwQvuyHuwAeRzuKswbKcfBqn22QQnJgap
PkFjmkyIgbP7g9sJZqVKq7irD8jRYumpSp/0dXdFvEkro3XTfyNbtYDSoCH6k5sTEwPLJtechGLV
cFfrYBawaDczAbE9PI/STFph/6ptlTDoB6E/CPZ+w58Jppm1zrO2pu6xLHrCRUqGoA/HdH83tgiL
AeqKvVZbC17uht2s96UmTvFEvYaGg8OgMV6qA+URg37TQ74fxIZlBKdjCI71F9TAHLSrvfrsFZu2
tQ+Db7Xb4hs3+705bYkiN8fW0HAJOHNgBLIGVzzXmWlwLifowYJHJtG+0CSJWW3J+cZxnE0BmWYc
yvuYSYvd4eeMdR1LwXE3jIz0ddRHlyZEUoXvXwrZ6VKVN5/uvHocNIR9vcfV0NPXH+Kulmn/v6Jx
FCzylJK/HyXZXSZ9W4/j1m1RwRiD0FNqVt2taFbQXLuP3tgTmmrqjgm9WmcOgeY6qTsbohJ+KDWE
8v35uir9F7MaDWkLYuRr14nKfTM3NLd5ylVGVDXVp/vXB6eoxh8AA/0Z8CGnHk2yY1VQ0bmS/cyE
m44Kec6exuIc3BZn5AVFZgl/FYlX6mkB1tBQ+HgI3Fs5cMOnFj+rSQTujmD5GFko1nRoVAo9iyvz
OGkZ0e/x8uhsc7mf0kSvGUa9vsqfMlzNx6EhlDv/qHtDV3YKx6IE6M31drMQs+lf/89rrEaOBa7K
fhfIwLoXyamQorYOKF/aAztH7Jgr9b2ypso0AZ/gpoe/XP2S/9J/n7bW3NQz4QPGJ3MtvI2X89Ch
7cnYFZyAhZHam44vnHHFNi1FT34B5/4FVPtnlr/l4SLak9TE1AOz1OtMPi1DRtm9oYbvWutbkg30
PwByivTLBoCBDB05G+8iH2sCmMEmwWt8tob+RKSzO7hFhE+OgnGbK9gkcEwygqprp4l21DzafAOh
xdlGFBEhW+kBpvDxHXZdrLT6YRB2fAKqGSPptRNAq8KvpZYzhJurQAl3MvWVS7TkFfZ6ozgxAwrn
XcYKNoYIrI1MXD87fP0Ibub3qPxh/gphq7WT1MeTLlbKkdkr3OpLo+4vxkFIWpEPKtc0wOG/FTzr
0ERMdc3Q73o9S/EWrB1D9dJwrCX+DqpYiwxb2Yrt7ZHHvCx4YYhyqfRCZGtXq4pXsbaOnDC6OmHb
AE7RxSZUNvYC21hX6EU8g7e6DE3e8NItgJFrG6P32sleu5DkIutKbZm+viHko1D5cRvAGQVbTb09
cWRyt9wViJjpTdET7sGb0ruZhSpdJ6VQmrGoULVCJUR3jCuSC5q5CixhbaokaHF9t21N4gnGU94R
rs3TH+UzgqG1DZXo8tuq+ivJzU001QbyrVGkQTpnSX0YJgc224OkxjrcI9zdPZ4P9wGk2/IwCAm3
M6pM2XmsR3YE+/qof25Lfnz8R7CwMzTRlfJViw1q6bGTNnlrK085MAa+NQ2Lvpa8LgIZ82+gQcry
MeDXYhvMFEtYreod1z2BjWDLUXkcYyvcDnXAT9yd/chrqzEPr+GG4dkEPJHTq4m1tmuc+ClYDiJX
daeFuYw1SFCHyKWib0sG/mQcvmpFt2pWMb7U+nFaTQ7Zj+iLy254dhypIDKIaMAbv9ODfAY+kZe+
YNnghpzW6YVy8G77ViuQbJ6B+7VUxCkkn0N7Zrt8of1DHk2Itawh2WV9oKFysM0QY6D6Zbbsuvtu
en7uiwvwBlYmC1EF2pU/xpui3Nme7s6HbYJP9fY8/8CENZd2WTX56DaLfoMSQ1FAKvRhvBoJ9jYE
C909eEpoGdsV2+d9R44VLnBjwxuwmzELbGlreI5j6JJQwLFwGTnkY3zUt3MPJNfqXzxDbcGKHrkx
fiwjNOBKFaluWtM21rqxZLC3uvrtNmm2WeAz9KKVyLBXkF1aUmUy2meWzXnb6PwlELcVV/DKAqEq
dSZQjdtfV6d2JT+enoN4lfOeA8LC2LrrcSIUPmm00eNnSPVaYyPXUjs0v18XZyjtVHjhn4SIXiYt
SLQs/j6164TTybMzb40WD2xjxhVrBWd/WjK53YbxsN1GYBFunRpt6Pc2ow8tK++CRwzpHjey+uq8
1gQaxtBeXRzN3i0KAkIUFT0loijK/L74YTm8+X5RM2VGBKs/oqUgTT7E+Eam2N2L4wHNdZpXhZZ/
/dU8ptHgieo98FjgBKAqBJ5YXHu0MgdMtFVXjsugENAMOOGM1EgwYoN0yZwlICkNCqDTOev4Kvf0
TIBH1CJS1zwzchkXHPFDc55cvCErVPDVg4TnshRSg0M6zqpmpji8uTe+eUpe/3D+7Cu6zTM8SgKR
4OMNkf/L3Y1Dpk1HWZmORfpaBQvLHHXflz+uQE8DE265X4av9yeqCyRe754qpHv2Xae3e2FWMnob
aMYRqr43BdDETe9CCHujHxcYmy+4ED+hApXb6Z8syNikcamq86o34kwRVr0+o3EIFz07dDvdEbNh
SRkRi9iza2dwa/+2VejDVbdCVX1mB3yriYdSty/Q67xwY91KohVVyAb5980ND5Zu+x5CxJfdzGrw
SZCtmrmr2QbawSF35Ogwv3PzThIfzPJrqTYWcH+GupCPVZe/zBiOauwPTkQ/aEJHIskd6Djv5b4X
OsLTl8mMMoc8u7WDhQqGTKuVvm9iEt/FMZO+cjLH0KPwbV/0TW9wdx7W/yHyVgKpAdB2z2pOydVp
na7eyjMeFnn0sK8/JE2JOEDbeplzofpFFJ0a36tFEhdc7XgBApF9i3qf9AyIYeb6EVj1iIZ18M2A
8n8B65C2+QFaBVEEVCIPgecarQxbXuNMjMHlEpzt5wjRRzreqnuKxX+CvXoFD0jsMAo212sOp/R3
I5MiiHO8Au1rJlXJ+SdEtZ0peV4Oiwf7JeElkE4wcB0Bzwvo0oTIuH4K5VNVEcts3GoUFZBrw1tV
pkk6WmHHR2r803DepBsZ0u2q4AHY2BwSURh7pvTyD3NjHO0nFe/Vr5mpxiZ7InETI9aPnRKTqPfs
NbfR+741MpNrW1TuDeLU9qxQSjRjXcjKh1595AW+y2VxPZhgLNYBVjGD/NN/LEaOjpeYCKnnoGWV
TUtwOHvZnmWP6MzEKRHxif5GSxntkGhvolj5SCGz+oKzrJ+LajscOUYIkGR0vAHYm9Gkbl4TfX6y
GRRmB7Tu47y9GOMTN4EWivWtaHEO0F0f/971PCn1v+3HCpMOAp4j6RIfQUNHaa6MTBVDUOvi/Kg5
+8TLR7Hgq3g3t8TYsKktVQw9wcVhEh0MATdtzgq8mBQmHRYdirOENb8QI44oiAE/WVPsIs5IlccD
zobqMcT7pF5WDOVWN+SIVimE/pPXATmHg982hpxeciPDIH1U0c9Cdq6geHVIGZCm8KAHYJAwb9N5
l6RZKZDE0FUWfRdAEfHADd2plwmVthuZ/6NT7NyejWhm16ObliM7LY/SRZv9RZJifyItyr3B+IsB
RgKzzhESLWaHrGBua+RtQXDkHviXCY4r6ksV6oBKWQN9tU83dFfKdPTB5E8/mfsCWAgghfoIlqfY
o6P7+T+QKd9RscJO64yHoUh/TgRl2aGlYjHPSWPXiiF9wJG7Bnapcuk/G5GP2T8DcGne7I5NjTIy
NbeRk8jIxW/dLPRcdDk5sSmsdonrW6rXmfc7FU4O2YBWMGL5u1IkOdn52Kaz5pkJxJC6xlyTbzTv
c9b44+2gAmpJHuMPPdvV8C4Sz3jhEPC+0s+0BhzhvB+pgAOJ5Wub49Qum9OXbQKA9DgEoz2uwWFa
xzaLRy+N7xG0N1l+eQs68pH18DlUhN1rb3An/QRddynn4WQLB4CemoLOGNu9ZNEVjha2MtHhpwAB
tM7ih1WsIpbdJKacXDHqSZ3R+aaHyClNQgR5N+M3tGyaSGnMY3M2lhBR8Un3GNhVlRL6t4dXW6YH
60g95gMZlSwzW/P4RUK4zavnbHakPF0w2dJYIRXwxgXR3iZ184vPjerSi0/UfvJIpmW6SWMW8MKX
LLjBIc615SzFK53OKRcmUSQTQ2VbyJCgNe3SFe+tvOzODkG3QvP3XViHXnw/3VVBE4mtRvScmfGg
7BCvogzgnoWwa7qjxGWOe9sRenX427ZU/fK1oTgANgp5pcVU45SMCcnfpp93UFZIJZCLnVqb+rIM
IaaoGBKIOtCfZlRM3tyh5+2jCsDKKjv6oQmqRisoxI8QJncReRjZm5E9vrogwaoUqnmE7BSNy+7q
UjGyS6IJlZrIjKZnXwvd2EReL1o62nrDYTvCL2P6vNIv/Nck5FmsqwR5dtFL4Gy0UDa7l3Lfd/eT
UmpNrrqZpEZqp1HErEWm07FkwMFgDqWjwMyIxCIyrUtM7TEpOujDDV8y5B6IViXhkr6pDpdD5qu9
boeWsy7ooApJTIdqlsc76zA3LQvKFF1OIkHfQdZwRH06fc/b8sm1lyxMckmNYCVkVHbnsZ1z/4oN
CxCYuwToWY8Gae61x3WFUl+DQblo55b2avnRC1BrlQOApsKEEvLAV+3J0uR/l/0yKhps412VRMoS
YG9ZBoL/5ERBaYkbl62HF+2KhSIVPc+U9A8n4JKStlpJwo2NGGeZSKRVKd47CL2ZXTZdGNtOEIEx
/FDhfMg36RMidOmMSr5U2ieI8voqGVgGARsvn2m89zBZbKix/YpeAP2IHtFO/U9zFZdrvmyKuJyX
9CmUZMcbp63VvXpZc7Wv8JpR5WkVlA5G84NkcIwTiJf/ILd5TmO7xEHBUmoIG+807JTAWt+B2IBz
yfw6O+zVAaaTksR3KEvihDh8/sbpuCsqGjBMJW8vUV4h+7xq5X76JIOVo0JlrkTl8eWiuwgPMKaM
qwvvKHykSfv6cCUwDu2SekQ0xHXPxNWYbxoaW4pxw/h3Gqe48Z+mb9fIEh3cnHLNFs/0+L4LXcwx
4DBA+alyEfHut/isv8lWq53I7kQBQ1w19qRhl71DF0BSFoCBqcaEKSefH45qRkD645VraOcQprpI
C+JQB9YEF+wGU1MNb5509FphDbgMP2eD5PX7eKgm3/F2wWdrbJZVFdoPnfkV12NqLR1TH8CLlAr3
P3BBFNEIEVa1D94z66oWyC62ufjzLt+JcY2NUgGMoWOJiPdPSpEDfIY/tX8Z6FJeveATZiJlU4Wc
Q5Pw75157Qw9WANoRE9VEFTbMDDnRKqL5g+HJzgpn7UaTiUPIFXk+8EN48msxwjYDrCb8rHz9v1B
mlR1UVU/Vb3OWn9R16YIALdecXXfhei6NrCz9gjkPnq7mREhcuE6UveffEpEbZhY7bGOlw42nkO8
VV6or6pFxEWri+lpsw65WMq3cp6Z1FKpHNpgByI6CesxgZ10XyuEPm0dY2es3Da6/wvSxlL/YKcJ
lCuKNfcyVcj2cfWqqkOkHwapJUuQQfT3QaU6/08sxifPkC0z4RAeJL1XqDrq0EXjNQiXpJtycoa3
qkmWehiplWKo8yfnTVGyW3k2bvzJYPasBrZOzrDNT6lBbIemXpB8UEqFuTZY6N0asF+bpyXeeif8
nyEYMcAQ6rp84iLRBNGmzDfYhZj3JcvnAzlJ/tfXe9iucHEl/cxs/VIIJtQ6DrGBU8SYft9F7ghb
gvIcbv3DLL8CSnUKJl1DXMXut8rWtA7BwXAjmObU/BpStg1jQo6dkZ0G6x9RRU6gfVrvEciJEWBB
ejjKOzPEqduLyQ/I4X0TR2mFTW9eKpyGsTMN5l74fD+RMqHk0C64PP4XEEgp5scLXu7HOfoPh+E0
IUa6qBn2nJ/Xw9/P3a3ksDeL2RJ/nny2KTcIXCb8pIjKj15GgMsrKnvSvRHYsvDFAYFcPeHmzxn9
ycgKFXxB8SWXqLlhbzeKQCtWElATcA3D/VWSjg6SBb67xrHs39E2rC17c6UufpeRJcP/h/o8Mzny
CHdvg1laG6+AwDwnsGtrmDAZksoTuwgmm+IUXJcXRmrfbrrV8/JqqMeaSsuR7M0b+3Dp4MpHeFuJ
VhKRlbCZ6+tJaDxVKwErzpojPhKscTEWgeJZaz10ueUNBKqjNL1wf9yfgX/wzcU/SdBi5ND9ytOx
3CJWNknSZRnHrSOQpXv97zC5/9DkRKufCpYTRv0Nf5LuUXquqWBlouDuY3UKlEUpIsWX2piBxQyG
0kUFx3BJY9OShZRuMtwhcRs90m8Gta9qScJa/fAvc1Qzcs9QI8syDn0g7s32Mhi3WlCsU3s+2fDL
+jKKWWr/mrzjJ+Taea5jHHT5wI4Haa7aR/SJQCzjDAnqLQt5hqKQbusr9xo87iDjPMNIWxVbRyWd
jNaT/wuzUkt+ALlWCUP34NyM8oM7mN49nyZ9Bu/85YBxNr3oZoyA5IKqQa3oaC7JVHz02duTkgCO
8XOHr1SsEEzDoPiJNNhh89zXK2YGZJluWkutnMUf23s1pjKgLieil7tHyL1JvsbINpaatL2zOY0Z
iWrD9az3v4NPoDA95BUmx77Ay3HG7qB9NQR755BvfFU3T9gZtgTvDv/mHSnNuOXXARSzkFfQjAkQ
whggMP6NpcwaNc8JWf+gtEhKbMgC04Owdbi5K7dNAePLIK3N78SCnKrpA2AiN2XME8ZHsXdg4aWb
5LRUzsF4yNV12sN6NR8RmsDcsZkjtgTd4vjrbAuZ7PbH+V+eanaryExawCuVLUyY8uqKjp2aokMF
MEjZGN/I1+W+R4clgkZdyjf/q08R0jQdd4+Oq9PE/hfc92evC/AYrTWvoEQjbxXaS2L6sRpjQ+wd
nf+jISFn1+z+nsRGxzOrXwAg1vo2TYVPLvuLSCHn4JSSgWLQbGJBqz/d2JHman6XvAqBtPCFD+Vx
3SWiFnh9HmOjsmjU3RWEtbsD06lC4qmDRBv9TwJ1dPtTU7WPTxE69Y/xQzTXA0Bc+5KI21rV7ijI
3HSMOZ8VXxsX8Gy3QWByGZqathy9/PiiJiTv5t5DfDXGkGqqWnXZmHHIC6iOCPwZ57DW3bZQwK4O
j1lrqiEENkNEoWE4wtbUMUhjIOfiYbB2XZT8fO+Jh+va4S4UcugUBMzMGe/q2xgdaEDs3ZbB5UpM
lHFcfQmQMZyxgxvL1K7/qQuxQLbOWaNbDlB+r28rC+c1WT1NAB5qFxxLaOvocdZYgzuM0pKMs1/f
8ekV0d/PBodgrT8a7iXVC+Y3uxI1aa2W2H+hX+TyJyfGyDAfJYlqRHVfDhZfTftMvp7QA0nee7fz
yXDNHFF7OEtyqJltVB3qjkg+vg7tRMKIdKAFAfb+UzShTv8dgMBFIKFPrZkutJLPhD/LSr49GDHk
zwUILa9k4FRY9DSoZJvkYZYvyo3rCFxJ7OfQRffQxcOgY/54AYa2eZqwxxOSCY+8lHPHzegCtwnG
IOioE2x9q1lbwaSuX/HZ/ueZznT1FN4ckvciGoQBwVL0rVzE2Fk80PGeZtdwH4Q/1J7sCgsYePPf
SkeVez2reSmVnPv4uSXu5gXRlCq6qmLJ/WJuAlmEHoKAO3pCppciz0cpTfM7pArX+NsCwmvkz7TH
JT/t/lrD1vRWkYSsFrUv8wNQTfPRmMQaySSP3T/ujlDpcai0crAmO/w1QB+n6Fqnbjv7z+3yMCw0
WJyk8u3KI/OMaZtbdHOv4U+Vi0r1xoTt0+gktpBWkkpkjHwyIywOPD6BakHvyjAn1g95Kp6Hz+md
EKa+zs+R96rO+r8BSvU/HHKbU0FpdKITiWQMQ7K9aifO/gaT3tzwqhDfCbUuDcBP5IA8R5xzwuKi
2ln7KfMWcxjsnWaz4bsXmwHb1hXiVsVUFVsGzlyRtK7BeaGn6Zn0KwWK/VR6BAvYS7e5BkJd7q6o
in7VVonIjxMP5SvnojGR+E5J//6oCI3Jjdot9CU+KWcPQVcZpCt2hXX+0rnr1J0Jl771YejJ3rX3
qw9PU8o9jXktFn/5hOSh8+mge//QImB/4JniyuUVGLvgFlElQBZmim1CVt5pEDPa+VB1EgsNSKCV
z0CzSF03Grki8A3QrbjFTlcbxNf7t918E41SSvVyITrBrIqx4rihJIRWRZ4yNiBKwFXRwAauJ+ky
8hY8SxR4amJi9jcn3cUA6ZrfDzu9U03i9caeDx8CWPVkjBnnYdNGMMiKrDxLsWV8kFQC1+vrbwTg
1VvRfB+T/A7VW1DFpl5L0wZa8FympCA1dB7LnmPHl6ASCdVnzevXxntU5JJ9z8axWBiPfHA+pF4g
/mSSqCe+YzAEv1pB6mFVBbN+QkYBD8XfiEoou84SFcOvHsI1QWlJCEofOpsJd3wMeweBUtm/QY/q
xGsXpSPonCUeaU5dGXcT+04PQiKYKg4J2MToZOsSLTscMXN5tHU8JUe2cG00qhLgyTjAaVsdp+gf
S1WkWIkDEwASIbxvMj+eO0GT1V/4a8VNIDyA4wCjDTxF+0WSDAfp+ewUtG3sv/j1ycaIJxGoJPfb
u8TDyDX2RZXKFz0r1YTMM/gRfK9DqXAbgqnqCC2XSlqCLqwQXlL1BwelDk5JNfTkTQIq/CiLWXNr
XEOE4NIsghA4dIHSOryvBMx5HX0Lh6IAv14y7SFXaX8tJgeWFjQ818LeZ3Kwd+ELSwrim+6ApG8X
dFTMhYhxp+kEZasl5OewWHcNn7F9q/7cUbCR3Jihy2GSPWk4c3WtesEm69cloW/48NKsOWqjbhku
dTw6v8K5dN9yg5MLtNkILSkVHWMywgndPWvFR4eObomqjjR9v8b6ktSRCMmkEz9NeIov7ZL5GyP2
PUAgW++5V8Ck9vInYRzQ3mpYFgCCsa/4vB0QPhn1Bf9GKzuxpIarET9BpEpYkCduXQD4P4RZYy8s
aVcsbCCYOiNk/TbCtwmOKIpOZJRmyBcEVaN4NBaPOl8e47kPEWEVwxYoAYCnYrtIXZwOiyo95/EL
Tw62m7qkqzA93lwOVThHCgwXV/F/52WEtHlV5Jb9kXdWy055WbqTDqGVR6xSkv97oBEbpoUO+U5o
8mhR6gI8rs5eyXdFhMYaXYew2ZCN++vkWQBAFlSRj5gwWmco1HhvKaa5qb/j5E3vxLKp0RT8qVM+
ESAr0Is1IslgraZY9E2sYNxLDCTIessak15bSewDhlcdgfLzbkIshSHmJTsYjW2GNCDL6/m+dWsl
iYelbaFHkgWXkAfOVaATyHu5VBF/vAdHZCmR+KL08GrYqEz9RqO1NF0VAL0hZoR+u/yWFtrre+Vg
IM7fQ+xWIJgnDBcfF805Ruf85LsWYNUVtnkh1BwwBHoubXMXrYRDmmykXDQgKr60MFPgkzBQ8XZQ
18zG+ffMgKTHuyfRhNHOdCvK6EAiSmyhxVyInKTnObf6UYOS5r/FRZ+ZH31O9h/0QlWzBx3rq6fD
XYE2LbpnWAaM6nkEhwCSnRMlEYxAZ6zsMwqlPYTn2neMp+9cgTvJCB+CkHlGFbuWlXMGj0aMGhsx
dgGXxcEzhPmsHHxClEKHOYXuatlrlWzKy8zbAkYWUrgaR099g3egoEmFuGZdQiKmKK/8OqnGYNnu
qLPqQBfrbwv96xyCXjSsoIgii8+rV0Gk++XDyQ5nnEkmif6ohP+Gz/z3Ha7qfYrBRS2l5LwAQo3y
7V9eKtzXPFqwjZTXhs7xwhdOvwkIMuPdNoXVERUzu/wVcMcCDGWMroHhiW7o9TAXgAyjgzct31gs
1NDKlpJmKuAeSH3xY3MBGXdBK+80Yl+N+AA9mFx/j9a7bcwHEBQlnwijG6yuOKt/7THkxgMJCGwV
n7W0hRXi2yGfWAMYF+OMgFSd/8KMuy+wNbitMKhlmvbGcpb7r6rv2GhlK04O0Fc31fDVDfgb948D
Va1pGVQowXLPyGSYFDliewELx/f0XJkXSYh0jPy68vjFRwbU2H5M8554HPmLUf3beah/dYktCm6X
aXyLqq53PkQokA7VQugJAL8tatdjCYbYi61W+uG/jnoqIpayaevDFFhr8Y/oZsy6txvnPlmYE2IN
U12cxOWMLEk0xDP9P3BFDmc88FAerVsAK6IA8xuVq850kEih9mxsGLumuOJtQtVbUSW+qFKgTH11
Lw1MCo4XCcgw3rUd2ucQN/9KtcS3nuPQtfKHrhM5JtNRgEY5SPhOYumTF44CDMUCqOUtns9cV8dl
F+tvUbiCKdsCDEQyb0FefvSsn4qxG6muSkCLkOmvsFj8lQZVxU24Kk8zZDjnuHNGzTEsYX7i4TgT
FRuoPS+TedvCz+Le8BH7pDWZDDkK7dWQdfm7yQz3u7+MbFhNhiAfA8xM8KnrV02zhWj72gLGHhFK
nHwL+G1Rc6cP6JKAcXk+oCTQK0bp1neNcb0OgGYaUMY2LXKMMxvy2pBNmU7DgZF2Bd82MQX/cqUd
9LWm/2Xk3IYsCqyVt3vFru5Ili0Ce47ROdDC87AQcxBNEHgmBv5wEgsKHG0xtdFs/OKKkhtJxSFf
ZGemI1Hje0iyFY8S69Ey7yJHdGpu9O6WSN58AMlF0mCUihqcqk0ONy310rLWc8S/LN/3elHTmiXb
q5dFgwrgYLKxT2UXFKVBQAAYqNS/c7K+m1z6idjqtfiw4Ci5t7ZDIhqSfGrHBVHM4MqVQ246anRv
KQKFwXPmnunSqRpdo1PcE0hnADCKAY2vYKdIV3IB5kSjZmlh4nabvhZ393jFYR+PjP4LiJzpz5Gl
BOrdAOf4no+Unm+13i7+mAPvtR48t+huSvSUAJzhQ9F2swOla7AtDGJ4xLJJModwMvF1M/DkdCO/
PU04CRviLogbldpdz5diFd+XPSQkzGpFPGo/6BCaNsSqgBe3tjYxpRUgbZmMOdLD8+pmiD/d0Zy8
8p/axpOS5PKIJm/SEqBy6A4KCB7F4mxk+MXe9ZwKWa0+mu6khU49Ysg6DrOT14IVJpmDs5yD8fzu
u+NZ6bFdwOZIZMjoC7umylw9UzmJCJIzvJblGJQvG3XWLDHnYgw6dQp8iaWn0GVuRIWM9VDCkKZq
gY9a7dknQtF45mqqJZPobAuEwMAhWMC6YDkLgCD6AS88WT8K7HjWF0RkQkd9+IKWhL2n/Fdo4don
AMcBn9AuibSBidjKZrPPrEtsT1u9FiyHD5NsvCadGhHCS5Ry3OJoBRYHYx6L13H+NZyZemNGg3eP
4byScBeHbgowoJN3xnmdOffTtseLKXMaQaBZqqp+BRYF2BIizHpNfTOHiYqTTK2cCztdYqMNXH5J
mWqVaS87xuYxlSdblVhSARgv+clk3p3ELPOorYPI9h0KHFOkcAD4WOkTHwJ8oBJSSzgS7UmKIGrh
KmfO4gB0nRgcdcFe3HM6rDdKDRnbwFMKXUx0dEqgqo82RpOTtzsPnjtwMs9dZHdlJSCPDBqJvvuq
JBmTLVQJZhgATpqdkKpfMyCYB1PV9uLaMWAAX+v+6+eObVu0ARWu9RoDAoTKjRHgj/YY1PiNYLto
9vUMhoGdMiQkbnM7JoMF82Fx7gOc4Q2jkYJ07Y4uDVK1a9pIb5qBzUYDw3EgZjNNwy9EOPBvbf/z
6kBlkLofOUJ30PnUo0y1ymTZw0zgrq5RsFzDarhnu7+CAOj2VZc5rn1QDZA3+F5rtueCv47arcEm
ynJtbn1qA4SjBdMlVgXqk9V/0UGkX4/Ew1YRgHi7sfuHk/2AFhUV+AKByMfyFpthwpW7N62+k1gx
dWMj/imv1zqTCpXFdRKfKV9H2ydJbGPVLccP9gjM6STqUDurr3EMAqi1rnht3jrmcuGAlzIXBkA3
8PuxLT9y7DQhfPxgqUXXPaGRTuUIKxfXBVUdWNiECjOPzOuZ+feGPKOrsZfzC7Cj/E+2Bk2XrCbC
x7PyUvbtTPSuMYCkfUlVU8HZNu9lR7jOm1hRKR0B90xr69/FLYIvvgj9xFy7abe/Rb+3+TO5UJby
I0SfcaqxsRRWxTG5EROLW3Q9CbTTSInClwiIycj8z2kypUOiaNxqDCZS9MTeqeJRd0QERRLE86yi
I8UA4Eyt1wxlyOVXyfi2foWen3Ay4UKavh2sLzOIosw5hfOOaMk/1ph27jkh2eeNuQL4Tb5bXEg7
XSTqSvfscr2xlFiaKeewWTJaVAhRCjaHDAtyoZzSBuOggRgpw5Rc1JbmcMbXE3Ez9B7FJwkV72M/
oJFpEQt+EVFFNhYI0pP/7OblUq8Sv0kI51W+5uVIhrc/+++FCT20TLS1cvZtXCBIqSfAO2cE2GMc
dNWaxmOTuhYqRd1bOQDg90+xOwuN/QzAB6Pc5s5ZrTLIg/OExjwNLIuUSMfWRjHmq0zAVnLKV38/
eXeEuw4jOpnsBxlnSke/pEKfsShYXjkI5+hhx2+sQXG6KoHOH3f9//IoqRVVZuzFdY/LAk2EMtlx
PV/ZMMFHNhDqjecn3eBZm/SrSbV47secFGbR8qRuNIjUQ0a27rcZlm9lOJCiaPFIzRKX8hxHIeWP
kpZME6GkxR0XhBRwrO0+rTcxktis/JxLtDVmmMCtj4ReVkpJFGBGQkuNsxHig6d05NJVA6CfBZVD
gA8c9tsyJ26qtWgi12mMA8YUo1Q/7cR9apx4op+r9I2tYy+YGpn8FppBL5iANPPZ+HOwA9zWuxg/
IadGtq22UZ7WvZRUw782tuSoOloiq44bFMks1MnIB3F7iQ24i8NUSEy1jwpf5DWB1go2t3NbuUdd
gAadeIGEqzIL+exlOBvzLrCwLVCq1hto0chZs5hBWP1ju3FQAGnq/BBBGJQ3pItswYZjIDNV7eqP
1moLTOIlUe7NfvGaUUKYy+dtllMKsa9m++uR/dbe6wcPDNatB9FEcWClUlsEQx4hl95JCQCGqbDt
qFyZ4E9E5kTGkZPo3Q85fMZf0oHOBFF5wRaL5J624pa15j7NRVPdUYd8v9rFbMTXd0dZ1+1Imzq9
KLz54OM+r4mecoOyjLl4znIEL/Hghd0+4p+2r6lVtwGLeHMHbNq5L5jyx5+BMwTullglEweMKkUL
vPOO3yq1+tGNz4uEjfvfyqC6KxgH4CXBmEDk5cqDuGuA+OI2yvn4cFBubYfE82vjj2qqtjKGn9h/
rqeTwx2GElHPKkKehcujQviGNpck348tgKDp1kAQc1dXSHfkuV4FMtT52oTpWaNLNMXPmG1fl3/D
YLZyqg/5rvWgTlSGF9eMtqxqGZT6NIEt8OJdRdZ7fm2yYMu/cFGZuTtrZB8PHef4T5o6KxpBY4w7
VplTPIHPZm2tNZ73SM9DIkUIzc5XcOiPUnd4cZMd9nEqK9DK1wjvjAK4lokM0Y6awmx41BOlBocf
YSnq5Tl0slQ4pDkl60IWXwBy11wp91PKX50vt7/s/v+u1CZ+psvMRqGklCywv1kXgcwSYCJbSZ2I
KUxf1djaBk848HJEoX0UFZ2D6KqTiM8ORjj5uIwuDDEy0bwrzMnlGQKvpu5cSmG9pLwmCWBIdmow
HjuvU2Ga4PmB0mYKX7VrJJfUDSF0IHbibWJ0gSJI2Jie8fi/L10Qz+Y2T/gjDJU5uM+poS5ZxNSr
Jlc73e+4yzdXDGow5S/gH8k6Rrw0xz/KGknB3vAXhvezHueOAqp/njxVXnSG2SXTZI/5aRiFTAjE
VfRIR7D1l0a1BnewK7gT3dIQK7KCERvK/sPElgZ05LMMdkmIM1M7MFOOKlkLLj8pPdWu5TfwsApC
Z6rmga0DP12+UlJaAd0Hm9RD8scd/7U7r27WikwfxMvrb1CUT7H9kLhWOtd9UGfPaJpbja3rKmS1
WXIp2eTURGy6OtxPq9CLj58LuK7DNKg6ifoDiQtYz2vPXNBpWKqGa+pu0ENxw4OFH1f0VJXPUrQ3
PPZbMqwwD53/8Mso8/mORFanI1Sjv7N7LkoqU0aWyRyHnRKdBcCci3etnbgtFOve0qlv0BjToFPE
SOd6o3VC/5Xzf5vUg2J7yCNGlw/sS3jaNhHQUwLfyaNcCsmaLTvvUd3UjFVMm1IDodJ/J+GjCaRd
JfLuQ6jfTduppm5MX/OfCgKkTKRlHPv8nI/lCFt0BYtFhLqJJHsLIGvnAcj+V7SQ9ARgpLnO8f2q
HJAu8Mg80A0lVlkGbVYVeUNkii+mIbtx3TRO+EEzDk7eVfNIlEGipHJ09jCo+3+AJ/Kg5aXaeT2l
bdnRHIFjHcQGlowhRpNNhlkw6KRi4gh8U1iq/NMmJIwR8S680J7Kh1g31sTb1Dgn9FCJTctE8K4o
zPnWL/AjtwhfmeWeshlmr4B5aPlkqkiBMNZURz9mgMsry+hu96xWyiE6uOu//yqnZZncN7q4zSY/
0L4R2y+tdVeO/s9QWFMa4ILPO7uMoHdLWe5ntAGYXQI5gAKBDbpyK5Ht42q3ZHAWp+RkV6+5P8zW
fEG1bUt3UnZ+l5ErvOAKznGxN/UC1GYNFOa3bt8FFfwBjNdD5g/Fhki9fNBMN7x1i06F8lxiWeD2
H9BZ7W2nMx1K4Lo/YURZR2Mr4tjqwhlGKm3Quy3+bxHodGdcX3v0xEy8lOlRx4mD0saRv40tjNkz
6qP6ks9j2Ht6CK/cSoAA5RHVGCn15NzjXBfnrXama9/krWzLEzaHMG9CME1NC0d5xv/WnSH3Bcb2
cO17ruQlSGQXTGQDkLs+V0MBUBq0raUU2B8UuVdAOP1LjMf15LdSDv6psFG6Ba82lU4n+9GhdlF7
dNRvavY1t6xetMxUtikbuEUwIlzCf4YAHMBNNxhpPghwM0ISmQ2xnqo9qlNsxZ+/orT9neebh97p
pl9z4ifL6Xo2M4VsPg87B7Yrtvn9ff9ZtU7S9QN5moiwh+sZpUfAtMqcmPjdhvjp7f2FFrs6SgIR
1vj7DEqLOAsdPESrOAMotI8tTBKvpyYt5sCDvYxvTO+m8uTJzTUGbwCdte0cz7ih2xy837F5/0YV
XpyMBCPoQDPxR5TAPYR5/Mp9OW26eO3vtsZQzJinQFetq8j9N9pzu8GrUsdCpwpbuDS71JMvsr7R
6KZis7FL+8M0aovA1Y7tQqYYo10VnKKVPSM6JQpLm9LqCEYHXb8hZ42/tjn4/HRrsigTOWnStE6p
ZOGXo4lOnMt1KYBJpGJaJwXMG2bP2UI8gNfrg2n+5Do9KZ5YQWSNf8rl9If7PweMC1v9k0nxfptI
O4Fy3z7fCF4KWjlX68ip4U8ncf6W7ITZlmPjhmEU0DJ160O5lokKWgbHBjn5kD1BMdSIAJcNqahh
d69tFKI24GnHcFulCTBuPX5ot7f/zYaP3bit3vSXhA1NDqvqWRh2OIsCQYv14A1Tk6h8zfmcqJ6V
s4AgzdowyqI8Cf2RMFlPKwD96PCPyVezSRKXUKO/vICW0keegbjxzi+SMpOz6me+SyiVTNOvr1PQ
bFt4Slo+3n1LcMVL2XWqcgL1PWldFtUaIn6x6ux513FY1O/YRDyddm5PLyRQ1agmPb1JjECS7lq2
n8tW7f+ibH7LJqW8rkqEAH5UrKJ8crCLNr6fyyvm50lbcNPnxPWqV2+zEhkEJVW6myHuKVVtNrAB
4jf90e4aZC4xUtSaNEcPi9BXVlbEgmZVCQEqanvbuYqrJUN5n0U/lzVTcb2h1fzctNE+Il5FYwMX
mOD6Ud6srwfDCC4FkiVZeaon6yC/SQ5UZitEWwa75gw2ZlzvR7hxldFX1oviUCrQpubTZdncGLDT
Ccb0XrcYwbPVbXxe+yf/3gHTc6Pt4n5dbzgNBFRnLtP4NO/cTW0eOCcYyZ2YWA8T1/+276hIDHqs
TgqNpRMcNUDY6VSy5VgpM/n8L3rS+Rtd2AUWD4p312gJPjXDbbOdVBcriWEcUNNIUtxIqJUfz0Xh
gXtCnsXdwPYwNiO23phOSl4kOzZph2rJ0cgQDfFU6Qww6keRah5Cj1sldfnSKTkiTOnFDXX90c1K
HlndximZY4+TXUdLnG5qgzNfXC23h60NMkzBvzx7A4+y7JM7Z/6uINXh+LvdU7tYYXV+bndOkH4e
dBhnC3doftbF/kaR4E9IXC4WuM8iX4wzhJCkgVJZ3uTdW8j52+SYduDrzHFqSB2cTvZcqhgbgxPq
P9HG7zfb3/Njz98wk2RQxpLPIL2HJ5/IM270Lz8lL8Js5A2PKBObo6ZVmwzICnpJJPQIEkW9Oly2
1rwuQH/iWOGGJgeMm/PYs0NPgEB0aZrgsH81EOWZ3eFwy75yA3DeFaJ+dKr+g7bs/5eMHC0acgZq
vPZeKLd6Yt7/r1hbLaoscY7BcB0+G1AyS5KhVS0Bw1Gll/BDqbLfso2RBlxFBo7LpJ19D1c28EuT
yv1OupVO/dn8UgeVjbugOYuqmyXXEWk/i950Tn8fW0v6pOGhk1okphtCd6KOgsvgaPvK6bIIa/EJ
vMFPA3MOcfMubWSKg2L6uxDhLgCYXt0lImp9HAb3NIvb3/Cnf93j0spWPbRfPP0yhKKF7D3NzFxw
jZVX1S0OkqJ8UmKf2uk2lTcaZYJ3TYEQM11slx5Z2jS9kZS8dGqRFXRcIC+E85IOB8rsm0QrOwv6
1RCYVlEGGFc60dgIIHN6CswN8qesBKJcKCXQaLh2tI0gTJIEa3XOX04TL64xxQTGGAXlWISlX4kV
b5K4FO21FljtLtzZKpBkRmNf8cBi+3bRZryn/m8OdoCZo0yoZA0kfNSzDVsU8vXfPR+EXuqe0U2+
2DzUKNKgnSHe1otwfNCtF/c3MRq7DvlWGwo6Gz4kHhw7N8fPgRrovLU0ysDZovDMxYKs1R5dWibl
RImVq9zZsYp1eG8qBTE+OjpwjjccTZyK6NTf0J0yQqM+sugaK14aHsLe7YA7XKbmkXR9aIo29i/Q
wGTm3psLdj2KG3fdN/9N9ab1GASu27tJ0AfuY7JL7MH4hVk8Is5pT2B/a9ry4qw7DnK8roaAUnMz
W/vPyStSJ+MVQ+gjhIb1pZn3fz6jZDjfYu9MR/d8ByvsI9g38jdFGaSQEUg0oE/3lv0a20tmFWE3
pTZG9+3459R0Jfa5ddOqoNdClMhA/z2LwdIriXxqHQrLMA7e22M9nK+U0bSOmDcYfCsI9j8ckA9l
Hdq+hYdmIxaYC6v+hhFsdR0lI2qEhfzwqknA+X/Uc7cX+xmzoUz8aPC98dy6Nrrbr3SP33TRR5mg
qcG85pM2DAHqTidgagXFZqA23wNZ724dQ4AckE3OXR2gKqNCG4UZpIFaWNhn4njWta/WzNw/CdX4
G3Tk0+hKKG124iVnmDC888Hg0R2eGXKbk7zzfItikP9J5Ca4gcCtd9qJxdpzMEJHVQawsql9fMsM
C/UWOvNbjtFl8AR95X1VqfSsLv3sasuyWn9n/9OeLDv8Vp7/lH5anv3iebqD2NnSsNU+4Hj3kp9d
wiEjQEfwr2Gp3uzwAyZc6Qba3T+Lw6gkc6mJVyH2/LkLTO6+wP8Eb386Nu+TSClyg/JYRNBY1J4Z
x8URftSDbhOLHXwWMqTTnaxD36JRI7EA36REmNyv70A8ZeryyuqLBRo9elp1NBH/zv1c/Ij/y3i/
oTNeMV35ltSU+3Bjap4vViltMOoDWoTqeqfiRRPmR8iYW6qk5ba6iV6Yu6D+4RdXkeULKUrKqUBt
VchlCJ8iwPTGp9hWM/Cq8w5rTaPICaB4hCsPJeJx4mI0fVMo0ORk2ATgJ3M2+pbM8679OSOrwhBB
50xdH/lhlE1rCcIzZrg7Bkt8W381eWHrzmKWSjg7d5gYBF6E3fUk918z0DjasYf/OUXdbEE+iJOy
aYRyDCo690sf9RCrKil86ipnzvUIGQW2oaAEyR1FFKa7+uaAMeRV1Uv38CuQhNYk9KICrJZVR7VL
XE0o/NixGpyGyDlLcbvGehSLWCwGfQrRk63/JvZhL6JaE7fEr7HefVGn7ufjo1oV9+nguv6xZ170
ez5PyVBHjb5llljbsPWT8tVHDn2VtLewPG4aujxyt3y7zl0QPDp/TpBA148QSR8532FXucmkh1Au
O+aZgnSdjLSPXPBeUQxBTBH2pr/l52wXlfAsR6dAtt1uAdEz4zMUn1/r7PRM5XyhdAGeT1b2ckgm
JjO87q2ohO1i7ONYcKNYNWz31JgHW7fFWPMa1+OK6aAS2xcrkuHlWm2IDNV2DfkW+sGlOZNu5cry
Tyyi3buQHnDvTOPjN8BZdjVrZK+dONYjtobithUqhGgwqJJYoWPB1nAm4KCq0ID/eBx0Fp5pcVGv
sSJsp11j9+JUwVxWzW+J9/ZoAkGEWyxx2c4H2oilJG5U92pwj4AtRENBAPk4v3WKmd1QKQ58mrG3
sDW3wbYFs0mDrqBbd8aOsaW3VP37wJXaxHH1W33IS028/D3u6oNYrPnWXdXVcjEvxPmI9Y2sfFui
Bn3dcH55vPvSEhEimO84qJwXD1BCABZLJg3AoWXqZh3p5O8mzhQC3sRDQK+vZhk+dWpfDcTAtZtd
T851HdRah5QWee1EBvT4+LcLrzqLqrFL1hj/AvbVLbMxPcFv77+HucJblpnActsR8t8qTK2C/XgC
JyCCGn1ZeSgwxSIqUfqoizkeM4jvS+fr81ewUCFNouNRIAyFFwUa/hrk1X28P7q2lnh8dV5UeTZB
w/mCegnqACca3Bwcxo8ppR1igxnrqUvCevafHzTSjaInvan72FzpMUIc1IHj7/f8jpIg/E5R6EP+
a5VIDDIMCsHkqGihN9tEpUZMlg/t/OMgRg7aJIzwt6iCchzTaQDC0FQO0PE4KfxpnviQae0nlW6y
h33uhargagVQB5baD/5/A6XrHN38eW4pLKA/jcmBpobU0Rt8OA8obW4BCwLAXPbFqZZthajg9bJx
EMLpYWNsMprxKiRj50KKexKPyb8S1iOQgzrQtJbMTw/QNHYK3Ad2D4cDsSVO8wjjWSqm1NKWqh1X
fYNO88W4JUsLmujwrOg0+GMVyUWtCsDmOkbAzFvtmH6Uj++/IdjbpFGOZgaMYFBwteRIavRnXt7x
gMJ003ND3kQNjZ87Wd1DTOcnDXIKvgSEFiZj8jGpyquVwQptiaN87JVA4OGFtAdPWJTZJDNsUIfv
km8P+sjr4kPaBy6Q6fwXlLvDbeDfjTKNafhzkJtAmauUYI4AioKUXl1QMjbC2mAXuFCRrNhIMoaJ
OUxO+BSWNKWFS0WSw/t1x7hYuNwsImUR5ex0jp42ssN6TrQowCh5SI+PBaMjt+mxqElmJrznuB+w
+sDto+YjP5L34wc4LnVcbvRfet5FjtDdqbxsw0a1Bmx7dyGFuwNhlLeTXoVkQYqsUaSMK4B6hiYS
T638ltrMWIpyW/1UTjOKNWB2eZDJXPps3Ks7eGlNu9MGDY4pDd36KckT7J+T3i8Lwd1ZSzUToMQK
pt60K7PiKfbWjTm+B8VVnVypF2QhSMGpRWcGCoyuM2zPibMhKt+3ncRxG18CBOZcKApW5mhotMVN
Hee25QsThKl104/oiGkQyQyJS2ptla3yCoJ+/dFTR442P1XGyMI9GDKssvjfrbXU5GacI3kXhp87
wGHGG+6n7psZDgkD2PaBUAEviEBQ7NDadznSeleI8WVWFIA63zR3C4j+g3ZrTx0Iz/QbijjzVq4P
DX2DieulHWpNkeGMBI491KKaBJhD8/PcO1GNmtugQ13xw/VHR+YMwym9fkwwXoWCmyUYmx3ZISMg
N6SuwN7gIz2pnwnA7zFlo6rSVqMUVRGneUjG0e9NkqRDY5CB4dGcprfAqmzjLRVvEh63jjsm6GTg
XWI11h8w9KPHOqCrElqLZPJRISHA16OlmoFmmU2+fikPp0qoEWeDTbUv041+Hz9SgfJUjJDZCFk/
rG0mSFF2AF+YjAHIBRwRGOsUKA4G5NHRP4uaj8TdYyrL2+Vt5kgTvYokyX8/FBwdnwszfJDoG83i
Nvd6O632HWjKB6/+4KB+3BnEwkHwrxCeP6UwDyz2GmDc/VVjaLHYvjsd4DaaJ1G2u3/4lEfZHmBq
BugahkNPhlGI1CdAQqvA/NCqoEeTjVGxiRf1y8XMs6Lki7/qwa5YCEvW2z6OhsGkbyeCt008k6DW
D1FfnSr0qOXUYsreABMDj/t4AVY7iNa0J9U6xyLeEjMs2ZK4xBOBZWv4r+0UnLhCXYSqAbSoUEph
wMQtRUbPs8UHxJTIRBtp0je55EPLGenB2MLCXynd8VzsDqwFVXJTUAMHoEyzfBKWqUzMUiSmimNE
lSyi659qETHHxse4cFUBAXhLKgmTWiPaY302vQKJN/KHpP27MMuCW9v0QSKW/jiXEeaZqAJjgWqi
9b9dMajNL781AXlzU4yG1gKZtDNCCtNgM9D5yXc4cikoEIYKio3zHgLv3tGpBGgCi0ycWeFpos+t
xZTurNnxjuTAWGExpcy51jTBxnSi169zE33s908cQJ9bwgurvs+puBgeUOZgh8a8yTVOx38K+5Ik
p7yX2Bi9PtD80Gx003qTN/8otWuRcr9CkDttx1ejfuIqLeb0C6hjpKtNjglO9XCWHBUlbcVAbdNz
/8+6h6/3fFSNbrbw7L9PuBFp6BrNcCmKGvEaGuZcyOtIceOutCzT6fYRG579oZMiSCmIZYoKK+6p
gEQUrzjoK1RNiD3pnfmC7JiqoJcGQ717Um9UQKg0dBa+ETLX5p1SaZK94A2i1HHRgaKDjjJ0WDas
1FYQZ4WWxggpzWVYkkIhLGJ65WuZLDAxrvJ8ZWIZZkgUuPuANjGgnXcHCuKJ3/4YCOgmcwLQ9az6
hpG+bXqZv+L0pgEHkCngTfyD5CN4/1HRQJKzyBYtmUvPrzD4cieM1whqzp2vtbbyh8h7/bbGtEuC
Q81d0YTUZiN9t6WSRaUVeOqVnB5STPHPZYOsc8OfEKc0VZ2YOxhoVO0q/kOvDg2Edz377e0nu1Ge
4q+TVMFyRDuZ/9995irk7W9qybyeHqT46/XVQFCsuCCU40ZVPPhJ5I+vrtXvNFdRztfre527C//4
Ujg3b1y/wwxPD5wLb3zEgAGbclZSQiMgqPPpCAc2Rm8jbTtwK0vH9bdT6LAxnRFWmAhMZ+x6TSEm
4HbBNGle+8RiGkTiColTxHfwQ2cgnUfDDfuXNnhYA0JOBInMor6EEPdX9xkJK7+YIazojqaBQ0Q5
avLdt0lWT9Ho7RNxARdfa4d3w24U1CTlkHlpGs8WuErZ7UK/phN39vHpjfGa2gx8kn3lrWDDjykK
qb+LWggCpRrsKhdQQVf/x6CGZNDylg/r42C7MHWE7QT2RV3jk5/yPN3VIgUVcal9KMduZIsIr/bg
AJFeshpa1ykE3PxYmwfqhmPfh1SBsel/qpNQUCw1srkLERulaQl5lRBoXsYpy5lwLViL6hrQ9haI
/Rb8RI//SfLuO/cZlDBz54gSU8+h3hYLLVm4k8jpY7n9FAMyM4cILmD50xcE4yqyOFng8YOFkLIE
LZHeg7YnKIbyBrWTVGLC7jzh1cXbJveMq80vbKnp9dE5j0vRZ0EVnCscG8SWVJkMZ+TsiVnAbhd+
uRTO5L/3R2NkxjPjTuLAudFBSJKQ5Gn1euO8e4MzUnNjuT9W62YCpuJDtOmhqyA0rJ1Rka8lUmXC
QocuvhLDbXOQZejGlAyFN6GBoyddpE9hTnazi3KjFpS8pJVUrdH+yvNAaIaM6KEl9NztyTcA4qkD
J1RXNAyxlpierp8GEGS1TvkAM+NDWqMFxEAoD78XzOmySDRbk16z44GIkQ0Cew8sbRakZOJMJ8ub
OF+SSfB3B94WU8aEwWIMP9eTAag7jQ2qek96+d0Knnw4c86/ESTT/mJ84fPUc25VJOw/2wFcwRjH
sHWnDbMr0BIEd6O4XUndeD9lbm9/iLePzQKGEvXnFNynxSDCNKJFC4irWDNvNjECHNi+ZRE3HbKH
w+adT0oq8LjjPx0i9570b9HsZjN+xvHRrCNdXwVx9W4YCKXp64zXm5jcKq+PL0PFn8KMxwwNsb7n
0OhpW3Gc//hh3L2DsM2cGTnj2Radp4P68+OVxROXUZ5Z71+KdeuEMJHAVhdoPmsqHbWIStg39GJT
Pgn9OTWlgXujnGck8wG9UAHevEl4RyBbG+dF0lSvEov6lYY65WoRaY1X21+qe7PiUt/weXn+ngkO
PhzAcZl9KRKBX/GauLx3/PqpvUgXRK3SRFJbANnRn40z+04DcH23KZ6jCEmDB1HT5DAlb2RDgkVf
A7hK+XBxptFtGoPGx6SPuudqddPMKunpG9Rn7S7BIT56erMoP5iDj3ZN54eAXpYsxzOklle3rnSO
tUBP4EQfJc9JcmvQdYSYD+sqqhHSXyXD9L6DyJLwhQqQuMTRD+eB/9XANc8hQw5EiLj24YlJuA5F
inC9DUyEm/cnCE3MXbPWw/UMpFkZN8ozxlbmTGnRDPkFbu9OOK1zBwD9qfmFxM/znydvFb5Rd088
1oAmwpAwdM/o1WprVhgwValWAf3iC5SVtMY57VJdR4FwGiCXcAsOC23MY9b/hNLnwpnO3CVGxeil
iJiS5fIluSlUkCAOJvolptlHxDQho+r1aflUZV4P3CcoFmmFj4jfuyCQS15M0T5N1iDrYdYo7iWi
+aNVOitMIp1+5URNfNpxiigVJPV+YlIKBgtS58MwQYbVqmoeJvXRwjoxQKcwXQNstEn1qZOwH92r
RmXPwsbUmfJ6c4s+gCHmql+jfqogWB8CMpuXWqLN2ebzmjFM0iHayR+I9IAlERjJ+wOj/av0eDD5
01Uw43K1yy2/p032DXk42mRt4bUd9X5FDcVpVA7sUDWPreA64Rtl7Ya2v1qOtr+Dyj7IbV1F7GdE
5PWLrbEY1Yt64OBRiqsZLIitO7DJ92YJMVhPuJZ9qA6oldG61maEZ+bZoIY8j5U+HwGRo5KGu+yK
iX5ikRh5at9sK6zp0AS1N7TwC+sg6IwOP+W9hKCWgYwe96HYm0nBvmBKKM3JRq14augDq1qCbTQG
LiDnB8LdAwtCeL5wGGXBi2iSz3PgFIMYXvJ27DdXAVHVCc6fbbCMrRcE2gnwmFAWsw9YbMoBFEXB
5/b7bVx0a6rdsE79qTs2Wn5czbcoqSkB1yeJItOOgOiyJLahFI9IClnSz6lU4A5xuTj+El2ofZDE
xkUXMmP4RxqB/LKYP0513PGY4AB2qDEXo6QYtZwqXeoK5++shrNE3xug4IMVoDJRzbVanzOBb32w
B8AcrzWU+tc/mxFuzCfWUClj1WGGp32CsLb+VlFsCZs+qAGd+l8h07Rh1HJY3hwwDDfMy3NwVN4v
quPWM6Z5TjRAmRFHTY0cvJsL7S134f1JHssWR1Kn6VjXj+eNzjPjvkGEllDVmBmZvczwRTREKfZz
wvZ5moP/SMsZlDx5zRaB+8REABwk0vQeBXNb7tMOoEv5ZOPqQiEbs0cX4Pr/7l930lhN0f7vDXok
yJCQLBuOI8nXUEWBr99vdrGEx6LU5ioXwmgEBhALKQs/3uUU1X36gt6ejNDAJcdyAHAhf3Wf18Nj
r//5lG7TtmMXiRR3WIhLryVBXWSgRqf9qKqmbucYCvweyEOUngFH9fU+E6cOSitzsc7AATBtruIo
I6LpGEvInGa7itxhiNOJkyWAYy1hn/nk55tVfU6pZoAYf6e7mqB44raY7APGRAOJ4k9zT0MjEm6G
ZSWj6wm+J8Dp4Th/yBEY18uhbbbv50R35gqn6/mAzyl88of6Xcme2AtzUvcNPXBzp5l5pi39eQd+
CWLcKgRVXgwCKiXemUtexlk2yraCV3ghc6ZtJRuSAQE9SBapRW9TuVz36+qfV/FEqVFOwUuQmFDw
iXkGb9kLIomuu7N/LgKzyCKKC/mSyYNabCytkmnyRkRYMTzd3b9r80rUEkiK5oFLIoPc3/w82+hJ
TMxF2iL1Abonj7PtOnjFwTt6+1icrmJCI3bXPLCQqGXxtR/FM8pEbtb1IWrUhrFWislfjQ9xNcdh
bG0JisJBadozyUxRt94oEK0Jnq7nEUo450aNwL1Rnd4A/sKvDllwHlSfTIVBaEFfh8mRNecBRhqA
uNDSSilU4dGxNvAdgC1pOvpDncbn0veanZXt16eiMD3Vt8xfqYp3qVnQucb9xg7Wty93/XnX/u6V
ZQk0LrzFLk0D3W87Ol+0YsXgeXNIHsFig8h5a2nY2RjMOcBJFPPAAqyje4dvWnSgaRo8QW9ifNkL
64RpeBOnXEe6dAcLYvLBw/0/A4KQnXY1UxE65BGt0CyJmsWpsiXMFFLcmHyASQXPWVBi8T0D600/
9YN895gDF7xtCHaxlaCHEW33jxpwx/zN29Kpavwy/j32oXHYe6GHq88OrUiXF5OyG2dui+WVhPXB
IfPkYqVX1vi8jGWlsYUHKx5VLZ0PX+d4vnC9/kXLU/xX4CrF/p5hdewjG5ZgMVckJoUObTtxAt2H
9NA1SmFeXl1OlukOjDtAxB3r8NaczPYTyYKDxONpluQjfPUNTYyB49Qob6kxbL9t4QaPh9sz49Ys
f45nsPwaMZxwWsv/rZ2VP3CO3Tg05C0Bcn7W3kBltKz00jqo6Yj7j6+umWnL8i/HSbsZFwe/J5mW
zb4WjsUykTXDd+wt5AdQUrp6EBprfUlM+WAqC9wCmEGNW7zLh7wcu+dh9NQ2nD7/dEpQA6um2uBv
cHt8SF6/ng7TNesfMXCQ4dpzL0zg2paWLyip3l+4CWCj3gHxZFXUuUwuUxeFxn71cxS6ONc5Nn28
MMaKId4xzteeRGSOCA9W8dFv3pTxzkGf2luvfu3PjlMlnknzYIS3bR3KjpMh3zqdMFlB2yDqRe7e
mfluqRDt1yrJyV758Id0N8Gh5qMSGdE43OVApjTHMa/DN6WoLXwYcamNGohcbrm1GlUweVWjLM/6
xGRQ5W/GtatsZ9DIr3PqeY7ISjvSFeOX6hr/etMlOoaD3/fG9YJFDAefNOfC+5bB/Orqcq6qNt7E
TtIumYIhVGYdEx/yCacSk/oYcfErZMsHTeXlGMeahWmdjbjzDw24duq5c0rtHhMhX+65STziD4YD
rL6aa/FYhB/39U2K8R6YeJrpZLMpW/eronLpnZPJKlRRrjHM/5AkRTAAPJK9rHZHFD2hsbXzfntt
DZWCvBmSfFMcI9ukhCqI8qNYf2Vqdy/IsNlS4sGmYYLTnQA4gEKxLU+Ma77XiSobeu2F2qkSuV7o
M4yJWuOW9Ewzfaa1ziQdqtzFI/io9RZ7z6YbW20ngupl3bdWZXqC5yMJQEphrDtXTxLirVfUAOhE
Sf31rzqspeV4yIm8IB6IgUP+GPonw1XfKXZLuyJQIZUAJunb4sCa3DFwI6P4HOBnbCz30YzR36fK
nteqMKv78dgGuhZ3hw736f0GvbTiJA59q+fFH5c7Ga92yNxvElbBppTzFS5QFnwIVN5+WEyi7a4Z
SNGN1FOfdtomU/YMDVNA6H9MxljqMuWjJYR04UxJjXj+BtYVDSh9tOq6OaRF0oIoheDncmkcqYdG
McRGv8x+NAkTbuanN7kZaratuvVJPIV+rVONjyi2aITqbGPBP1Ygn6yJCDMSJyN083/S4t17MSeq
DAP03Nq5M4TyB1skir9l+imdJFWzA+QJrKSwxgfi2EOnojfmGDpYORBx/F74r5iR3+XdU4P4bpuE
7Gbg11HG7pwyfTLvX+eVlRtP7zD6Me3szWOl8esYnjhqVYe76b9cwk+zs6rfezdMV1Kl3jPla3do
t0+7/gnmIHyh6fmxwYnTtMkVI1DrXNvYMsXGz9CBlts2N5BrRubWFrQbqTsJNS/TT+DY7aKrn/Pr
ia558m8B3fotEOKm44rgQf3PIlOEa408MNjyNYOR6e7ADxpTzp0eSLHXJiBTOxuyJVolFmkK1TxJ
OyDe8qHt27WisN0wPTWn67csadj1zYEDPz46spL9Gj9vnGML7nevecGoxz9hErcTfWdKpiwoxGWH
t38Fx0Yddn96dtPelmVnNwOfCiv/7oBEQ9FDPotMTtwMjkJXzK+mhGiyz2ilf7206J5P/j6A5qTI
Wc8js+YOhWh73MYVqwPkjVihIEDg3YnjTkZcJKWJyUEPHIws4XD2seabyon7GgoWyIZLrwqaoMxs
zdNOFfxRQkFZL432pg0YDgtVSCvKHSi0wLxEcDXpVOXY5eWgcfzwXm+85qbXNZea71PpiHvd6bcr
kI75lpdgZP1fnbYWUwsxO9zNfSsOPqiTasMjG2gDbZ+mIu6QvHmL7/tO0xW81K4aiGKpsgJRT98O
dp+PJm+hZ2heuKpCfdCvEVtREpJeQBtCBeszdaq+nzcsXgU1m1Czxjgznnx8hrMpL4d+wdXI+W7N
ZQeDt75T5upetwOX703EqMHurZFiKZ8HtmKvegonkrFvlDQfx4jlwjLqXj9Rr1zu0krvPA2qdAWz
bZn6QX+Rah3FuIxjnOhb7VcQewDCW/N2L0SCS4gROjt0nvQRoT8ch/r8bYzUxrPgm4dlkiXzDYw7
HYzJwTYHR2CI5ad5g6+EiELgoj1IC3d8fNgoSMdQHDI4UKX6CbLmcSD4ce9H46EyEce27YUZpsCS
6V2dUy7mYrMh45KWpdokaK5Wf5gRAtiQSsMKAnkqNF0Mk8b9AuAGGn9pV3A9DbwldGkfDbglf8Vs
tnbu+WPHgqkaL6GLgOdrIpDPpGd1a+fXx+SddiD3yqg1uY0D9AllnOSF8mXdLUUtcbo8vggESDyo
ktyvjV2vXSwTYVGXg8bTawVnt/RJZ5e03dO0tI8zX40hDGIT81faQOhbGl3VG4UV/vma4qsZ72Zf
DP82BcAu+QS+kVfeEQvbsR5c/tOz0cwuihRHnfvhACC1N3LqmN8cIMTKe/MtcqFS0DA5Dd8iXAdt
f/mt6nMT3nPSjsCPABq2u583WPW32kAAsLa3WucjjP4dEp4uKj1B4T5JsA6qFfZS0AoQzccTvdDz
+EaHzsHeTFa5S8AiFpZTvLv0FYY54ZtpiI88W6ncQN9A53DK1dJ60LqIbsCx8m3QZKv2Mt4tMWmP
q7b5nA1zetggoJ2KtU2Tad02/dTeYb7+vfmYMJH+4pWS3MNVj1C/8lNq60n2IYKjJGomXV2Hxw1M
sXHmMHh8uMhwrSe3XILhjDFambozwMVgTccYrZ6AMqWwB1PRza0lXMMUlD7htOmxxgejHYout3tb
txl5LpWAkx34DpNy8pXmzsZ3vCrBcyf7bhWxbowLWUmRYGxpKHb8zFKCyxfTuq0fpPRyJxESHwCr
SUQicmq25orRSXtj6m2X58XsAOXJUVvDM1Fy9ms7MSadSfgN+ZNrkutiVbqjd5OV93iQcVljMaNT
EaqS6eDXgYjVhTbAKkEnh4HibWGBzMuXZlZWbhsC2s1uyEAERZs9jZDObDIBvmunJPa2hoRUrLN6
oNUgaPtwBzEsCOFsvVGzA8nJI1ILHOH13bxUr0faGnDb7FxxjpB27tbbZZgDf2g38S8osdzd0bEU
CeqZpupkMjdWsCaR57oKsTy2znflbDqdycphK61Ifq30Ln54WgHNvFDl76caRPDU8FimxNGlLAnb
GNWzMejH4thv7SA2Pw+of6lgZLsq+UT7WrGYcAYAVt1PFftZSXI1XgRd3b0Kv9EvrInoEZB965o8
cjQYA5DncQF/TWX3nrdXLjueaLrWHyNgR2wFuNKSjFgvior3T9PDx4iKi++1YYFW4SchwJkja/1/
5tHGyDlfPuHIS47Mj/gETwIDiBbEF+BnDpl2xyiLSQwLAxNd/da5yIrHrgC4GWOYs3U8CKvfTpcc
Y8NKDhpEd/pYqec6+xK3MC/nFJTcrjrEPv3RJDHT1s1R/lVHBLYLkTalmK/zcBuwlAZb/F3mjo0o
LFUVUpOrTA4/KYnxzSaz/yms0Kn/sNVzwtfC6WjcXuc0fgkLZsuy7fBgEBbWkVqlFSIlOKYQoGrc
0oc/NBH0HCwzGYEHuSNcMP3hbUMjCdefD1YSzPo6wDBtHrCuiM8++lZY8Fq8Qd5gGrAnRx0IAQqq
onEhZLZgqdEtLbRCbY6SyMwHBf5GnYMEdtlsxwBCuQZnwSdhxBHejKEa+YWUVIi3DwSE1FF4GNff
KkS3mDF/jXtEZ5kGdF9baYzkxZGGSgVjo61khSXjwlUbj2th1E5atNw73c0J3mxZrj949bOpO1gZ
i5mQY0VF97WYtM43Xhgv2mhJXW7H/n6TY13AzNqed2a63+Qcj0o3hauZWdgS6+R/bWYAFIO+RErl
Ne9D3vup2xG5wGflTJ98AcUGyfjU8f5rSWY7nDWQvSqu9oznvasyU2z9qjSCKxOIntYktODT7Skp
GGc0nNY70qFO4+b6PKbuO4+5iRSHqbMWuLHF1w4iDku8d+HvnCagqKsfoNOl0NdVo1+nj5qj+MGU
mp/YKjKitTCy7I26e+Fmev1tIyjQozUFKTh0LgX5C6Atou6ygjAfrZNm/9HdWJD3XDhJ3NNfbHNp
HNRDkxeFg2qTR5On8KR4h296FuC4fJm0afK3IbHqisgJ2fmGEgxTmVvEph3kFlJ0k1FmqsQb3abU
5YRLbCReoYTIwQ2k1XZ9DSbCaDkCFcS5R8VSZaXBzTr9yqSDSgMZUVUakhGfwtGZ/ojg3ybAqLeX
D8s/G4/WZ+KLzk1Y/J/ovsl7hpDDkiYeEBuZui+e/8Pa0IGZfIOqTsubkd3sQLUQXJMmojjMD8aO
Ak5PWunngcGLs4RlLIlHJQEOsaAppJmRDzsVibkwPPeZL8S4RW8n93+ZpIZmFppBg17FUhqBHhcg
r6XwfN4cdPU5ZcvB14OU8S5ywI5ZyB9zqXjQiESgD9zI3jM6+7mLNjFGTgpRsQ8SCdbmrhJpSe9B
193qZjxVZBttzsJ0iglxl1RqUl20mH8NbSB3Vx3qDO+H8eDa40iOVzK2ExCM83byQy2GafYo6uOr
iDK6Axn4Sd2LIJoytoBuAJ4+zx4Ags5sYu4IxUCZaN8MhtCspXCGfYRNTgDdXIhAl7hDSb6vANFX
FBb4PpIHRjByACXwYCK/hreQcxvjC1B6zrfZ5Ll4Ry1OOA5nyFzGWGBcGAsN2Culxfma/WVbQpfY
w8W9wMahny7VAVw+VX++6UEhPgNuoJg9RHk7pzNlzuaT9RT7c2VYI23s3IoeYnnFPCug2xLuhit/
7Jls4WCNuTdOBhHlGldw2QwEoaVw2RwLsk6e4j04b4Hyp14isPqfOeJy5IWbijQx8Hv4lmX83xkr
1R4ZS9dzsb0orv+1lwlgU3k8qJ0IhCeXM5VNOWS/IlfUI5jw8i7H0YBQZfc2YIkPTDXw2HdWCgTf
GlBg0zbiDkMkbEcKVTz6Ep8ZESOLcRRNB+sb5xKSnh2Hc3a2tYE5ymIAsek2u2yOetPdWtvlRnNS
M9ztZXUWi7yhRNf496HSfb2qD8QR6d3QM4q2n3mWzn1mbrdIM0N9tJL8gcdFSmToFVks9B3RaUsk
BrwwJuSp6nghoMGhaxIAaOyzV0rxHMWeJrC2MQEGLDWqorJ1I9WYDf1rVUYqc4SS6kFxgzscDIL+
I8tqIZ4bX0TZ9iCwD4OPuXts0bUSSFPdMqhuhb9vDz+AnH9yofVTl4ahNuKFeqPBVfOfV+T2sQla
UVr4TowOsSrOSmCD1mvNuQ3WXxX3o7ZkzIwa7hSajP8i02x84YT6E5dHSwJXTi1dMr45WddxmTGP
14pi3QFsXitDZaLIMG1sxupOOVmmZHH3wFLFjMaEPxsX/5ChHc45E8PeMgOpZZGndnkr0FNL6Xjh
BV2ypw6YOVVo8LKS2oYWwdzT+64hftNcURaCBsrfH6VKNevCgFL5N0AUeoog7AtU6UJhhzTiu1+M
PLLypDrrhw+r25bssN0eOkBCocTYl4x1BoQLbULtb0516RuyJPdM+2oykPFN8SKOXYvQQDH8uyhN
UcCybXqvEn+/OVB46kOmDF5Z3blIL1/3SiQnv1snb1cva5wAa4jlJjFUioM9YlmrjxzsgSRunrfi
i4u/LVbmN9XTyn1S1mlkD/mRL7A51Z7pbQb15LVn/HQ6jCn4OTVj8UloVADddIt7lCiKQcA+T8bZ
VuX1zRs2hDRlDCgVEgToaEgH7E+zTl4UpxEkcg4ZSUDF5XIIjWPF6I2tPTv0cEK+i4NujSFllJeD
WY6qHqTisJhqIROpSg7fdDNlLHw9MH9zWy11CNFHYcB9aBp3Th+uM5I//1hL4TQtH0WQ7dOg4wxb
ZpknZpexwVfKl7ItiB1gwwx2eL+klHRt13asLoCnkFKYBgUOZv/favnjCd8ME3lxz/uMZ6RjNuz8
OVoDLsLZk/aXTatD27GPTah7jviSfYlwbQxeaH9Q3MVlMp4VGVPibBwr00kxTB2Q0sWXNqbkc2UY
+S/YliF8lpvt0GR+guOxmZrr+pG+MTxIQCN4dD91SQs0PD1h6IYstlhiFlW9TgkR1QDBbZ7qfTjI
z1k1bSgXlb3tyA76psRGb8WpzT/JPWmXAf29kkg2rBfI4ocpSLu+cmFU3zwcKku9a06QX7q4M/CA
hZa/CHn1pb9PaiU6aa+epyLLCv5dW32rRqneZTs6KQ2DTUf87n6eSQJQGO+AQXzN7SvVSy3ahgvJ
7/FJdplBnf7tPdW+/52HJnIu/G1Zk8oNB3CzJn3g33bPBwyEAGU/DqQAMRXFsXgSA42cRwvEyXu8
byVf9xEOzajKucu7DoZvp9Ntxej4wzjNwiLmNr99PM9qOWl19KO0dxpr3J6tnyKvhzhVJNMTp2G4
BZ0BmJPtGJmf1V9GZjnDs3w/91kXh78POg+zk8mwpfWymq/0alfl7cnHODsxhUUpCUE6QLkKpdLY
Z6G2nMglvShASx0mQl8YR3qg7oe1eilExgfSx2yPryhd8G4oIHw4Zv2an9dx9IoZxEDq/fr+0D8U
Atrv+HYbxOObMqq3EumOB/eRpRBfPVRXEkumWZnyFlmrhcL6XzfZne0YMtVDVVDrsYvlalQ7UzpX
kvYRjnPmpvM6Cp3mh2Vgv3YYxTqXZ0LeJENd6IPpVusyHOUfgnYTAanclD8SYXY19sNAlRrpG5++
VmVRnFZRL6dJbglxyh2PN9cb76wiU0pdsQz/C1MWE7mFvBjhV/z1BhX+q2FyW0TVlcD4WcmzU0wN
UPMBtwuM6xl0OGeFLx8YnQpwCNId+8d/5r3GObh0hvkfX0zpGZ4H+dOU25A2ALQCXsJQ/mOJgNW1
kPA2YlByDrV7fT4Blwzz7QJYp3T47O0LOjzwfb4Ogt4b35FitZAOe/5TvDHpOJEXvW4PMCSro9Zr
r1/Rk6qaoSpm2eAvoW57y98/JnJyV3NENW/LlMTMXqPVu1KVHc89pfEcgFFmDy0z6fRG2FAL4TOM
cQw9ZztEJILHaRbCF5shmbQYC9z3OQsGD0H0++j59TOvp7jPjKxnw0otTxpBghl2OTvmdJYalpl1
B/7131Yp/5kebhEmPQU+BmAIE5FVb7/sAy5XP9uoOvU0d44MRMLvxJeh20Qr1Fy0GV1oq6EIGs67
uJR6ndIfO3SOLFLX4GPEQbR7w10U7AmVo2HZ9WBAPb3sAtWkjq35TkYAMSIu5Y/m3Qoa5KxfgGO9
e/fM7342c4q65cO4e+BMIB4eLSKpYWSna5YJQwBAF9th6VASRGmp4SabbyLON3ptrZ2aGtM/pBYX
QS0vis8I33SnItCow6a63qfLwIt2acKxLnOo9hNUpnyGhuOw9SP2IIXfr1pTiKcyMShSbyaFnkQi
wmhsIRD4U9kfN0Hpk46h807iPn4hcQU1rt8eirn4lI+o9Ys7kITyW9jG5hZPiYM6rB9zkSqWcjwe
MwCFIQ34fVOA2TUGl2paTdhF7MK+pzz9AEameUBIXFRVQwzLj4KRT5CT9EIbGRuBTiPCACkIaQjo
ngsqoKcpUvsX6a4ZF830RdIgC/b9BIc9AH+WJWc1cX+FjKY3dPcMASFYDAmmZN7SfurzoDphfTlv
xXgWmeDnm/d+kAAxJ5VaNxTS/TPAK/9LrCq04Y1aR8hXnJY/v9gquIehVNPcyYC92q4LDEy6qOyv
65rh7PSUAvC+eR2ElrGH3gdPUCZWS+ts9BrzPrJqtL2rCNWR1IR532RQ7eo9ja6yW/jd7weFAwTb
rqKv8ChZ3CvTR1rVy1Qymzgt98rPcnBuVeyE2v68oHaGdZb3yWsV/CNWItQZVroTuTKn7CNN4K80
eICH1iVO3VEbgn85us/Texq4pHuj6y+xxhbqw06NFONIzyVBzIQJuy9flamqzSZ4WylOMvug73n7
rLXJX0qe8za8FgMpGLFI/rHjax/kvZWuT24IiojOLp8kVVc9aAm653DoCmYxMaR9BwUNPw9d8U4N
fI1cnmSesqvm/42X+LAaKdAxPsC5FgYHQYHLsLVBADx7UrJfr9FgQPipc82dm5o09ajuLrL1YU2A
yW5rLmHOP5F0ZMRXCgTylltB4YAa2504ZmCrXwLEJCg3w1D3istHtLxqe1pplEXpzTmPMCsHWWx5
PxsOEFW0hbCJkZZvt/jwZOlwupc9XzsWoH7h6UlXZt3OdA+gd57MXtYbk8JduYgppY/h8ZtffYoF
AReSt0jH6rb7Y8M2cBmE+8/2cHJdfUovecFc6TvB9uoe4dpgHZn82G+S5yD4qGMa046oHNQy9VW1
LF2TpxiSES6jfdhpDa+bujNdqftsMzNoQklZCn2gLLppDkOk7qkEpn59qHqasx1VsXQrHZjS6Ezd
MXYcpQsMWVnGGTje/BxQQVOIBPgB/JC2bR5XTs5ijPdC57l70ha+b3WYQuaQsVaj7MxCGUirjBDX
JDpARMGx61HnAfEMMmY/N0BV9hFeAguPFp8XHNrV994ND8xNloLAFUQSDV3GOHYGYCjETNoxXskd
R/AyBn0tOxU9ZDRkAjXsljAfSepoCKDzLfgmeNBgLewgpH9lOZ8RVra5klSVSYVb8bzc6lASqxQH
1EF17IppQBAr63u1FMjmQfVMhZY8diO0yJumHXSPcipgJQLQXpVYfD2Q9w+8E2nl4VYB6ifoEzIv
m6MFbphchJjopeODenKaG6w3+6qAz0zyqM2bvrGSf7Lv+0o+KLX2Ck0Jt5akBNKHw5hInxP+/FG/
Nj1GoUKbsb/6udn2k4+zZKPLAdBCEL0xZfv1OBn5ZaeWO/gbXon+9KajxtGoXC6VO/LrkrQhxm1n
nXebLsFJvf8TJOLPUPbz0xGhP+ggVXaKO0qfNYu1hKDJrJF1zb4PYe84jfKhRjkDQbLqD2c8JQNA
Ha4XBEkWvt8a9mdZrnqEIEgQq4WARefsdX3PugMkV8lJesOxROaTN5kXFsybxUU+5gQrVN6KGbCW
w1ey5s+BA2C0uzLQO+A7NFLloWne8DvofLWfbt7zEXtCPaRY8NemB2nKwOaJLWzc05Fa9yJFB1GS
ZMgmVUFb0yEBNQP8YufU/gzE38aUhGODkNTKVZ+amNbIbkrutjQRISTVVc10Mu3+3cw1VIqZ/J17
iGmHunf8/T9ybOOBp8AIfNzJ5g/5jedKLSoqwGq27zILApwNyf0j9ZvBGJluJVUlIx11RKyMPwZn
ltirZ4oGtWLLee3L3iePqIQbza0opXpOLd1QhwLnyV/BUg9NdXhLH4quM12wHx0Ihx+zv9AsstzN
rUvkQ9WL/ZftfX0iaQ+BxdcwNTLPYAIXewj4gzAFHjq/x4jyLRdeqOHr/R7eEYu+hR8LEB67cDKq
CpeZu19CZaxZLcnAWenyZIJMlhhRSeH5FLe/04v52uYfh0Dv9ybwOKy3gKRAF593n4Km1QOlss8V
wotgTuw+mDL4DR+Ekse5jqUbj+n3psECN6OQUgeEdVzgaWkO4tr2tJkeb9JVcuEakvrF52LHvWH8
9tBDbN8gUt/ffh5B549js5OGpUr/BGnkjKoHsNHWwzLw+9eS+/s15iSVZuZkkZ45V4Wev04Voxjf
+t63PjslpUBXi4690IFgsylLhZ4D2yaPwovYG1lzJlbATnToxgSMXtjYtabzDKE5eZuOSHwj7SH8
4LKODzqWy4SiKzOtXD/b43lWRbMlhOCcmu3tZL8zP14f9wGIOvJ2JWDR/aQXn5XMubGQ7UGNvW0p
p0cfhUu+RO5PTkVmn1obhernqaE+nefGh9xZto3b52jbj2MaXblYxS7OhGXgc3sOWZi7YDFdD2Wo
SnXGAwWDC2M9n7gikoWqsp7wMXu/1HiwWg6buIvemZ8s4QAKB2FANT4Z/VO30WzS2ETXWacX1PvE
d1NUU07GIO/f/+qcfmJphQ/ydg1Rwj9SPy115QcNPKka7EaAAL3Qg1BvGAz8YeW3PswpbP1nzAQ1
WgydL/KOkrG75V9JCF3ckCHdSI/+Ny6tgwHVgkcwxgWpeAQeyb5lRTwiORXrH3vXKDHgY2dEhEdf
J/DAHJRdhfxLo8uiISQTWZ1Hi2RwjWjWJDVLOsHobszHKMHmliCciAIkRf6Yk3cci/AjPMUoOZ8S
gNkoj+vNBjfYO5NxgNQWsD6NaOtRXD+Bs1SWgsF4pWevC1zuuCNpf9GJvzk0Iy+R6MD4j7ayVO4s
+7Z1O+Gf5fY8cD7QQbRfk0znLrHSyIfAaeVzqs9G+F3/FmrzlNKtzbHk29SXTtPcnyWDxR1AHzQ7
tmaxy2ahCJUI29//4JAVuWgRakKTnDaG2Sy8MLAooFBz1GMtEEdXGr7lqts0oLxPbfZGkFufwM9k
qwUnX2UG6DTX0HIqBAh3IMr8O3mHGN/qlRnA5EHKwN8/pAGhnHRTKZuSrn1dZzTagJVYhtQvZLzq
taE0MlmZ4fERAykwo9LbWfxUyk6fqkruDVWuzKsAt9Iifx0wlVlDG50hpnfIIAcapd9c6Tj6JE6F
+RdUoSv2Wla/JLrHnxp3NmLQSTSHP8z2UfhUqZ4/wgcAZeANzWOBgQeSF5UoWaQSsgm1xh8flyVr
1+TP5WAM5pHzd41gNnbMfzRdtZozjcY9xyLkImAIHFNU9l4ROvjoeyeGXVaeEbsv4Z8w4VW8NMqy
SRaFzAl/uXf3AWJuEUQeOMEtcLTsQQ3ADk+3vofrZwZYqQcfm5myZoOyWCbvMqj9XlmUZK98j7CB
8K1XM/GDaV9A4seT5tKDCbRAqdFQ2QWUsLbdruEC6I6T1DjmiyR2swFBfee/onlBfCqn7GZhAZR9
XmmcrpIGHr+u3SLgKDk9sBKfMVge+6BkLUDITm1dlO8GhqCS76umoYIUagdSWkVf88ubI6ke39g8
Su/UyOZNkaHexcpZC71BbAzdbMRBOyKq9TCzx2Qv/kELBrLIg0hs5CqYndfPCmumZKEv+Fec0zSy
fyCDHmDwsb7wPqgVQoyMixBat4Xup+QSc1N6+Jwid7kxSpcv+bQKWo78xDaQ9OUWEayinDSabbVq
hpi0Pz9h3vL0eP8UK3CZv7k6ARv3yOYGeURrvDqJv5PuRktiLHXB/kMgojFCUikDrcM0zl+Zp4Ez
jNv9AtzQf1kP2KoPnPBstfItyVFx3mr1GAfRQw6S5hUB+iyliRRsLZjEo0pOOOR0cZcBehPESldH
X8p0xMduELgBIZyD6Qt4U+4vBDtwLMHnola7pdk6uzMru4Pag+JFppYjIFLsHYrsZajI50oMYefU
r79PYlLtTwCXM0Llrd5lfxgjY6s33JwhblFDPnmCO94/rZYRa54108H0LYbaPveev40zWGkk81BW
u5rpK2nIXDUdRfEJfp4qVPbs5FZlMBUb1ohhzRus3IOdLj8zsRyt3zXWKEewp1BmTN5IMRQI3Pnx
1BjdhXDdVQw0o2zT63lkJtwWT6wX37jODXMLxwvE1EJ2np90+mmVuNbD141EOK8AUuNQXgU6dcq5
I2wem1xWVIVAEdhR3ZbDaA2k91VcFuvbwNpLhQFWQlWZenc4BGhz83IPhPW8tyJLA7Y9B/Tinfa7
6JEOvB9MYj4NqZ65WohyyEHmo27CwujgCikhT0CG7C3td5Rl6x1eNlQkObCj++Vy9K3yzdKHhFCJ
kVHly+86dvd9ixOWLBOKA+fHds547e/yCfb6a+iGocg/F9eTVxolDbZglga+o5UEhcvmXfYKAyRy
/byTWb/Nh+nEWAj6BUFRyXI8Eygu64Cw3LhxqlkyDXFw7+FlYpcNcwwuLyCboOfefi3JQNoLOa7y
1jddfN3CTXaCDQY8km9hAidobholcZZBXVsZsmVrUD+VYG5z0AGjoO62te6iCmcP0RTrlLV+NCsi
qs4lrRt8eGuyoYxE3MwFHuHKazW+whA7+LBgyk3aSz3nW5HcuO+YmCNgAr9ckPKYMOyr0ij/oD0m
o7uMkonqUeBPt9cHKzVs8GcPDBRM0/QyNsa7KOiSMO5+ZuxNX/fZAHiEZm8ah20iANLMdh/nMz6R
L3Ja0qh50qSBX0aqs5c4MyYo5hWgzMTnRVvyo6993mApHD+fjMeCz8zo0XMmDrOulzUgp/ffes23
N0+CSNahYwFwbP4t58ExcxqbGEStyLxD+nThP3tc21d9GJ2WOIH35BmigK9d6EyXSdLycOWKYJRY
pCE9845lkSWe8ViuTBfBz+I/ukRsWzxx4mTrBci92j7RNNJoFl5SlkG/t64Z++18duyWXvNtmGYf
y/jt+uLGitD+jt1bgp9BKhJfAgXfbT6SFfnvPv+ZYJ54vGkPEYm1zXa5u8Pcgl6K2eA7xs+0pslp
kpMnE2KJ05/Ky64voBoTqQWHWgIkTh8A5v4sOler/tkl8wcQylLkNWRFv00Ex+F6Uw8rpBE1xlNZ
ofwCHyidTUt8J9Lw9a9hfVIY/Aeagtw36siYrK/Yuc/MdGheRLAnxAO2wUmdMSaLLDPaVn1PNvcy
U4TisHKt2f21mO5PtHKUUYhQeelQe0evu6LEGTaUuRLbxc56TuLN9j52jPCFCOcKsl5CsdRZV1jL
9Tds9fORgXeqYiRQr1WrILyHcxqmYzXdm1gtkkiSOmwFtp+XlvK0ut7TqiF63opm+ZDRvYMyKNQB
dixZ2bno8SwsSrfm3v0kFVUrYdE4/KpMUlgwLsEuoVFhf8a47Qsmdd3I5sF/KDd+7A37vtMsC1wm
GOio9ru9IXTUewBpWuNV7gYSVehJysTHqvdt9P1O8eeWiHzvAlFUsnu3OtMjBSuAyBkdbwqnCaRQ
0AFOsBG0MWr2sYrhFzW7Gp4i0OWNuKao6qC2L22BDIQ6U1+4i8vc8JfliMQl6Nv+4H7pTbtFl3P+
dEjMARgwDN3lNZz8VQJ1V0hsb79r7PmEs6PiUPGTI6MusW2X1IsxJgdAWzaRp/kslJW1+3jCdzbT
WCJJCTTSSMzYyr6c51l4YuLCrlBopdpoSdJuZRg07YO3WL+Oj+bu64TbDSSVK5njTnQ9b/MIzgoD
1qq6Yxni+JzkP4JDg0elamBM8jQMcXHnql6MBzgyx5VgSA6gKhiD3kVOtS15IsRQs5/IWl+EGPNT
tupfX4SMEPBgz8ACNODlceRluV5j2T3VJLK45Nqt47syt/TJtY4wM5d2jpPBASl8l2BPLK5hPIBb
9zZbaEET8ZAJJoHvTkHe+NBG6tgmiwaJ9Utt0W10oGJz+z6fp7nxBY/rBnvug7wKsK/Qd492dbEK
W7d/ossSD3871UiHaxzj06kp4NCy47k0ziEIq48FfkTsgvY3iLbM8KHXoR6WCH4wsuUlbdw/MGZA
ocisA06KrARht8VQA5tlh5wHejPnXA32H7K54+avBus9QZbxWfsJjtRcSmZZDtuvw5OEwmoNIKIn
CcR23eKyNP32H+T9qOYYid6EEn2rbORBaux3OEkW0sZ8O/2zGmGmQfGRjGfs9TPbLg34f0YK4KMN
mJZAYYSqz3FyMFDt39PGSltfKQPHmvAC94mfiA1c5KHtKU7t6cXkBjXZuWjo61EnIzj19BCqgpmw
k4u8q20wSCYdMQTA6QouSny5oqkKdkL88u50O4neup0raZwjVUk0sp4vxLP5udsd/vLwhfXXNZyx
xxiwdqZU4QHQmySuL/mkApLHdOXAuGnkztrSkwHH9YIFfirprZMey305KhEbfyZkxLzt4TpbMyVm
H0OXlqeH/QOsTv8SylzC3KpdJbDIEdI17jYN3mMCOGwoMY8juFysRR+ivRMYrp30LyFI/zIP34NZ
76ixN+yhTmqOfyYJnho3qgy1UmfeOTNg9+SjBhqa2kWiLMsF8xhppmBxTL+jezhGyfQcP/KVu30V
qZZkMhDCzOD/PqgVZVEa+p7TrVjbOnhNSuehLDognNBSVXMzjnQx0UVuV/vGxzlnIPmOvdbQ5la4
QHlzJdCPDKwKY2jznxFCTdRfkv8REobM5k8fsQOcxdqopUArpITKR58yQ2ye7KCcNQGul50evovI
FPkQuJcMelZreGvJVr8voAA3W5Rf7vWZlF+vkOhd/UjTvXbs8Ns0pxQqi+Rfi2Vl6ed0QVaBYKeN
TgeOgzpivPTjs2yBsuqjzunA1anBvFpVbWmps4AaZRF7FmyILbT5wnnWM3FjxuoEmL3bqDg2Wtmy
i8EG5UxkiMhaQCSly8iz5BgeuBvh+tM1DSlVEaT3sdFmhBJh+Wn6dUyoW4BLNx83N72uH3GrUnm4
CWCH08FnLabrgZ68bYQrU91XseyH3aLa1VayUptIoJcDQZefwuWW4O9gJNOpbdf4cnVIPt4QZM1z
lRX/792VHDEpUqUHm3mM8iKXqZIFnBmYAPQM6OhJPDMsLqv+cdo9XuBX5fmoEdpWydGhnJhzhl9Y
50WSpZc92zsvYE8M93/CKlhwKMEiNXam4awweRlR7dRvo9E76QQ2rRiN5xC96OfmTj1xaGw0zLUw
X1XjpC1UhI6yYz2xZt3rkWiwMJhP1Ig7HYu/hoVszBmSnJ2KWp74ihZ875lD9uHC5B54/DBSZdpY
BcDBFTOMFoV5tqRChd8Uyvw+9ZhxzgWbJgHhZOyyqGyDxamEmd9Ufxq+xiVu6aBBHYrMY0gsbVic
3xMgMXuHK2PFXX/5jU79nEK6PUZeKuqmQPJHE84tmhhE2maFdhIc4LLrJPDUSspSwkArvNR0DF3d
Myy027U1fhBOVat6tVJQSS7tLlsr2MF+oU1AL8B2QDnMSLmKL40EV/POzq8Uf47UjS2gqJw8SE3/
CxWGxCumxk+gmXgE8oB+6mwahTW2FRlK3Z/MmbHqa4v8l4xGXaGry8tJAvGmYAT8JSDDQbfcoei2
GUBUfe5OuJPxFElz8EI8CYbb5D1/VfFNA3zKnL1eXVcppqaHhtaauviu5Q5QVt7xH8KGKCZyobaF
pCZ+neb4yx/BoTp8e9qdAp02H9/DID1NJ+cYlsNlcgUWCYE9xWYj1+ZjtuJ2IanpwTv0uXCrrASp
A8bWq7AnFKMcfAyyfYfx60LjOADyocfW4ty0KY4Fachf5bMkKjyL+mapWs3jKajoCqc/icqmztMl
B2PUoCHlkJHVCyy+22mnJ3VUh9Tgwqoz6Dmvy87mEh9KK91SQ3sLUL79XqvWWXqudAd+TU2nIj23
r3JqDGtWxdZ+d6USueWEoH6xh4AeJGk4aT/vmasFtSPy4/F/acXZt/BDqPFqBJQLA+rP8n+dRBMf
2KcjG0WF7R+8bjgwDnCmYJcZGjo3QS62+sQCtg6FxiYLPSVLh34DxISc5BxKVco0idWcBIls1Gxr
0xMa2tH8La0hPZ+nrijkomJZozVjGmavRMpdYjNNb+4YviwOsOo299At1qhlLyRBAuEiTgdiE7re
ewdPKvuMiROK28s/lWlozJ3SybR4ZNG4dQACgtH3W7v3ipKJB+Ap1k3gLWM1h4rsJibZarwQbwjW
h/TuR7METqclDkhwQ8jQyxO39X8rehTrljaHq0x5b5Uw4KeOymkdYzkHloMEJu7ojnjtOMtGI7vA
00HMRw7hUphCQ3row7uqS9/ohHJrxEPFIzM8AgrB/eVoVwrfqjuq7/NFHeMwqnfAykbDUizvJtWQ
LG0Hz7rmMR+bzwetayschBo+JksG4etFPb7VHA2X0wQ8EJGTIogBAOUxaI5n6WTegYVLNRH1HrXN
IyBD96PNIqcI3n2jm2+3AdxRntxZ06JuY9wbUbWLFw3nFP4L26yDPIOc31UbFfmuhqjSu9dO5i8i
5AH/ZF1KPKKav9LxYD4xdp74eIm5RGB8eMAfnulGyKfYsKwSAITor3fN6D59yhUVVwF9rTrHzCA3
XZ1wL4PGDNNa7nOLg8FTkrYwBi+/Dn5BmgaG8tqvZ79dnbjEwyMDK94wbA+aiy/snrns7vfnrn9T
MGLHoZJWRFyoXjWmv6ckA7MPJpRPA04SiRDpCBsWKSA6FFX6vw4k9yxbV0RDJLflFD11TPZU2alz
n/DJOMI+1QJ2NbqWYda89Vy+JsiPo56HgjkqtoUTVqht5kHSbHGAXr3MYw8Hj++X2CooCjfuSVzZ
gM/Ds7jpRaC6yEsMhBDCkuomv7qOMnbjxRqj+l3J6Rp2bZ0aryf/1yMAmJwNS73kc2xh0RNyBfPc
VebPOTVWEOvEChjDkI+emUckJIqcc7iLb3BmAiljm/6fJ0tSKQCTzMg+pdUZyPpEPjlwSascX53a
zbfl3WvcJVETDIoR1uYY9p9rMkiYjvE+5SEdw5xLubs1y45Fo8MN4iFQpvSHeGQlNNLP5ejip8Cy
5IKo0qoT7bmoOiPq3g4D2K6vcIEBb3AAz+HdG8mzsXyW10B65tCUBG3zXaMVYkGb3bZw+75nbHWJ
et/3IHfFOw+2NSu3huPfDPzUIQF8efZAxlC9A2xN7QhhH99T7SGQOvJ83+4uTWUQ1B/9n+vIu7U/
lXKQ6LNgpCgvdw6PyT4Oc2KJMGHcnBfSe5KWMItKcK8qa9k6Etb/OzmyyYo5l/UfMarGYWLLPSzg
s/OnMtmc3eWNmJ+OYrV3g/5hKSJV/S+Bsl29y88zSddLA8IFpq1rXn9UPJo+RGR5Pom34AF66dUn
kAP3R9fHRF8O2cz/SVEWG0toaaW6aLqYZBo9NQ+QzERJGk8ugfxgTOnkS+xprlYDKberDksBouNO
V6vpTe+ER4TlW5eDe1ZNfdAOD3B325aTpoM4GZAjBjLtPXbjjhnz2D1xl1YRY/CJU3kcN77exd6Z
5MbLPEQBCK5D+d9OB3R823JRkHh10Q/KOt1ny0onqJ3zKtkdshCp5xxDCDpSEnyLzoBi6Xw9KkQt
Pbxb1cg6J/P+G58+VJ8owazYC2XY2UntVEiq6OZxcjaXlqAyLHh8g8dldWwp2msgVEIjBtWPdE+y
gho3r/y+k8TQV0nv1dqSgd81IGBSWsRyYvVzyhVzCYyy9OmhFs84DWMlDPzog73ePGJ050KjF1LR
wkScTSZx5bUuqFEg1fQP6b7uUDHbXM+EyHSbXnOjP5L9bSVsSmYcDr+KKwDH3+sYa5WUpnXriMYc
+ZwFSkAMCG7AKXbvgNdayHrYBE115ivqdXAZuzDKdyCqYnRte7hyObhbczVvjCrYLxThivGsrzEs
m8ebwNQL0Dchr9fdFnUrc3bv9+WbRn24CO7mXkAthah0rQIa3Cy7K9tcCsWJMy3P6mEQ0rmLZJck
S994IDP4XTW7j2ASKs9+2uYw+WgCI/cta3diFYryJmE629CFkNUyvsSiVCEutT1CAHANHEJC/Mr0
/asAOeALEgC3p3W+oQ2JmzjeVwofJ6z+QTzsImoXVzPKsfJbpzXvMtqaZD+0WXXfg19ZOtLK5ivl
sBY7DtCabNp5ceI0u1V9zqddIylB8Ex8GglBNgaRI379i/Ktj7mGslV15EHPstZOjTS4hiWH4bux
A5MaLCznSOf+2v9Lq1LkzrWfanG8/+Hu9My1r+KiFI3PZ97DTzn5DLbrmWajdS6OtrOweh5s1IkH
Xc2IH2H7N3i0EUBt+avUjSCoJiwMzKxCar3c0WzgZwoG7uF0MDFiNPwb6E90zuxmdORQiupEAGQz
2XY+SD8fPHLRFpA/fjafFFbKShTnfm05uGArFeVvgVaEyY5KISCjgt2e1+MbDFPQXRoqFd6f+E+C
+fhCNk0wJMTmxboPouJ6cq6jvkoJw31hnep7BkNkmxKD6zG4mwOkyLuNq1YhkDJpHqodLvZcOrkP
9/cAbH5LuqpVJpKeLbveXEZNFUYAAvCuUj+lqRgwnNa8YGwqYUjm5xrKGJj4B5pG23bKDP+cdmwZ
+bPIDuen4w2dZLJvCljNvnmfjJTh/MCeh2MjJB8dr61a13dvT6iREbPHIUwv0OzR84287S5aNGhn
QxOKXtFUSBvq9e/qvcRwxmqIDWJzbRMCzRt672DG/QcH1L0eUNDCY/ru0FNfwLruTq8wnl0WDMjh
X+qTPjuUMR8DBZ2tXbsuWrHfbjQf5sUiAm835nC4tWGcXt2QeHNVCc4NwQY0KO6go8RKHpShGuDi
yhxuHVw4WN7nR+GPjkcf91W22Tn/ZJPHb06C5mYgLGA1OMGuFYZBb66XE15P6LWBl8Xi4VHFFxUs
2jB+JXAi11utXsC84FZpI9Ti54lcU19lEgm4Msbq7jA2m+jbdCqthlcoZGqPDJJt6NccyRHe9B3A
c8VqfdeHLLwVvWpgoxoujb744X/zT83fdIJheHmFhj6lO66htl+JyAKBYyHGMn8PlJzsxuph7rkd
pw1V0OmIhPIa71smktglyhjHB5HyqHahspRxqKvv1gO+YlZ7b3vgMe1mAnigjbctYNUmWu50H7Mi
Tt8Q4d+aTdu2Rzq088l45SD93WWA6B5otMx0cS0tkKKRFOIUSvxZHy3e9+1caZn5daobnvv9vLDt
5OZMmwrdyJjgBnSTPC5DUr2CJQnbEn1KWRb8O4Q7wZyTcP9ePYtj4Gq5m38VM3pWFRQZEgMwMWv0
sxCvnBVfT2ARJN6IBInenEegLyOKXb9Nlzon4MkGSYW7fRKEsTgWW6Vz64jB9vBV6sEv/5rOgrog
fSMUfY6e3ivg2jTm67DQD2udOSV0bAzymqN+kkVXBGE8u5nnuQ42u3kteAdX+o0irS4qwm7fTCOX
uY9/Y5keNFo3X0+cviIQ15hmOH6t533pBCh3KAqYwPoZhonAVeHA7wTeEEIUiM48sDvI2wxorO+l
O0V0I4AkjJfDKzf5SI0Lfqo4+ugk76HyqGNJwr7rTruK6PkTWgKmRg38BPc6h8GOuPzelCTd6Jtz
Q8QYeJa7KCCNBwFoj4kyqSXH/UJMXTPLjoNiQjA9Me4nFTlJYnoimHxkyyeFjAve9ida1upG7gCa
ALbZFemXEbduF1WPnejg5YCvkUoK1LQt3vjN4wsva0U2lzkJz+0jMILK9HjnTVDxktpvGYADx5R0
txuW91y8bUDB3KdnZjyI4brCvA+FM/G3uKOybWcSb/cUkzeT5gQAYj/plLDTjbxOsOL5xcN7NBlu
5ETm4D5Vp6EA+vJbB2iFVpojl7AuScWWegIQ4rrEbe7GZN5YypRMcg3M4GPcmWqveDh+JJgrPAa0
pFzhQ6xewyfafQTFikA8bee1CkKcz1NnZAZEqgX5rLOG/gnqxy7fgWokzJQHXjRzUAJU7BZR9eGZ
aMHoB8thANCgnIPEgZOekmprD9evouglulNupkEMk7BoZCry9aOEOomkvxDVdj3cTLwDS7IHbV7j
DLtTgib+aBTSG/Nv3pgF5Y80u3ln7emJS1teVaxiyC/tBUMx7Q47pCuuPsDOaR3L6yzZxWikaX6F
29ZexmcG2JrWU4niPAODbkBm1A2hFHaifBfC/EMLhZnJ5B6Cra99XS2gR4Iw4TYeIVOqXH88X5aT
5P3mbrEdCE6VAR0q+LYxZ5yQK2AxpGVSBsyoU/ZRbstjcV15W94bzwqCg1fHc7iO249bzqARr3bv
zPOIIciV8mvvH/jjMO4aqOFdF682sC5UhFysHIJGI8XiMOW1TtJrzavb1gUNU16psKj07SUkYvSK
edquKfQhp/pHE/IE2SiKRFh5jLOsJCR1+LTLmkdAFlNtGQ1q1Jgp0H/4cOgTQtdIeH+ldHWNPCBF
EJBPFolYbYkIzGJVds1WmaG/TZz5P4Pm7W1+sFc7O0PIVEWHDhQD7xTTXrcrn2AEgyZPv4Rw4cSI
zOE28aolsD8sMUZWBoIxmXfrEBleD8diR8pjeEIbTJbdoXzGGLtlrqimVYNTSlRr6wfcbzO2QBGd
4+oXqjFNreLQe2Bo7TrC+mT1fP+OfidRmhHMZRRo5PbZDjFzsX07njO91SYyB/wztNJxya9ifhLs
ytGddwtKl0R+XEx3/jZ3/UDoG0T67lt+aEslnekSsLCNVlPKEuMyZFXnps6LeWgnKNg2jeuBEzbS
13mMRjmFqbIXwuw51Kd8UYpJQpsbWAfSsTt3OL6mINZwMEIhYHbUWKHRgv/kXcfasl4Xvtotdodp
9icsdgNsI+3x20ZPJ5BkkTLYdzAJeZ7Unj8kd2OY6JIoycX6Z0pon9++hBsRaZNPq0rxa3kNxZOk
miUSRY/DycPc17r5wvuz3NdDGvngBvjXVPVamIS+ibNAh+4Q6u9fekhxRtEqF18YZqMiGRwJkPrO
rqkKmH60zOGdl2dMsbun0/NOPexD+jULFeWi1uL3q/VgAknw93IWrr41+g8/gQyRBNmvgkcI7uHT
bsvOqsevK8wVowzYXPg6oSA2pAk8uXmqY8aqmE67Q8W3jjOn9/DBTmubw+xfGfwA6JcEFyy2uVDs
j28pdC6w1MYWj0haxUukdBf3wh96lhUL6oA+PvPEyplt4MIppuosnAGktExzPSZak9+9uYqrJqlS
GMl8sLFlpyOkIzEx6fQMJSUuxQ2KPFKxFq8+0m7dB62G5Pl48DdkrfiTeVl/8iuoO92ZZ8eI8X1P
blJp3twK88lyyYsogwkPyvEEdSzISmUhkVPX4l5c3b1SqafnerNmkDaLbH0F6EIpDVcGVEgSOak7
qd98f/pnJzU+OwJN/Kg0Fpa8JGN0cHF7Bz9Aiyzz5hMq9fpwEqblRkh1P1gDIhy7DdrVhHRNEBd9
4JmBLB/m2Zba7YkU7DsbDfJORqLdyOB6Hidp0se69KBETXk8uB6ZysyybmQ5vj6p0Zc8F4jehW0g
afNaZm91FLpc3Z3nJJ0ZmRZbT41fyT9JXh+KDlEC9vpOKHy0S8W9dYZc50jHSrukVFnOpPOl5MCm
m7TTtZwbBAUVLIzL2Nw957BuMBxTaZE8qYQXCFXwiwebN1uGEzsASwj1zyIS3+WeGhySsSIUhxCs
zwxgV2agSNYpM6yahP2jLyvWJDEZTL9ZF10aOMWv7zwuOxsy1Mu3s1ZBWif1UYnwYVt4YCg3O03W
im2seRoqB6sKdb2HFDIIBvIVmBvbLaxq5rMVQfVLskMu+dGwoH+J17kcBpQuI0FNTZbSeMHD+8yY
KCcKAsMP8kU5oNHQXP0QRoNxrpJ8aCvFC8TaEHs333c96p6SIyYC1PIzCg2TezwIbn7Hzp55Zb2w
rW7J/XlElHCBqEy/VfGBY7RHIzrLing1MJPTk9H4rz862n1R3xnHe/S+s1zJhyeAHf/dr9tGgZSX
9QGGp75R9Xlr88vW/ulaT2qzc9H9iyeO8Ad9V70neIWDabjcFWv/IQhlH2i8lWUnPZgPHlN60gZk
V4itpkYfJBvAffPapAjeDD6C0E+zyJZV0RcqKU8F5zxKbGFF/hDZ4k7YkBjlaXLq7cMBdOxRqQXz
jsmmSCtPBQT4+4Hb89JprzcPrPa9GK5zHszlFBN+yE2xjqwimojZepNUsfA1UUy/85GJJHHFBQrE
/Ul3/PPIC5hf+ITIuWXFtD1tP9tePnlSEpfJOo2kxsE1a+aep07ihIlzcflDIf867p+6DhXEWdeM
HgoDy7ZGYJ/jG0I8HLeaPvzVvpCACl9+rJyps0Bu/2i/2sR1jbFxMtJwc9w+Y43bS8noH1B5qZMf
v9Yb+rgSjJ2MxVnsLqbPuf0tSB4UdoJs7HH1SPviIXLB8Rhs7sokKV4fxl5lM/x5bhrmMWNhWIB8
5xVaeg/kjWwCHjAMwkXqabDP3LzjUYfiD22CNp78wordyJXK186DyMfBPLq+IcADD1gCamegnFTh
srsEvM21PfnNtcupaYFEARH5XnUuioBMkIVpWQj6pHOLJ6b0UBDgygocHgVlkCTkci7v/hfHKbKI
5/+v3KwxqY6YZw1jj4Vbwngm1z73DLUAwxZDIcCKRTHHel38LaE2aWC3RsK+ZUiMN4uc9035Q7OC
lR9QsWSYku17QbAUWNLlXhIlWsKBFUGcn4crg+T9aN2m0/ViWvmqiemGemgwONDLzn+qNHirey4V
cEJeqDncsEP2K5e2t3IjyYt6yHzuAK1l878aLVUnKh/+c7U9InmRC5NGnIO+oV1SdmX3NjaJip6Y
zZS7buPYiHBKqgZ7RUZyreWjVK+mT6RH5WCbxzjDH+4wu9rbau/KuV9P3VYR+LOtmtU3jMawesxd
He3MDdyJ/H+Qrz/oYzacKuPkRDRD32QlJZRSM1mP5pBtZLkofz7TXN6ZAB69l4lPwx9IZQzKf7qe
keJM6/b/Pcueem9G8spKpBRrl/Rois79iAH3zCp4OWgDY9a/s/lQtJGVfmWv8449VgUjDqGBHcHg
xVModvRXkNzm0bC7YJrRy1CsGjHVOWgshW3fYSs1V9ujKJh6YbY8Zb1UHFoJBi5JRlqoapDO82rg
XbI/NtkuYhRbDrUOrxg530oyBISsjN3rsKPlVdS4WJyO7l4Pstfn2SGc0y9lxnye4C5IAf7Y8Dyx
xr8SHPOIlBXo+PqV2432Lu+eekOYcE970/Zp5QRt4gkCdXGngt2Ax+6252mShmLUXu4+bFSFQ7yE
qY2jr3/OlGdha9FTY2yjgxQ5A2klSK/bywA5paMvBHHS1bWT2grHNkTYJnB7WH5JjWQ+2nxdV2bb
lSYtPauPSzJwxTzROhL1cELO3wTI8aNzUlen1RRqjla3zPh2J88RVlU6Ro9dKRpO/tOnTSotLMvK
ozRkGVN7RP7/wUgoqqQtbHR37opagSoHdZCIcgLoMs/vkmqskiN5dwmnmIYyqGgs0gth7S4ALWmO
dW/2YMCE7oBzFTj9BhOXG0JWvWjzzsugg6wJiFOhpVhQUfrThrcGlulz0fcL+hEp/QYax/sksAPE
XcwQjuOzubIlwGZo0NWehrbSC2gZvxLcWfUIQmMC0XSYgAnxX6Xx4hLeDWAR3n8TLtTcNe6lOlyl
ZtlXwcnxIs/SfFcV2QkcTuzNz6rNpJpFQTshu+KUyMdQHkH8mF4i8GPU/AARNaOrapkRuR5BtfHM
dfSrUi3nelcpZvlmZ5fobYhBZ2s/iKFG/rtXRBrnaEjB1M4uqMK7beCCEfR5xwHmy3kXrx+ypHXX
ONvu0Q/xq/z4BUnWDsZJ+qC1un3n/2roEmzJdcyEQLxsV2ltzaKecYkN4bUR79MBgJGWnJuCE7U1
wk3G38xP46Vc+MKiMHH2JUCtpt2iUYBrhaqCRQ9wAM4OsgtcR9gb1gu0ZRrsoS2Qg1MxykAZTtVH
Dl/Z37tDisaQmbFYyFdoAWtOuL2b8l/lD1RX1kzI/e857CqbF4iBYzbMYcRwTumMrTRXAkUufyTO
tVkr9V60cpkWXBMAhI03vR9w6OCffO2UI5WdunxY5wWX9henwCCQezqISaNEeqz/7CgyXHyfjlbU
XKpObKPnJhQJeNG/t0CfL0VBudW17jFxCZyy1aONu2KBllF7mRF82QMpQ0esD3o0u0XlBTDk9nCa
vZs2o+5/AlcPNqLVKVZkmFXuUiaQhzSqDFQaJNQ+vpAEiWPTwCsW7JpJrtLu3iG0vWXDYrkmljbg
l1iXVB0dm4uBxujanYd3SXroDEP2sP9hX6pjiIxuYsVNBxRE2nXvQNkWmtmrG/u0wHrCPViXOjV6
LgGLq6QUvnJIkHUtijovmX9HjfQ7ZnsNO6cCyrkiNKKJSxz6GXoP7NFICZV/eYEHDlvPMQaGhOam
XziovRE/BClABZFV0TVqtNiLMw60dATvJI7FlUqtbjMiWiuT+VoCj7z/7NeQ644kCcPIJ85DvQzf
cApihiU/ApAUtDfQH/7CvnMIB6LOIk/79seQAs7TfTwU4sWeLMmGmltSCG2Gg/riy6v99XUWgRfU
gFeCvyVhYWdYlYWcYSZeYYFXQbgL9XxLSoT2V013kGKn3nBHFprN8EVuTBKTkpOwO5T48x+Eavhu
FlVgqKCYwIMAyC8xTDmd6FHo1knMnIlsySX3vsWAKC2IYgee2P3kN6revbzaX3As4plYfr0h28OP
TRrmFSo35L5cOJtzgWiDjzmfPll3538OG4qyrfg2a5GVYdjx4GQw5tg+7GW76ciwt/6lthtA/chL
rgj2JWam2BCcwTzPelZCZ4J6tFeg9dJ1LZ0NMYPXHSt2+XsAaEbdx+fvSuhddCTQDYWvvqpuFFnx
a4tlOZakppg3aXFLe6VQnydcwpS6Y4aJFDQCRJ1rGQtNif0hspRJ4QwEIC1I5W2rEncR4pEo+wqZ
SVWjszAUSmziAScYJqHjEMMTtCLPdr18CX0DETMzmoEL5rFAZyoemENoJjOunvFyMkjDAUr8MEwa
yqxuUvMOjSYz3I/o53KbakmqRfb0IXfE1nK/iyq0W8VcfQbhH8ClUJPKJ5Zd0yIHdlnjNL3AqsGb
LXECYXVa1nQiVRfkgnYmQ0cn1w8KR2aF/m8HfvJ8XUtejjLwQAMFZ2B7LwjleenvDAvFvtVEiciO
PzY/TDBw17ZV3GGOtS66ALb3/xk/YsgTrSmf0T1M0aWKQDT0Xofzd2Xf+SmxZFSiO0cS4flOi8my
bRftdj1Oj/KG+9jBaO9fF/FNHgr0GAnt0h2pTllZgxfyaioGUGgnyj4BvvZPDmFdJuRIGkd53Jr2
JLue1MdD/llNcwXTloSYUCWdhieaN8Cb6JXeNpAsV5j9wwNN96HxPh3L+UypK5e4c7YlZBRb1zqR
lIa/BfW+uDmJXArN+XURxgqLf7f6HQuBXJdnMHGiCIT6JhWfisW16pZRBDVjZy9gpjMBTgD7KO18
ArXPXmxIIL+Qp37N6s+t4JZwe6PSNv8Ks/A3JDh8hE2ZX2euorptbMxXUKM3GY5B08jXc7zFheAH
uHb5PC9nqnJc003j7zkSaOt2KMiBSN+579mCpLGhBSfFo35m4OXOtqvn/o9sWHd8fN/449dnmZmT
2+VP8hBJzdoaPRQTwt6Et9hwGVpg+zBo+VIpvhFxNbGOSCNT5nf6E03JnUtbfXHQkKk+tnhc8q2S
AxaErtjA3Vv1meOj2c1qwzhyU4xzUVnpOyktXNsnd2NSi/E0OEsLYkPQ+a2G6O+4Kh01d6evYsZ4
ZTP5db7XVKGlcmbU1W92h+fZ1o6CN1WsJ1hYdrYWQhzy8FBn/4U4so5bYOecdWqnm2kaNEnFLrUA
6ZDIK3R96M0Pt6eLGntSXiH3mKJBGcYp8NxpKFTO5c4CleftdGHSUcuL5jFEym6DYe27OBcI4pfN
R4EayeTh7huw3xmNOgXgmAkID0dAwfKOkOgGsSy9uCs8ROUslGi9MIaf270kK7HSZsyTkuouzVMf
Y2fhDuHumz5IO0yCjuV9kh9xOekCg7cT4ZY9PU8mukGFrytmSxRfPCp0DTvXzEkvROB9AxLIbYoo
k2eeg2v/UlUtNJDQONf3ASq6CREzQhtd3QrWwR95GMueSnwfk05kBP1UWg97ZPa9nLIBqN7oFgCj
S0GLzZi41Usbi1LO9pIAsx3kc4Rg5TBg969QgVpC0S6oPxHCZRjk8Z6Gv2WbTXQzhOFBkKlpUKP8
ebqZBM4U1ATlpevJOqybOr107AsMuJo2kDAfIcDgeW32lCgJFgCnjuNA0HAeMWrs/m8Lrz5qvoCD
g4IpWlTi6xitT7zmC4Ng2lf9EZWyfVmr/rale/pZ50/FCEbjobSWgKlsaku9icmprRGtEOcHKtSo
j/59pfKhuYghio7V9xDBfR4dl7bclNrqd1ZqkdImPi1skZL5e0dUS8I1eTx3H6etjw0G5OSGJAIh
TcpxIqJGAgVfNf4h6PZNMDf4gP6JW4ovApNd7c+qdBED1IMkpYyHyiVsj1hCn6vF2EVlOQ9TnriQ
DbwtwnH96V/UGyuQgs5FSae95f6o4ux7tj3zXQvOsXTc8Pf9nkc+bWBCLhB4wGpYYRo/jidOA5ow
Lb2BadaFBaqTeBIAA5NCBWs23jLlU53wG9HO+sJXylHOvfEjVYAWk+HRKQBSEeeL7XJ2Vikb+w5J
CKV5aUH/xkIJ/0aigi/AYU59H79KGqXJi5N8hMFblwysobisyNbJqxgKSDvKDTjNYw+tNO+WtRIE
YuZYSb58TqPgNK/P/vreE4sIvfXxeXidrBPd41qkvmPai/OfB+/7D7K1Tlnk9qiDtjnWHKFGhZeH
TWQzj9Wc/lFC7p2vv/JTE5ujC+1oJUK78z/hg47cT5/6RVsxfe6kN+umTthmc1BQruxPM0VitLit
bWmaNaXykr3hCmopWJeJHzDwlrWS9HWlVFBVzql0UoN7rLMKBlmeXGSw+eYaS39A/y2tIF7usoOk
Q07BRgT05IWQaIusg+kOjepFNEYLEum8NnlCFSxvITH3YTgitSXxV9fU+w/fphNntR26oDPNrOLw
5gwP5SPwVjVGvmqbMbNo/yhcAsywRv8GHYJ5nVePMRo6NpfJztuq2towpiyQDjkFDPyfxIWBzwZV
I+u92BWXXC05wSTINN2Wfv8QtmOmV8/+RtSqCv8xZcyMj5DN0Am21Ew31T2pRbTvwFNSt4jYhCH7
fmDewBjjQ1Kk0bmanjRodD8So/wTIKq6USeMUJ7lTv9vFwLX1d4en36hRSYdCLeY2mAaklk+/nMT
gZzsWRVcYSU7SZw9rdA7cUmR+7+LKzhdmvRBtgjlh+VDlx10pMI2zSz6MiCLH1pE4bibWbFTjW/4
PT0M0O5RpQ9x+7Ns7p+FOXyZsd4nb2+nnVuFMpqsWZHlxVkUdRYieiNDC31jKQXb9BWxxssPP6oe
SO9BX0Oaa7hANgNzIz04KsMjDnX8bM36EkabZ32N1TonSthRjVGGccDQfJDDcsHdKhlMrsS3H1/K
Rj3I8DlsqY0ccT82GngRYbuOLxsmH/V/A/DwtqWmepMBJHHHfPywYejFC/ocg2OEuRc2clT7lfAm
wfyvrG2TtzEB6sJk5R5lNOleZ6qOCwiwwE5uW/6NpEUsEB2GnBqr7wppckSFsfEWvE52HitauoI6
frTVtODgFVGBMOivtuWsBuHEbUICPKS72tRoMImEsV9KJD0K5L4JFDVF4HAy9yHR6zIKjbmsAJLM
6kEzRog3Or7GjRs1HQJsAiF2XiOZoXKXzTXA02dCI7EdewTcpTTc/nemBWLKFs6TFcekldYEjr+Y
hWyzgK7LAgjFk8+dFpk8Prf0M0O8Lj57dvAccz3iKn67Gv633DIznvd6VypEgRHgNiRVChIZxDK0
1OMFvGK3Nk9uEdJB5/MC+QqqM97yE070jjumtI3218sTDGqPrYhtrvjw2UMcNfEd5zKnPDQdTOtZ
0q0/T3D4dKyy5kiU62Uu0PWM6R1tqn0rNhk/tuyPT6mPrqJGzF3hUyQCmw/pTSymr06em1ACtX7U
/24Kb2Pms1xMTv+fWiod+gMR+YOMzMdNasxGEhZ298QTyVT3vKIcXm/tVr9obaNRYvqpP67UUxL9
FFUGX0ne8mzPX47bQlsvtoPclCVoGELDrycI9uBDFTZ25sfOPT47d5E2XvZugCILcHwmIPDMm0ER
cFciGQO2vBvnfNLdsurvDk4z4VBgFDOXJCyHYVnKBHSPKytjhcLx89Mu/L/EZ9AcIqL6TtRTL1X1
X2RPYIP5Vulzp441W37uh2HUx5qjJDOCQcLhN1pAAR4vQ5rEhRT97qCvTNpOK42khf1ZhGGpwkVe
2/klmzW7K0dhvpWH6RPpHnUi4LWy9cNcBPxgYXOyWp0GwzagQJSfJRBFE83xNoqteScGSqdjW18C
3bnUkXjlIGJUrJUABQYGTwpPvsVrKTts1RntPhPHPUlAc3lJ3noAzha0oJvGLeC+vUonC7wd+RPA
pOr7h2imGLkkcYy9xBOwOOM3AUKytB0t/AkW1c2VwLMLCh/5P+JJeQCAYgJtfYD5e+o/QZOtyJJJ
0k6x/BTnlhR9LDZhdOSywJQy5FNoI/rd1tLGABO8o2ZT3L6i71xiwfMDiU2fCGqZGkjjsqQRkeiU
2GW5X8BexPhUtG+F/qC07pN4ZOlheduZfBqKrtXxnbTjFJl/xn20waH9yVqmw1LhBkGFfPlZslmk
I9fbwWfQhaJfcj7a3/DA5j6Kf43fKJsjLdVbuCDZ2LlJ9bKZrl5rlSg+YJyME9DFvdMV+18Hu+HU
AmGeMftdEViKCiMJLCBH94JwqHEEy2cY9F9Y7VQ25C9ulEy0X4RvdTD7tjvWnW6aGBdv5BrasGRa
4sSlvRYkvr2YOmX0KTB9Lq+yg74SuHYcMSTCeTrZh1J3g2y59ZdWUFG8DgN1B8nImoAEs1l9+oxW
em9Wu/vHCgORD0d5K+DgeyCrxtY1sjcfvFARaFkS31aLU7hmN45NjmYcdFATM5Qbbcm3Fh/XOuT4
qKx5hS4TdNUM9N2j+y1JzmRmjWZ8+dxcu9Zx5Fo6Kn4VnPrtTnZUiKVp6FXM6k9fHD4fzkr4vTAf
jFnsTfjwgaUOjm4J8tAfcnGcKfVbXPjFEHJZJipTssllXYqvzNhRxsJHmQrIY3CdQKM+PtFgYf1M
mKAXq2AjeqWx2bhbg8jdCMrhS+Ab+77n+t96XLimY6CxbMQtXMpi3b6NklRCyEdZwUj3+Jyebu7R
Kl90B0rvGpgP8tI5UdWrZMm/WLk8bDBPio1mLWDmNfUckneuKBCQKlhHh7/IESR6yKS3V10GcDe8
Valys7bBGCKuv3PIQgrPmxoOnVuhLKMtRA1H6yg6tkLIkDXhHwIM6VKd/OlUsGWl3q/MXexszvko
yZKLDgLrF8q7W8hlc45JhJjWXgcajWs/D2k2+ZCIDIGSB7VfC5NcCsEQFCAahy5/uojDN83qSCzk
Ai9rPvFJbwxbsZTUhamWTDC00Bnj09xR00d0f6Q1kl1fpz4ZI6S9QIRYQzJoHUapwAP9OJCf7xKg
5ZCThvM/FNz18sl6s2583imF+sVbFnj+Bb4drPKl2cGShWwiEGhb1x9NMYi+xOMyHSvlF/pA8XIw
MlGCQuwpJF8+BbRmN0iVSCnlInaZZj1AyDCUGQ72GZjD09QVMoiBmDy/vWhliDnzgQikYnro48sp
7Ng0TsNm1h+2hnGCaiR/R32WhEurCXjvwdbtP4TFH1nooDX71Mc//PbZA/Ig7MTQP9BLEMhtYV/a
f5TdWYMRdgMJY8scBWvexTdamIMSzjxRSoJ0FKe1XMgx1QVYHxts9PlVIzYeAyDdjd2YCWPV0l3K
DCabyALIjbP/D1QXrpCMwkQCkjhSEdfaBVdWn14Q60GxUE7oYYnWR5QvC8sMKDqQtWJViH3M6xQZ
58gNFsixaJ+AN58FzpxHvPqhlwFu1GmdwRFy1uDJ0Ac99ZWTgU8lWGYI7TvKwhF4zf/GAS7IPtnZ
jqReFUvTaclTG8JDg6mU1EEJ3+fBhzqpMbIxYT5b3dcNjjHzsH5WP5dF/KIj0IbFUkJgDdPAdww/
axjI9NGAy4yRXSAJQuOmxfIKmMteyboVo5MQboiDweubp+YY4MNbOJETqjfIgwSJQ4bajU551Wgk
lHNyh+MZYWFaCyu8nfhhhczCrov9G1A/9Zk/1lNthKbrmEKahmscPf8g2Fkh3nZ4IwEdVEVK5unx
+j7C60QVT67k5xeZTatGMB3I/L1jKUQD9jhAOtxvd0b3pKBjsjeI0G2XR46XmbQbYMzhluGOcwIn
1kHSLew5kS0LfiBFL9gLqGEfXQHn9w0KoY/Z2GHl2Zx1IcFFlZSWVg6hCTV2+IKZxRs26ZEcwKtM
r+fz4FBCQezsf1Jp83Ycrjl57BrZn8VyNjEbVbAr3LlCW7I6WRjAuOp9ZY97DjpRDoa/MS2f4aXk
SU0EAwbdZo2s0QsBWxTZ9jp+1uOXzghnGbmt6MJd/gEejyJfTFX2miTkyE42EAy2OgwPtHM4NVfD
aUjSxw7+KAsexCgdCy7J0Q1OCLHND16GGcQ/fdntLp8flPvfKJftdAcpdkrOrCn1wL9XJM+tA3V3
R0fbZ8aQdPCzwdl6GcCN4iHFitEoRitMYq58lfvt3Ii0JkxKls2lWmL0EE0d2qQwlcXkFSjVfRU4
dPhWfSO2avrnLt6d8MsGNGgf1UcaZV1Y6K+SYt11Vwbo1RPBSoJBsAxHJ27GcNwLFviKEaJ1MyhT
hUtC5CiMbNQgZlR6JvSxmsX8kV3M4KP2JzrSKGpBm1/7XI6L86JT6EankLq1oUAMM/80Csfj24jt
qZy8xflKzxHwr20MWcNltUUqe2m1Q3P7pGxJvPToLCxdt6KvgNJQVr1fQs5f1KvNNBb5rP9nZ35S
va13OhAkMNBPnropGHQc9gm4DaGiT9sKFAPk8Q9v5r9G3TIdMkvH37BxCO8ASq0qqtL4KHQmWyEK
vsGU/TVJ0zW5kG5fHJ+0lJT4RI4JvPhL29uGH4swKh5Q5Iw3MgT/YHBzxLhlev+54Lsp34bCxLB+
nBV6WvJ7uUmEObz1yvQMjOGiq9KHHoEr5Kk1e2BvzDjKBYRC/kVaAOQhsx6EyEC4vsfg1uxyIrya
ReGy5L+CzxLz+fZGuGrGP77oto39RR/uqpETIK8woa3qibU2m0Pi3SvfVuJTzPtExbiHMle5gnjq
vzJmbTFQX5AOV9GNBU3+mh2HkV9DOdyX1lWwF6qw0Frhi3qHo5tn2PVRl6rKtbQ2ot8LLAH+WJdi
HyPvvGKFnt6pGy1y+WG/SiyreUyOaFIXmuiiZc5VEYZvfU6EBC9iEeLfd5fmjjOykw40PKs1gf6y
th/yJtmG93+aI+OBx66E0LvdleIOYnrYgph0lVVYIHS7iRzJ8z70WRe9HH7yPLWVpucWjSl8aEd2
YRPHvzMaUr6IAJ23cAJItr0IpBXpMtOaIjGZ2pvThPbG9mkSyYa2EPFubEqQDZ0pKxB4ZlqA/x7Q
thklHyOQ+mb1QZWOkwJTj1P+ZYn5x+KUh084dFsKDH/thmYbHLCpPRJIq+9kCDkUZDIopPCnKvZV
yEuVFPQq5vQiiC0GhSyrDIxM8uh/CVzE8RcmAiR5reK3PHCVVdKGiBwKMaU9q70zZHw+B2xwbm4C
IH9WktQQ9abuDo57erhnt9lNfTj+VfDhVvtuYiTZ634fWUsX0hw67FsbVqvtfg3LoQ/hbuafkPsd
DfDHNV1moIlthsWY5bU/C+LZH9ROBXda9h9kNTBWMW47rOsQIjePZkwkXHQYXxkNnPGiU8WokLDu
4KgwYkGMt1AU49Awn5nRUDO6wzoPX0y6GxLiSyb6OU7oJOBfbyohyOddEDdSCay63hIckXUjCq9A
iEH9JooZ45u8yDJxkpv43HTQY72W4zierK7gBKWdtq2IVfORW1mhjs36erikiVmSscE4pxr5QaUB
LCeNPkN+ux5LcuruzScbVeVelZorWJq90FJqpM3rx3VzE1SiJrRdNpi3FOeK0J9FuRnBz0y4WIj0
Ig0pugw6x+DYwR7CnbmPpGiEUD6LPqs7XhqBUfUfdXa7xSiYf7BijnFsAcgUJFnpECQ6OYijv5bO
rgjZFnGWYLUc/E/8Kf+aNq49TkxV2pKjXK4ep22FPb3mjejW/Gx4N+eurXyQkQogu0Ih70tJ1OB3
Y0ccVqhdzVW+AfMI4nsj8I9xqT7bRChw5sR/uVZXzxY3IvBSxPR4/BabMgaKvawEEPymgPTKC0KU
j/PZrImcAhSMRV3BWNsvrVk7OMzTZR+/5XZrY13bzJcDgHs/1y1R+BUmbJhC8Tc3hUkkOo8YhYV7
6jNmJzHsMf3w+Izg83RvCGaphrl8gy7XsSwGbXsfeM1FWh826QLUM1sqk//04bE6LiectSby2jdu
Vmb9kf5IldEX2B1HexAfI4u4+jHqaEVBpR2BUfingWp7QE50O83xZqDE6Vgx6rSxRqlOWMujtQC7
xWmjGyZvjFnfuVqlP/P7d2pR8nw10W1id6vVRrb5n4EQjLGZTjAStx/fm3bhwrVq49+6Bz/Lk8aP
/NZC56LAPw5JLBPS3jZshGMG0PLTOsjikMb7++zerMHuOr9nW7UPmTAj7Mqt8BAmfzbM3nP5b1f4
WpvPvP8g8rjoRd8T+9SLqwOIU89khwqKev4t90Hr4kNzLk+VKEUhCLIYg8E9nPJ08QTrpugylA+C
aRZE6pAReXsjgxnFra8+m/io2WINL8/L4ZCpFKhgs62kF38/gec8KY3h+rb0efVj5f3Z2cnKGHvM
viwAtTAUQi3hi52w18SR9uBmiY+OQZQ+LOu+sPGoQcDvPNca/hhAWhG8o7Fvjy4jW5J6zHBOYhSY
8s+AmZ+bUX84qDxZNJq+hmxvWMmY64SBBcFovuokC34vmfc7huy31zwogfp17X6h9YljJezKaawt
LAn326a4RGFddHQBkqq6yCEoEb/n6JAjyxl0tkV3YKl2tm54cujz9wBR3Iu4iQpl4d0mpp0XGX8x
UfnJvTzK/ITC4aZEiOs3zpdLSPtuf/GsFIH+skyyYelcoyw35LAdRhqVOk9HJ7WjHaIN/s9IXDrH
5K3i38p6WOBqZ62KyZiX0KhKNGxitV/gIyAcRBR3NN9QjBK1PKfiT3jh582hn8YgFVry0NvvYdOG
gFME9brrdLKS7iGZczE6Jp2iMcmOK1zk4yXt0gh4hH+3lxyU7yg/8cIvSnWHZbxGBiQ5I3d6jdHv
6/3oouWochs16tR6ddjanTBJB5uVmcwQ/Dg9KGj7uwv3SThn03QgnyjSUng/tQHC83nClaQwZsow
L8ClcRgLe6/hS4fEP/9r5dOqAuTmti/eXrnE1l+Kklm76LopwSj92WWjDdLkFi5xeTmIAy/Cvf25
tt6zuI/UGWBRlbwfMIQxfrfmWieTORs6nvwWDwpZ6Yl8FAjdnAfqKfe4v3yv7Ql+Ejq0NmOaXnsE
3nTUcCwqLhRHUYcne1He4Myh7HGnuKdvA8GHNJ0UNiYFsCG3Trgsv2im1XlTK8Wny6K4pStK+Q57
5EOSVUNT0QDXvyJAcUCcWwhlaMPT8ANEnzE7pcf4YggvwIdHBJCNF4wSxLZsDpEW9GScGbJG7AWn
KYBZpKuZkdWxqtyUUyXEOZsB7a3X9aKJbZPvAa3dJLOfN32xPGgtRU5Eg4jnIAsICwah+dhFnfIJ
t8ReEVy5xlWCIAtAdHC2VxYZXGiW4Gymx4QDChcPw/kfoRctyct24ZbkFXDYT74/l7JOIr0Ywthx
Gn+GnCC5O1C2fosgc+7dE64sTZ7aGWzzJOD+2BmPW/sUjKJeJsyUn8c37XSbzSt2mTaPmdL4V66b
CX6HkybtmZZ4Io9/RejUjFOdznxUcTMPbIpcf1WqBgnZ8TxD9he8bagUnf+qhO+mBzxvfJ8K9D32
QWTM+TF9v62lveXbpnuTmNbEDxQFlYa7YPHO9FBCfhMkzOWmPNNdS8oR8E0ipFenmTOPP/gxmxgd
x+f7uFU4UHkvFvpzxHw5+orgkwC7vD0PX8RxU6BnneDYMtE2AnxHU6dWA7oqLbwCz1uNKX+P4GwD
cshQzL/P5AoS5b2bylGBDVhU1RGhoRJYVvRRhOweQmIL1Whvx/DI4WmJNYI8AdKyD17aBoECjNhq
EFVo7QnmvPC00BZayRGrdet2cduBxUgNq6MnF8I6UBX54eafKaNLCDLsdyhTKXV/44jh1siXSgri
mOJYHLRQIRekGKzhaBmotrmbmEjAiDOTTAQczHyB8AlwmK2km5dDFtW6nh0MbyyFUfc9Ef0Vpq4l
8An1JK64s8P4uw8mpqjuw+sOX3s+3W29AQMxMNPI9Ki33AaH5tk/5or3kzPHY2OAuINxWYClqQZg
9ROnMKyPbYF9VGTuM4EcF1+IvNl3ckYwNdOYVhbvSOYMPBxkbIoXJdhYWPH/x6XP27lDNbDfzKAn
ceZAgJ1phjLaecO+fkGs2JSqmZoHSa3MCUsB0kTHpdlO6uSrazt6/Z9X/bZ4ixlQkO5RnAAZG8bw
Yyjh8rXka6gE/3LO6R21GQH+9Po64M2xw+jEJ3jFrxXEm8d2fGQNZF84Brs2Q0jSaK1JTfD4vV4m
BlmEnR/WaeO8N8Fvs1LNLLyOGllqxpeq7JYy/YqIYJQGnucNOwP47D31rDhdzAlsX/wpqaczXv6z
i9BFbsYRIMkoZFvHuismdYFWYUOL8jsvF6bfLEWDcGLKmg+3qC/+iGYa19JXS4Yrznjo6XS7MODP
qQH2Y9wd9FfSqKZWHXOj/fBn+PVhtOA3SziILx1jCvFaIXPW8cDLgNp6XEvKepbBUXaQhIP9lFvM
KMc0S22f2cxejwJQ4q+hZu8GqAGOrqvTI/4tGNd2iMIo3jV9IyLH95cTN8vrgOX1LvOPH5YsXDMP
cs0eSUvJMdTPVkOxBpNHQrjjUcOHsWtNncFNIDr7zaI2rEp7DaePoa3wvMpq730ZLZi36qi9XETp
f0eCoG5MNhxF9UK96nRuU6WLQnq8puX3cFT7dk2pKngg+ztA8YymFDNXBfqsH9CBEMgpu/QC/e1Q
5ipWHwbBdd1y75xaOw7TkEmy42m8n3tWF6lF4Vsrqz8GtVm6KpoIybM6DszNCY9SiaZcxRsh/5Uw
hnPuD/1H9zQ4YHaOwnLVHyjzCOw91Ebg61/kzt9Wnwz8wpibMmTMh8k1cWSalMtEQVHzfKEFhyL/
D7kyvYx0pMkCMM4FBc7onwLdakLGNcaXdR6Z+9AnhHBU5JFAf8MMltaakb8y4rke28zPtQpEfNhe
9WVv5I5qLfc//MABDANNCIRJXwGTzFGiojQlVqq/j8Gt3cdoh5H8DibrDXzMvyP+CRda/jWHFIc6
FBfUeBT3NJ1iHOnNSk9CnHk8TjMkf4H8+1Xc1L9YPo0PPSUBxGmQLb2AmN8Y+SpI177ky2fi2QDT
mSFf0N2YenMkM9/Y9KmIOfE40NpvfnKPVLsVWyihB+YlIUVn5/P4qgykqpjLKpsdfQ4QylKKBK3S
RoNYtqylrIxdTadbDnqaoHcxlBJPhus3zn0sbAr45ZjH+jG/Xr29N1vMPzicI99cF0jvNCBDWS4E
+VMoZlM2Ad91TkVumlv/9RQVDlPsAAgUa5y0qSKNaFZpv5GYLlbrGSzXCUYvdvcqxRNkuDHPOyvY
1nFH9ukisXyLaeKePBUJjnT9gtKF+L2eAajL3OHp+cExIH6tuI0mXcjqJmAuApgK0j2k/YgZze3u
wGrypF6e3BEDGzuOoGHb/Md364iYPSlBLGfrrtPe8NeceFvDTX2R5ruw8nOHR28y9XrYu+1P9kGs
URryFpgB25MSvVG4Y6gLr9wGGPUnPWrFi9KhD1rGYeETVq8cINAP90KDDwJ6hppqJqrJtL5nbKat
i6t7VU+3mKto37mewGbx2ix8mX9ihuTyfpfAuWl/nJvlJEtX/Jk3i34wLIQjavK+LwOhdtQz3K30
TfF5Xwo+yClL872IxUXStyPWuj9Vs3JE0u5GaZ8ZZbhrm116a4renUxHOjy3QoFcU8R9BXVdES2z
WjsnUR8JiR9n69QDEc+v4PTh6TkiAgJmeaKx8YbGHy1L1NNld4lA4K+iHPOBsSvEZ4P8Pvfit/JL
A6gM7Wv+l2eeOnnC8jerKC0h51gNL5VD+5+aQkQed58Bk4melkWcAoYk1OVQdT2XA7AoopsmYOSu
7Zxo4FE6nAfSTpaXgvEDTjH135RQCjTjPozgoYtEB+YepFCFt15eWFMMlU7vYjFtxbRD41zKzGJC
7bPTouO3BnDMLmc2fZQmQmW99hlFv6Z1gmBxd0o58lxG5BFfgH+H5wUqhBssDxSoaoSJA4Vt1wo5
zQoMgw+KyxIhv41yB15QHzHhEt/WeGLGC/zjxe5Pt3mnpBxB+NkEkIiqs3Wyoc5amN/zPoB/aCzG
CdE3xoF35TI44rrvCgbvwKkdREeS7B5zBYCv8zuAmlhPWynTju/wuOIhPi4kaBYzf9gZlGFKAsqo
tXeiydsiWiW6tuYQyijWXv3jsB5ImYRrFvriKKcFjfe7xa1xtgU6jVOISvRI6mKFI836pvifsIqe
QsG/0kAhaR6qzfeMCkl4vTPjg+5bhLQarWDAKuun4I2xdE8a3tOxNyq/aeDgBZxvG2aaWPS+Xxgm
VbGVORdYI9a9a9Cqc9MXK9cPicBBUk/oFi1wawZBtjWHKFCv7Zzl3jRgShc/p2/hcd6detA0M8jB
JppTgxYdF0hsG9sSTeAn4uM14ZZTA15zyGb7oU79fgxLuyQXXg0H/50C3i9jyPx+PnsR++edVoE3
/EZu1UExqE15FXJrnKkPbOsiaFXK29qinErIKL5sGbb2yqPPxxsCx3RfgCball9hg7Vtv3BdEJvY
xJC0cCX4I8p1A1qoAvxX/Bt61nGWYypsr71yZFhw8ER1LvVnhQxk1Za3IHiwfs9yEXB6NihMsdE4
eVXk/onWXQZlM6ojjaG0VDtyrFRXF3lZCTTz7m9uP2liqdvaDc4JmiyZqF7j8QTou6dmzkMGGM5Z
FAng6M7bx7iTqFMn3WL7ku7AkC2FIxgRgVFrCROnQk+Xr5ndgJihYgbPZFx9FvDoR08vycVpRsQa
NyrKoclEZChylFWG4RxZsrTZ1ZXs9iJqSyq2e59scIVsA07v7sNnqKSjH7jXe/Br62CXFFkvl9Lc
yIdQ00VyLGR/3hbX7ajOlVwyhcP1grY8m2AYrv5K+msQPeAVZ3WuIeXn7bfhZxD+QUf5BajO5mvT
DMwtZgA+d//FSqTatUKVEtghj90kvw8mVlDm5+CqonDdo1UtV6LQ6WqiK5fd9fIJK5ONDo4cG2Xl
5TY+MM0fQ3dIBV43ox4TAY94I0B0KMVWFS3qtcrjmM/X7sJvsGffpbJJz3a3EhNIfvwpfU+GzNtX
V27BL/TpFuhHSVNeLE31JDGuTlb+BUW4p9lZBWuFmTLugIlmGnjD4kiqieT+oa87npnUdZwRRSmx
MJjo9uBTnXoufGhj+gmO/uaL3Q62iKJpVttJUcPmj9dz8O3But0vjn4FNZIfX9NzMfQXng8J/Q0M
Jh7A/oMCuA4TGvSLI7Wz9g3AgVz46F/ly49BJSJHFTy/BFEfhtrjqIhzB9FwDJcAG3asr5LbmVHI
ifWVfSxFSp25Z/E1hJZLTIhIg5CjmBT4NxNBn7e7Ppd5wyVQasPE4ZjylBwnxoD/QzT9Xv/HKbgT
cZn4PRp3KbgztSbIYAmrzNcLFA15mT2Qm1hoYfJSAS50/Zn+DqNsitEpzkpWMTMtHnoiP5OBs0wG
WW/WcT57zuyRsPosCJlFoAc5denO+1gQibQApiA1bjN2nMSI3dZesxfIw91e1iuX7oE2dypmpgBW
lxOiDjylAwSJuZGv8f6fofId54nmd4dEx2QCLTKkSIScr6Qf4vlnKEMNZPmWvGSwfzLODYT5eo/p
nSgKdTnpw2C1DtgaG5OIzhdDe8C5f5w8WZxYXsYL6gIL9lefG+SRupc9byr62d06v51JbRLcw81c
+ZamMZj4p7LZGiC3/VSfjjs69JRh3E0+TUUOXHu7S/AffZH9r0EqwwyGMJAP3kjNBZGxZjvKpjPB
8yYbhWGozOufGpkoKXvgO8vNrwXaCd+SXKQtuBNqgdyfaiLZIQTcP7eauCFTigppyXbHlfZFi1JA
xX9lE6T7ZFVkF7LzL30Qtu65wFK+yC5+eeHNAuwjE0WOvWdK+q8D0yn/LnS0d9OsryfG6CA3WVnv
bRx6WiR0dJvSgpJnx90sJlVQ6yLAqHQTrZdcT9Wra/QOrPjS8avZ+OBy6NCYxkRM9MATC6ZR1hN+
YvoyYeAeoZeEpqBw8JU4QtisgwieMdhLo9ZqugFCUUJZzYkPR5zjwSH354p8wGJkL5AIaxLNN9qk
QXIuG2kImKgZP/RZT0YgVsvbXZXUQWulbwEu0G0yCaMk0YiHod2c/J7Wer1RdNPZ9QvwyxFNgkFj
nm5j9YA+YXudbJ3LCbU8yaPQ1JV/2KBFgpDW8QoxDoxOlInqqyQ//hAhl1AI47eJOTxZmmSFwPf+
Qf93PoKmoVNFskWAUsBUWy8WmYlw2KUBlpLU0tYfkEsCo8cAE1NPC7nFgyA6lC6Wi2OCHLXMNW7P
CJU1i3Cg5iVK2yvRxy3yNx/laAx75o05qLoLMnA5W1TI02mxn/JiNzpvBL49nglAa31+UVuSnBhO
GXmTubnxyPUbKp//XZaV2R5zsVsuPuFk31v9dWF6mjEVxQFq6F2AiXN/Y6dm4zlbxWXSCLEcy3ln
yRnZqU0RiMRg29qlS1Gcpst3ealAQXeC7nZAyJ4sJ7AWAnXXoWqvfHd9zggud/8QcVBfuAf5X5Vb
ru8JqU/dY6oZALmfLrjoRlBp8dC1+eoIalCBmqkgPPCjO1OJ2BdDVaWH8R/6qZTQ0QnyQzfwuGln
W8vIklOJx+NmmSsrQjY9YimxeeVG1U7wiOIpOeKVFDu6WHSq/mtVMc0dDYSiPcv6ddbmRaRsKE3O
Usskzmf6tk8sI1lZRsVn9Mdego7TFpntXeqfJDDnR6KR2FltDO5GS7K/wnF0HtGhof6LtcL1ymci
AVzl52YDGsInDAUvENj3HPZ3KZUj/WzXflXkFtZXWP9yruVXNgOrPCzUOOiCRZYC/XQ4CeBmk730
2IKZI2z4zbF5OU0N9GpRx9WBeggW5HKZr2JkRGLrzf3q9xfqcF3wkJbfZwoPudY7hqM681Fy/YBm
t1HJfbNtPJ9PaWK6X0pfw5xUrZZ8osZY3+dNFEe5/376QLgK26xl3UZOTkGSib36twkzh3m0hIEq
ZLrcg3dDDrODWXgo3v3SNlQr5btsf3rlEig+8krrfCYiaDDeyMzOGH7PD03GOoyA/FyLxR4qwOiJ
ayW9XtovaPLr0j6RyLq1ntRqxkpV1pUCw+K1bLtWMCzA2Bew3yRPJzoNBAmKfQrwJF1DZypRWX/3
6RvgjFLVSWEM/15cINN8lW6L4zmvjntRpc0n80c6Z5/fmWcGaQlKibRFQWsOjLKhXcnWtLjuvfOj
GPDJx0aNkJr7ryw34tgBzNav111+XxB/lFVW/kcLsj4DLyTEGzMlSxjbFyqww+Vmtdv+asgxd5wd
CcM23RbfisySCDcB/jf8ZmXXqxT21W3EO5L0UPLcFp/j/NtVci+x7KL10sO+yWQPgYdoWRAE255r
K7KSXkwy5b7vhG8lM57MJyT7WLEdF00pHn0YUm7VHYyvzRU41eFfKfJsfOfmXpff6bRkSt15E38Z
peVxgCEKz0RQh3gDmDhT7fnZZLtcBA2hUNtHh3n6/HO0qf4FMzovrwgRnfnulszgoyDbDmGEnZik
kkcg1QN1L9VfhH6CHZMSEMh9yijSpORW0xIfZ8a7SxUnfthVndA0C2OmfbQkxZ6eIxrqJZ/ir8d5
Y2p4J6Mu1O2gNp7pLPQPs8cUpl25ZtM2KMfAoUB9E12dy20TQjF1fAfoWGvJ0aHHV3dxVnDbat/D
qLAHN/tKnZH7NIcgXh1VCtEmwOCs0//gyTecFAro65NG3B2UbMfQZfSd/w1TTReGjniqKGt5Kiwm
CoHuGiHjdUmFC0+fJZ0QGlvMOYE6VGwzj/Abm88IfWNIt1qsFat5hNMzvQkYM1ruf6/h/4pvmluX
fjmaSrOf5rVJv5SrEMY5oXCNkGpfjp0P9iuV0MOFAFi6w7BC6ZOiqnB+M2iYW+SlTBEjLKJAeBMK
uIgVsBmGB78kCTTuoAygFGsEBlUfZ3lVjrbtl/qLzNaqivWfWtrYakG8H8EX95PhBNi6kyIsHs/b
aniXj7ELpfeqqSLrJbi7O7Ng2Cpe5og6YETc1ZsGZftl2y820NBTjiU/QwSd6ic231cWFHcUAtX6
sT0o21tqCnBmpBW7VL+G8nDP0y8eWkrVFw0pc+4TB1DFM5FJQz+dADc15N3ndYa767uG+lVSUVvc
e1WEGL9yivJUMFnaoY8nxHq9LGW7yF8ZTzFPzF/8hI5/ZvxMxT9M6d8FfhNX/N7MCKrzUiuZQ1En
hkvhIMEDtiBcJnW81ZD2c3S65dvAXW88ychuESfJboVpWUfYBQ0oaFsXJMDdfvxMFStCXEcsCJCF
SvtC2P0/zob5SEl6XrftLlf19LzQRzyaVk8kfZEzBimZJ7Ofr/l12E5y4YJuu1vUqXAIUfi2OjBm
HnfoORX0B6o6ewp+MtMJu15iDKKd8orh8YNM9v0hXirykUIFncmbXQht6RoVrJLvNFtiBIMz+TXv
m5xpZl9vdDmSZ8noPt28oEKPWApKSMk8iiEQvlYyr/SeMi4SvO+5+UR4gU5mWMU7z7adJprYYYPe
SdhU8vhsQf+swoI1JlqB2IZ42REdJ9Fo7Ahq/xSTZRmFT2oPSN5Snn/sS1R8lj5Bdu6vFwm5UDvC
oMHhu65aCMvC9wTfVVfTHvIcjhMs9DP24V/+g/KJn79N3v1SNpMwb6wgfPxmXehvUL2c8L+kA3kZ
s75ANny6c4UQt1ol4jdv/0U6hJp0HEMMG8Jd6BLlikMZUooFaNMeBhiXVTpenbIhStjMZVjyG7sc
AlQa/Zs9veBGlWk69hC/oR6uN3Jx9RToG4x6ZwY7mZGpt/ZColhW0gLe0eB0/aOloO+LatqHmEaX
Pnlh67vAQqqFamhecb07qca4Pa2Sj2V0YZDoNTQHaaCycdAFfsxvygQlTtK2eagNcPfGETRJRs6W
oCdWjp/bYMtyBZMMZbtsPyu5oda7fISGzpOc4wdIT9ls5FSLj9+gYupk4ZwyY29ZndIBcfqFb8S6
ptcbDKXmQGKtzpNoN8fSg4IgMzjRiTpkH3fyHMQ/HfSYMJ7+0uslVNWitQrOkdVhAaJ7JfmIOLp0
gHs9jh1/nBDQf5VYiLuabM0Zywm4M/G5ZEtB3afHC9fLHwUGbW0jb7QSawbGNcbYWh+KVlnpISgi
GJdVpHfL1Qo/fPFbHuoxein8O9o8uwqikNezp7JJVOZHXwyc/1/xEtFFMG5Hw77hIIDXpV8Vbog4
wA6F7iMdBN2FQr+PH/+DJrMF1Zbh98xwv0pg8oSTUpDIizInt/pxYmvCgrhYyMjdqib4ErHRCu3e
NDpw1aQfRPgenAPmGkiLy/9NHXec2oCbHpha1ugDQkWyzsIYZTh/eR/u9qtz55A4O3E7Ngc6z6Px
+9+GS5eX1o7xR4iHTMVy0ndFrg87GrVqhwUw/BgZZtPkOGRMuEvQLQJNg9+tJ1TSeI2hRQJRpJQ4
4hhh2Fvb8daCM+EYfBQvsrFaYMf/P7T5zi//WpnthquXTlKujczyCkPLXaTI45Ug+549LS4Oy9v8
PuYxDuFJkhFn9bDWaoNecsoF8+0mBH44SpEhcswgVdGZJgqW9j0CK12VnOk6KAndv9Fv5F6Kc+Ry
jxUcHlUiHlmqvfpm8LgbKyrpiJgy67jus1j3c/ITpwfnCN8ZMVj9ZBMCshVs/+sh1CQgONRPmgcN
bLb3fLpGEQZVnfdfpdUEpDOvgd04YfboHAMkAOMe/WxkL3SL927WIZx1BMDcOK3tQN/tYSO5hrEc
klvmxZdyOXER/HmceUBCuERdJjs1ca0b23S+Y4hcn2VjXK/AiJ17kmhLNZtd3oTH9WLJvMdGXgwf
PN5EpoCZMZt7x/buSP4N3RjlVFytqoXXXQb/vGtP/yUjFM8Zx9MDiABJRdlUFtFX7CClgMqyifaM
P7Lfsz7rT9exYb+Mw67XWc2miTx7p3AObpUUBXYLkQIFMyYi+TYbGW/pGxWWtiznyt173e2F5ErX
ISNL5OoL1s9um3gYzn2cBwLYN6C6bMCiyI01/k4l+N0eJaMKzFj5aKxLR+NjdH7b8R0zA0mTDJ4+
yRHk1fXz7KKvUCtuTdvplANxCDOkHQpxvWhBgyoVLMHcE3BU81qKkmghxT+048ipttmFnvh+B9zI
taCwRs/CRmZ0wQpRAT5wEVLw/2bs7DNFfJAqrOQ9M4n2SvECZHDyF8GFZArMBAMCPbLz8QVLp4pv
Wb8LSqdfIhpo6n3Dz42R42jI1qy3+m6/lV9SloEwx//n4v7fPA+261E5SobAs/NFeFNs6D50aqni
QiWgJtV7Jgr95bQAQpo6Zh7Dgqi1AYeg7RungfS62P5X5fiychHbJbTNuaKQRLeppSmEkdH6y8hW
80SUqRz5FtOuQO1jSQTCmbQxjATZDZcMdZYtOF7B7+BTJ5JdzjtBU+xTVKADSRTzknN5hoQancLB
WIcsw7bj0YmCz8Zpv8WHnjM4nuR7r16jbWzcrpvMCb90L/9KuKhVcTO49dV1L3wZ7U9eM27t9ngg
z9lFWAz+J79mvcvBE82iYfE9dQ+hgsdHt2isnCNGC4fHzgAoUbcFyI9ubg8bWgSxgrlNqNUR0hHZ
4P12SnX08WpeRSrcuVuBonBZh/6nc8XT3B1qO5YcQbEOwehG7EAj7YhcKPoNgALtXbJnCqdiUsQt
46xWZa+Q04QS4uUGGJiUSfgrhNs2EWksols6BvCExvoY3RIdcqLkfUvxTDFRNNafR8UzW82YFqi6
HUIq8uwpZxNnpGs0s88zLGCblR5+ezuTmRxL94JKTorxkvyaG0dTfHOxZNEbFavtDgYXSzkPzold
BfnXUfNEFo+wqSzLe6qJaGz3WxlJkF4PiE70p8xPtt50vh+kY42DnrRFwPRPAxzI6i9U/fzROgT+
cI/dUj/QU38iPdwRYNW4M0sFpdGfwSndXrHhXj9au+JYL+gd/JQCryc9G8aRSyuvkor/FM/zcf/D
0xMRlL1jqE0BQbxGZKj3gLzOLUMLQk83FrlyPUww27NZYFHqagcGWgG7yvFCCcld9fcFUQ3/wn7p
D9zEhx+RqU9MZRiEWkLgMBenwYR4cZFgeKhAT/8NG4v3/vqb9qqHHaalMtjce7/OUp2shOrC1e4S
BC1aKVkSPOLgH4qUON+2eqt5neYwfnDT0dQSWBMt2WCBOWuJNC49P/SwACg8rSn1yUuY5NVFKnPc
oTdMKgELMyjoM/zviD2DRdXGWNn/R4P0UEK2P3aZA1Wj5M0vV+Ktpwseln04ZqwnwhZWc8PzdpR0
CnM89O9GYcbfjbJTgka1WSs+ZTPFkjuGsRFVaxBG0DZjqWwRRY8qBL/uAInxFheGQCE17Mp13lrf
uLKdFBRGHqQL7ODJljVKIIfZIzLe2GYDJubx4l7zDm5LQLjyqqsGRySITO0hcE6uh4Namnml3+E1
Zg9xH+/PiBhR7vkaKbGLjehJZy1Hjcb/WLfJ2Wcpml2Ihxz/7xRzPii/8Z/f9YaT+ORS20YnBjf7
DeB9gFcCx25m/x8nxmQuuf4mpYRu5rcsQ/Q24PXPsOWtV76e4HpREXnJvYEgk5VxHyPuZY5p+oUB
A7yVmdk85gult/IGIJSjhWOtNWId7xIgexBsj3XhGof6yJ4VWKzv1PbGJv3HYoC0q++jSKNTabVg
R1Fo07E4nL4Dabj0gPvnpqTcWmeG4GvZYd0v/fep24NCvOqZbLTURA8e8kY5dhrDq/vqnnTEtWAZ
boqRHB4ERjhQMc14P3tsnPM+DN4n1sNIJoy8+6oXA5WG9Vq1ExThi2FP2z6jTQo7ZZRE5Jcal/u0
aSE+8DZIAt/O8JgRbJBAEewTMIjiR8SU12ky9QwSuITQBex+8Vjs8YSUDj39GUtxTMCoONqJ+4CH
fUr4OsALOWjDHapFU/hrUHiLE31CkST9qbIeJAqf1Hr4YlPm8zIfPF+OMSlZpCiAbNSiiPcRAM3q
Ft5R0rs3W0gu9OsQr34UJwcAWx4zRntWkCdCjFlg5ON8ZKP2yDrPv6cScVrH8KVCTEm7msGUNXIw
kp7KAYRMFYgelfSjD4c6DTaZWWmKOk9B6KxQH2Qa9GP+D77SnZNLO9T/mE6vL3krFgbFjEI2pRHM
4FkD8QdAcJtz767zndOJY7Cm+0IsAfb68U9TnJqxodue339Dviwn1uEudMgJbXt+CxIa+3rdFMeZ
6runuWYWcHTm428MSlVrPfCZRiGJHmxIdPsdeDevkHVNhscSAO8dD0sI6PpxXjAllMUHAXjvkqhK
VyVjMhYZ5b2YwXmBomAccmSn7WWRDOaoaTxM8DyPCd+thRFp0ApIovPLbsGLP9aUyKhYjR/xkdbD
ZhrqSXbNhcGYlMuzZBaRVec7RU04W8HruWpFqDkyIaWHONJnSUVlKYXhYpMEL6kaJYy7S+4a2wRv
7NdBOzFxxNYZIX1m9d9SX5uY5dZ/QMUmnO7TucTc7/vjntmIcHGDwUKMF1eYSZY4fzl526QC36zw
+/dgdLS2/FgEGI8r3zlLypzjdniyqOoExKFXby88NAyt2dy8aY7kEuzidIX/4IMNucrgnXyzYran
rakuWjyDERc+zKyw410NVsdB6C6CX2v26ZCvopF04245EBS3/9VPZlQ916iUWwjMagg3w0cmF6dd
vdbjTM5rLAXzhvFerpAtmbrP1bnIzn2Y3FfNivYKITuHZIRQeSkffggyA4Nb5MTPPzRYeBPU9BCc
fOy6wQc6UEcTpKqvdMh2hQTFCzOtaRPT38FTH1jRZWGpvTagT2ARgR+Vl0+k/9+UteniyomKNksD
jad85Pb03sHKUUWkqXoKXXYqQVUpZ65b4lquUl9ZFHCgWc8eJ9F1mXwyZ0gTVZgovb6/e0nM/jkD
dyPHf3oEEUtzcQcfa3q5a9iMKBOzsLXjSKp+4lOzwLfCUtfZVQOoOpGVbZX3k6dUytSm4IrQXH6l
KNtH9HU0ZOq0oEkb1lg3vbdzwQVh1JA7pe9DOB7aSJW1DehAnUfD/K3Ec4ICBllYKXAH2etYBdVq
erH3cp7X03S+xyxdHHPzae7/h1ZR2G4VQodIntnubBQXCe3FTKh+/TcNDiNY8QhvTEwQWEz4TTaH
BzwRXri4NGowqutjvemZ5s3q/TAyO5hx5f3R0WcHK/s7t92ttoxLF8dmdG0gx3XgmbPmIY7hXGRr
ML5fjq270yNCQPVuVQONACZYUSMfIvS3dBytH8qdEbzXxTKQMVDRAZQV8jhnvnmAGjomRPojbFaj
vvYhwQ5vhM7GE20KWmITRDYsC/FxWfsqEgit+lO7wFXPT14djILF6lFN08uYYeDm8buh7Dem3Lbg
rtT4ZISpkGdEfJ3bY3IgWu2stHUvCeu5DNYbrNCxcUJL1s+lbTLjZ4UPi+UDwdY53Lfnnuh/NFkG
znO1Zf8OUqqg3P/jnMNAh+0SQQXARHogDSrozNtNPVEYeH5e6TMSytzBIHt0tv4Bd6LTYpA+5x+E
7IaO6ChyA0URIxDo9RBcMeuwWwOu/TSLrhX4tOLyRsloV/lAMKV/576sC+drXvRfHZSWIKh+D4ac
CmGUTCxyJOodSTep2e9VA1+4Bl2nVt9+nWsmZZnWbpSZwmUwk1UGRlxw2NHVgBPY5wvBlirIXjJ8
Xv/V8FoEs5WXCwfC+7OKlK2YCasmmpfpJUTA8PBNtrq4kWO68J9ryNU0/X3ahbApj5lhFlE7+IUN
b7/IiHeaVdm/1Bf/QcpjFiovWtjp1GXPRxWFVUvMMN9GXmy00Uq/8H2WLH//PItSCH8zzXRB8cdN
FJDvGjQFkHDNKLzIYCFlUeqhKgUZNqoSGXt6i+EMVs0QfZMC7doHt0U3I5nfFrogpigHF99N0WEI
bfXfQ6tua9hqQKadjBTITxGwqJwdEoKyp3NbQWZy3gF0Z+U5rVHbUTrjvP7aTTaUIt2YJbOLVXc2
oWNQNfEkRQviWe9NvOO+gxyNPwTamY4odKBvvCGi+EVcNudZmAMVLI9VPjjvTM8Pi9FHkQdgxfLc
2u1ejhClz5gkWDLt4mx1Y9kiBdgZsT3NVNXHKum7RtJ+6fHi70Y9gJ04P1En7otLkdPNUpPqaP8l
DRjwz/Kfhm2r0o5zw51agjKCPoy4V5URTmAzcBQ5Ya/raOk51saEJDDnjd/3JscBZLbymrBM3aU9
zBuUDDTB+3IrqzfgLeQ6e9KQyn0HgDWcxFUTfGFVr1YSW4Medq//arhrJKGJsrV7y8y3OJ3qVJC+
KaDftFUujWe6ZhbsBhpv79dt7LQFZrUbSr6hl9LLWkpGLJ1unakkxRGd0aAVEzRZm0Hq5BTNDeZj
vde9ksI3VrEeTsSPxSjegku31BiKDj9FcmZDKQhiHHtCZudsmjHiWupDhvZmo5VGi+pVatPX47y2
Aa/cMBsX4z4IQTLlXZ7fxQMrqQmVSweccYkPm9BRPh5xJoVIHR7IJcL1rZn38cHbLF9q2VnlKMes
fzNpvBZgn12rrKkX92Lr4CjVVPp1cABs8bWzS2aXZDcGdN2uqJ7xspiWkZ94VOUv+eUSP09kxM6k
TtJA+DSJusrHY3uvLPHfrsfSf8qbm9WQkIBBsKjMvcN7ld9m+jUUuoCuuw0fb2/Hk8nnqr9p1Cjm
3fbeZjzXTQAV0OvnR/sAGVZvG4yKdrxXs41kC+wQAUcL4UNnJ6JeeLj02v4OfUuD7/DO4zb8evHf
JLxCu8FgUE2d03KJcIPm6OjUi6XznWzkKq2UIjXb8SorvX9MfwUc6IrX8W13UK5zhh64dJOyf/0G
HDj2r3g9eXquhXoOiFYZtSBDqLQPz7sK651ezf5neReZH9gckfDiaGg8w8ka1bcdJLmZt3chqzdX
eo7uRNE4NFt4/eq6KChvXcGdi32loKYIj0gC1jHVKv09NvUP2Ac8KGIVa9lNACjxSh0gmH1RzbeW
ZphJ7sfoNBom9XwMrqZ1Mopfe4e/CzzJelrfyzMew13pAMlS0NrBhVHserZXYj9dpbB7+M5qerM/
9RW6Bi41vv9bfrcY9btY3GZ77xk+AXdHxIzfxRXF677HbCUqNmflOAAV/7JW1WF7FSMuPNzgjRdX
yDMvvYEXxSZnATAcQWDblnK1laf/NVc/fSFk4J1UYQ9Vooz6hsPM0LmltkQADz8O7A8MiFfyGCo3
gv89cUfc0DV++GK6sDcbxinbKWaYuZMq05/lSo5zngBwndyro5JGuDYYCX6FZ/VDQ12KIcmHVlos
XkDQnyvxuRHL5YFM7Rs+OsGxmNcK5ntHo7rkuAtSbhkztQ793vl6IDNhywiumUjOZO32Hzu/3SbV
TWgKETNdpFreo/adPrVI2D+FJCjFihbCaeMPZn0ZZLTRtUg2F89VOoIQvOb2opSP6LqcZg1Pz2mj
8p8vaLvQjngkSztUOykolyINHCT7P9IGBakKm03kFgRkfg3hq1LInbaAtd1/JZ2huf1yGhWvVeB1
vnVWihJSMq+PISJ0OfNAJGNv65WHrMlVS/hgrOSby+4GPr+o/pZjlG7XTdSNJbOZVWSkgv0CqXOl
/gDzcS8xmj8PpiwOhG8/XMwt9KIXQ5B2/Uj1bHoNtDkJQ9UMOvOVVZivN5Yq0hp5cbgGtbRzWl8/
n9fiPOctykzaMLzcTbyOkS7vyW8tYsOy2L9frBJegWPPDzEOqWg3vXSqjmL9zVTMbaNEBS7XR7IP
i4nym3h4Vi5EwvGI0RKCpMsrTertQ94J28denD1J4/xkbJcVSeaY61lfikdnHGO1I5FhZ2Ic24Z7
OqeqQaHSyQGamSEB1hVA3ICQ55F1W+y0Rr8+lXv0hlBrfrCjvVsPDNcKI86MgkvdmtK23xc+hTwy
P01LRpkcmE3CGdcNTNLEUWPXDaQzpnwjkQ8Gox/DhQSc1+g2fLnTK3VTOPs9zwnqXcP87kOj3EIZ
VJEDRV3m620Q55KDAVYLlp4gBSt/RQv9d34N0mU+wh760EIh3FzI00k5o9FQOTsYFm/jtTYMVBLy
9m9399crAyzLuIlB9hiiF3h1PdL2DKUm/B5jUsWDsybP9/maulPVRvVAfdOsp+GikjWsYt8aWuQS
C7SjhZp3DHvHEvu/JmT3erHFnjzkWlqdk8mp+bd7Yo/HO+mAoe9VVqzEgsclGurRB6dtvOtSMWW5
/aM3GBYRBCFwXUzAk9OU6ubyNpW/Oyp0jdH6QlNnr+rI5RCOXZZ2RcJXQcnJIovaqc57mpc9ZgJP
ycbb4zats2clrL45gDRNEomFNaBQ13K7jRgwr7NPW6Xyp1VcEliGONghxGczc9jjup8Xz94hfohe
mzsUiEFoUCV1vAT/hWKCorRsbgKWWEL5fpJacWK7zSzeny7Q+ML1VjHwuVn/2/AyoJbmB88DGisx
2nziJ98J3xp3HTV/CnEiA38m0lKVn3830eRz8Nng1x8I1/+Plwc9BzraBzEJLMkkA1UmO/18ftVC
ASmNx8+jXAK51nsWmmnsLQUyi7lc3Y/j/+Pi5Ch9nqcTOwfIXxzSKXBeINa0A70jdpYBFq9WzKri
nIE8CggF3sAK2giAOvIFLa/immG11ITVQtaPi/pUCZx/7qx6aqA3ieRaFBNVMMs1QrWN2pzEbb9E
LjOdHEjuKLOTxLNihN4q+9qwq5ilaOo+8plrLEHd59vtnSPNM4lXuU+vDbnSN4XP3fHKcNtAd9g4
wN1GVOkrndYE3f0Ym8qlVcbOLM78qbfTb8nHzv2ifUhgvRUAmE4qgmseb7aAV5MSPxrCuobX9KA9
O5Iay8YCPA9MVxPit1vgoSNYlkfF4Sdk8Xp2seQA8Hsbeb6GKav8eNsuvUYImCHZJbq8GEHTOBED
meu78TIixFNdb1SbcxMV/m4OonWhH3BBWl+TLSVn5p050W1vBkDd6ahXN94xHTfa3UQBkeRkMQ0A
/T40B891seuWXT6JNCn5oUqgqJut7QfN67mERj52eIjGY8jhZJ+QJB6KVDv9RRoN6swu2FgBFRWR
G0GWdX5B2kMuvQ+0fwd9/eeM/99l+CnjkVeye/K3JddKs4Ligrxmu3zmrBQcUIshV12jKelNebhy
AdhuaSGhuF6oDB4vybUqV8JGZN118uVRm6AsR31cUc7gKCXLp1otJC/Yon102FLdVrJWwYIDVb4L
3EFnYo3RoJRGFpt7bDD//CaPc8RoIMwwiLLN8RbMQl28rpuzdUlVjb4i2cKjRYRmJEfUy/w5brTP
9GMlC9te6m4iKAREi7BgigJfnXkJa25lw3UJT3HCE8A7UVx+bCXKp3M81anaEaGS7HbSb2sOpXNu
j0/TTjUrmh7xRZXQEvojvTi5XO07hcNf+d6XtCAPDcwUR9fd86uMRciOLFRKJNbW/qmZDeGxSdXq
/bgjINdthPbDWL1ld9FWkr/eMbyCTEUvqw2y/b2ECEntdrjCVtUtgzVglg3CCFwmi8V4M3KoC+Yj
kTgYgRtOJBBM/GOnbC236O2Pp5Lju/qA9FFRg0UwsELUaTvzjdRscDbixAs/ItmDw7Xd2pI+ZkGe
5FkxjWZjBgdIGOXkEpb0Y9GaZhe4x4K84Qvu+xLy2ORE1bM0RgtswdQVW+5mDFaNPamVnsFGM2+Q
pFtmrDw7TS4MbC4HDVtbQGtdZkEL+q/FcwhgDnonksk88SqVubt5oCNSUyKupmA26aJDOye08vEB
tmGjFl0/UkqqW9wO7MeiomdagcWdYx0baGdsZTklisSoSPAy/GvD+2pzjzS8xTBagaXZ6EGig6xQ
VgGp9Wq/pMoDOroqIBuqYc8xzJXfSPSzvWXDVttW/05NJnGpMm2/PpPyAhAL6rXMOn1Gogt13Etp
0g12NamxdKBBzz4XtR9Z2juYVVd8GJdp1if//EhhNdtdqdadODS40GMpaXWdCCCoZKGE+54p8Y6K
1uPQGtOgs6iVWnXnBYv2lOYH/GRZ3JwpfsYwRXtDoQTg+ot5S0t4EBMtaDNFVfS5HMJYnQBfiov0
0azMnOviqCh0qWmP2g12W41x4Svc/vuy2NHMUe8sP23zH5HL+8Cr2r0f6LCRu+3BRxzE3bMFFfUS
EMCXWhmkeey/5GRYmkTxVQviLS45odhtoSSbtlIuh7TACMO2BUyJ9UK23JnI7pMQ2TR0Y5qcEFkk
WzJRiBv2NJ0JOvYfUYuYUCydj4Mjc3AuonbGVqFBNZyqR9qXOkg93CeLlFJC1LPLHv4U2kZRokh0
V5WLWAvUECMg/rAIoetLUlmaVfKeZRN44ZfQwQdR368/rXRi9/sxL8sqA+Re1TRfqoFWgT8seeOg
uN6pvt0rM2l4hK4w//XfKrNQhtQYnL3+nnJF0zFjKDns+eXgxcgG574Efge2/O/hBwvgepKcPj7T
taBSxYW8gM6etbDMF1VZ+QDlfEz0/RmqWAa+B5w0QA15SfTejDbCfFsT+igZeuUWui2EYUBtFR5x
SYb8dIPe6MCJTcHiBamen35t6EHQcMBGmo7Jj1pPa3+p0yw/LYR3qtZz+NqG4hYAdrvkOyA9FEtj
8hlqeVGyRXbeEaorh0L+fsG9a++FOg+F7xRXuUHEDM7bIMSvmAptCFxCqqc8eQvgMxdH9PTW99rJ
jRn5I07w5v5V5GQ8e6bFuU7T3hJJVNs/xm+CnagTCGAf9weqAHPIRZEJ44j7p+79xkrEFh5vUuzw
B/J0n9f8j4MF8pHpswWQt/QERy42x8jyA3JmVkW+c8YBoILOTyDVOdDOjYVouAxwS9crhr+XZ0tL
iJfXt2jo0fF0jmOyWMpSSxh4wh8HgFZKPfgyjzEzZEhOY9GRZLtuB6a3bzIiBB1iR4qkgpqW7dAk
2+HJE2dEHl9xfINgRGnrHZUYOxRzzlQyv6aenp5eIkd51oeWQu9WOIz93SwgfdKgl/GPqvQVltXy
wj49mKpSMbFNT87ZjL62/6L6nO3WKeVIItWiVuCnC+DXanfUFeQHpOAKT0J8q6A4XFKTULyBLwWL
in01YMUyTztlzJKCkwdECpvlxP6n56fXcNk8eDsi66pS9QcuWcYbRVVzoIC/aGzjRHAJkhnYw+YM
7SWrDMzKz0UU3iPkTyyYYE6DikLQ7Ir29APhf4M1DSvIdm3zvzpJryd5lGIUOi4600ETknix+rbL
klAdnMWkVoQauCObbQuDb/uvpS8Va+pCyUlTSAhjC9OoQZAtsamnbJRx8eWJI0MUWeZT4SZUBugZ
tN/7+3AgoLWc3ZJ5RFcpBYr71TjLNd2tcUjOYsiUv8iGug9+l3g42i5b+TCsX1Uxc5syVL/4e1S8
I1kbHsw9DiYenEchUUvmnRO5UiK+NOJxOOofgcb5xxJ70oiYUWstfKu5AMXC5c6Xe2l2bk8LMerb
WEzfQsMmY5MfE3EPMMsBsBXasC9NqT8FpkxldgKOg6897xjY/vBoXtXnEy5RGbjFTmtCIVKUpQLe
QH25D1eutRZ+rzFbkg40Zq7629S3djcHp+RdmnegH+XKqOozuaEsKQqsIfkWli1w8DYG1+4MevlZ
mkxNFdpCW4vJGb5wNbpvSzbH4kvCV9Z5fonlvB9AiD7KT/94xMSHz06o7tM3YkVdFyP87Qu4kZbI
zGezQNOj7CZ/tQrXLhRexAK6UutttK0P8lRF1H7eGWLgDvgUWKKFWRTnvwyTeQhZqpDMKbSPjKHV
pNYQYN6otTo1klM1youmEOpP+vwiGXVzXLnSuJM5uHH1JUJrIa7Ub7LMK9b6C1MFTJ2Ya96WT64r
tURtB7H2URInTxsRt+ZIbKbkfFnjCys9JisGaUDRWixx34ANd1miA0KCxwBhqrcxE/c/R2fVcnos
FYle+knJoWx+BzJqo734in30IIbjI5A7mGWXRj2n36Dy2W7X14FqxQTZYNvEo7osOepchfkW3q5/
eRaKNDgWFlBWwc3XbGPCywfhBnlW8hzdFAESpFfWm/8RdmVoDhflN0KIykFxWrzgZtITcfjtcYgV
71Ug5jY20fIctuGkvDQFMFuXSEt7DcLRBbKXGJOI62NEEUPC7RbIH2G6baJRyOpVwy8O4r1Gcrcm
oQt3kw5VkIdOjMhJ/eNG+b+JSyKLEHGVGk/63vhBaWc2afpS+MqAbD/U6gJGsMPkJOrfXGlwifLZ
j/tv52FghjYideMuvLquv7RvKkayvhQEiTNPtMaMcIgCtBBDAR21fmcJs0+BUABQEADAdt93UnRf
5p4IXEPNgk+kzj56QlJ0lk5c7fNnpeUv5Uwr+1SI5fEaaS148rqkQlCqSWABSL+2ZecvLhdgCsuq
qk/9mhEEZ8ShR5gzwFnd8hKx9TpwXw+5qKj+QKdKcrfK41p0Rrwmrk+FLyqdkFB9afVVVKo4F2Aq
UUrdilMgpNw4ry1e3LbYQg7lPyTQRuFk+Sw6yVZxdttRj/D2sYuO32tXDkqnTYfBSlVCrzFFMiOj
XJdHqisxW1Md+SS91tdh86gu5/xrql3YQ2aEu0/qY8PcO1sPuODmJaWizNA5phWUIippkP/B6j3O
n42ABRCmIw0WD0GRqGDoR9zMIHBy7t0/whYT4+jAYfsBqOHXEQ8rGJIIk4b9NBb1OLxKUQ6LPF1q
fvpO1ggkIghGXXcA+6Tj5DVCg5FsEMDC60pmNuqmn1nIPLlZlaWo5g0TJI0xgstCmpQ9kG/8TOS7
R7SChxGJ+riENj/Fx5RHEMV426XCootRLXKpJWQVtF4iU/+HZLpqc4EiSjAlkuzUiPPwGzb+Agjw
FMICM+Rr3cQfE8whobMuM5a+ajA7atrSP4J83ryl2pT5Xoqtlx5wWEyc5CtmB2fAoNvzGyXMIlBL
GtjLpjP44lH3c11Htl7fXmjlFB98prLEzREckq749ccSGdXFfBI+47pRTaq9wJWKkr3Lxodfcfmq
HOZpNElGoNQYj9gxYSyVznD3jQnhT7e59BwFrOV/aEMst9dGvtYkyiGeU48FHg3vHBvqJqIbEL80
5CfaeaTXbrX+wQpSAcG952dLaZdLYIHqQZwESW8pKBAcAYF96kcWkNu7JiENU1zd58sNSMdfx+f+
A1S/FSa54QQLmI8STFTpSrSl7KvgENcDrjHWQC/vqCRxEJD0F6UVONDAqwzHqQQstqyBEDci8lqC
rfXPH8ydychUvW0L5lifyQJXx8cGaSVInGU1PZEqpGrFIO5eKd475RVZxCm+IXbblWe2m7meK4Q3
QnLEXRebdYUSfNQsNUjSr7X9Eo/HGMp1Bp5ZDAUPJ5OF3Asrusx5SR0BDZsNZ3a+B5xxkpAk6OPE
vSICXkqDvMnq3LzUl3JXkurqMRZwN2YcmlXy1uGT+x2VRcdmYF602Bb5eVo0mdUNo6Vzoc182BE6
2LsdwUkytKTQo13Z1qBALQCzu7CsRHJIgpRdihue4NDgSHo59pP19liuF9Ns3xVxMrPM+ErhSNwX
YofiDOjDH9SJ/HMFDfFyRDDoPxG2aL+ZObFpBFvE9gbNMAwEXeq3j9ln1OxmC7xWj0onZpbwtlSN
0y5lCYBDTxdD7uAIm3ZvDCyJPD43vEs+FMU3815xI4SaJbmXcXd4tWcaghW2D6Pyvo2WiqZTUzq9
3455yDykBUXd2Ja72fbWxZq+04Qv0bquSyNqnspDKWy6jzIIcSGB90gITMo2Q5sy95z+q0pSxXSX
yEAK8qatUieZuTbFCgnHzwfKkQiK+ccBZAwqDJs/EHuQbVwdccSPMxLrJiaEu645QtCIRiRQnrW+
9LQTheN18QYDhRwcOCaDiJu7LQQ+a2e4YOob+yRkOpJobN7X6ioUd1LguNp+zarnHdknJuYt/9mF
pkiQMMM3qRTXRSQInioIbSVK8qDDddPC2tK4VetpIU3Oe5kdBVhjMehIADKAkBrrpJdjIapjqObI
WgOqRqUGxI3u5XiyyfMwkOTDHMnSqYK13FwRR17dDgQOao76Ln1zKqBiMvMm7WydS3E5T/VOrfQx
IAJlgPohvkmvfD2I2zG+E6d2gyDJRzQYIRQZIjPHhygt/s2G3J/22AcP3MKkizEeqxnbCjkR9cOZ
7OFZbOrC9Sr/oV3kmdOSvhKDpUUo97ASduwCVQR3KNCHRotwTDZPY4sdAE4DY6lC2P98JFvsgjtQ
MHdgDVfMql9NjEQjojDnYt53gmwsyrRFLn/g/g3l2SKHqoD1wCZ0Ww6p/PnVJonA5rTO3TUSCE5a
ISAZh+E81eh4xZlyrxtUSXjNp8A4VcpyL31fqlwv9LFgBaloHwlyPQvQItLU0jBhQsZOEqAuJJxV
raFfM6kiLBqXQBwrWb5RcXHiwRchJL9L5X0CqWGXU/QAgDcX4bp/u1efx3oKIJCzPthO9V+ryR+6
Xesob64KFjdoLcbMeDa2ePazcU8ARobfwr+i1xNkYMpDtWMYuKSAIlAru5pEhDYUJNgzAbCzdOei
lTi3gOzU9fgLgQfoXcknzDYqj4qhlxsX1yWT7vQdvunkvp+ZzKCNJvoMgZJ3ZYZkHoFdR8adoEq6
rp0PxQyB9yfzLJHnz4MKze/AM7YF4tr2BREvCKbrcGSYajTjTSpL/VDINIsFFmcNUoNLmVfCYyE2
BVf08BRhKu2u+LS3KzvIQUMmB6n8Xk4PSaJFxCUXTRMzJESZ9Qjq1dTv5OqzvEcv1gDKth9ncHXB
7YF7DOY/tjGDYyKQBBHcYd3pY1E8gu5Liv3Ujq7N8qVNyS/cdma7EuApP3Wfz6nCpg9EnDkVQW6i
HMCKynKJe0J1AfZLSsl3EYDW9MXCIswHQ7r5VnepJqtSdP2ZGyWROjeEyXyGBru774aDkbThKQG2
8WmCqvP0NzTzSS4vMFTj9naF0gnc4oizgX+C79m/+oZRJ/VNORztGqBwTRKJPlFGcFCJ90fFvxCj
NLq+a91Msr85FoywyRHL0+NDh/CjPhpWpOsB5S8wa0orjsvRsx5j9xq9oLzpek/vFd5JLBvhRGkS
3NykUfnGfX9kUvwNCoZsMjtnBeI093+sNEBze23M3XDyAY0Iy1pZ6PkwARPhkX4dda3ya5Op+0Li
arK/vm5QDFNkiz3dwjudLVCZ2BQrGyhvmU+290RyyH2Z7V68fbkMOJbZkmsv2lBVeApMBKO3Wofe
OfRO4It06GqB6ENPDzWEOtf29iv+qQ2B5riHOr/0GGUgi+VJryyA/eC1SNTRvJq7dbuFpU1BAf6T
0Uph1CSeJR+Wo4t/XsNi71SBUplZ7ezF+DR++rJPIsnxD4sKQ62Y7S61l/ZqRszjbe+OiMVuXcGo
kQAku1AOUfu+5WJYkog3Zcldvw6fNsKyYSv99h1+fFEVWPC7GtJZgl/Q7VOPEY8mkc03Ovf9mO86
+Px29YEXXE+wBUMf3LwTVuENP5ByP4Vm9gwGtkp/VDE8svwQjn+LX8Mh34WT3/T+4K7HxrBL1gHk
xm/Fdyoa0F1+aIIxJJnENMQG+/Ggd+QeTlQvMfd4i+LZYmPb77KAqD7o3w34TMaECn2zWYCzvEEc
8t9DIHOPSQhGXTc6M5LJ+tP8PbeaPZFsKHZDOMMcH627xZYtLFx7R8K/jfyRlPFhoms1p8H4ww7s
D7KctYkcu76xQ6Rax0ZS4IcWA3bk4MMGP2pMfrrqGshLg5j2A6bvhkvAHeKkdVh5gCeBuxFqSh/N
iTHTRFnecAe6g8QESkWPCahvQKYUuZfGqflqE/Pcih1p7F8x0CvWLE6oXvW67o5ZyaMaL5G9KWMt
DV1Lk33Dm3PSw23bx14KHr1ol3NhvgGdpbqgucYONLMeO41D0ty9uFodkg9KU3mGffTbWxEzE0oU
fOQoj7neu3XIs5KMFtWFjkM+g6GNwasYAPnQ4e9Hn57S/z2RCBq/rslPbiHsgIgHQhAdEjEx+V2L
g6WMtBhkhQDyDadfMrx6W+3AgvKqgBAKacfY0u6s96dMxf9IGvqpXkcMK21aaIYkiVi3TRBu20le
mt4HH+DLoHvEelszIqXTnESykprxB9V7+hELPhy53C7BO7maU+y9uTlWfhGwZu36TrN6YHnuz8Lt
7KlqJ8E2zgTu3uPlnEKnu/LV4Vu2ZkQU9HYbW13AVpUjRDbnTAy2sKR+tG4SGS/RZVztYvYM4a6C
xJnOU05PH1EWKV+Z0ht9hYeLQKw92uEKvpnIV9bKe/LSkas9q+ADv/yc3oGf/T48500pEPpEpVry
EsSpwHVzhkTpWQsvJsMgKPBqs0+7dtv3bQL0U/HcYGdUPjHTEuNYfrZ2ahCac0pNvBepj0VcLptb
tB0uJIFh3SrxWyUsFUwrhhaRBmS3cxPs4I2aXuV5sZr/jJ+vofG7NRyJTX/B/PS/ciexgFZ1FB27
dxQACHVrxKq0YOXJ1ezqOYxP3oE9Pt5Lumtsc+KuDefqo7Zf+rDrZ0TFvOW3rio5oRYeTwl1ss1i
zysXQlz+5WN+Go3Ek8nyKkRiAAx38RaIFP4nYXe0L2RhYE6uiMXfihyAlphk1iRqSp6jmuSU7wwl
PMtkeAMv+YgzZiK7GRUdJk75g3sMmyGzo95bMEKqIXGSlnPrS2pF+xSZVDiBWNJTU4Y2GiFOogDy
ZU6pKc3JotW+b1plxBYFBL6joxztqSOjvdGvosDdAcFyFZf341y5NH7sBHEuMIhhMvTXr5epXTSf
w1qrkGgVADHVQidHitVcRlxVwUE222RsoFyoH6bkR9I05leJ534HyviJj4mZGE7FJy5K1pSJlyCL
0DONTB7Yq2IP+zmLHqa31Aie7+Wd6JeyLiXHy8fX660tY0sWfD0Nm79Ea1LKIhfn3DLj+UFXTJkC
EpvzjrnemOPm/k5aAGgPrqV4ecwUG8Lp4GIuX+izRbDgywKvol6XMxGn7gkF9W8Gd6mBa52/2LHv
JjsT5fwnN7cE+u8ESQhX3ELgLCyATMq3AkMzSGqGxaXhs+jA76SXVUv8ejhFNOFEgKCH2WXzgH9D
Dt921H8e6jeN7DT0+gIRfGiv1u9C7hJOynOApRxuYXbvNZoWACWOxaDBrhQ09CccdajxGTcyrd5+
EoJQfvKOXIhGHKvv5VoYlWnSD6GO2lgMMQUjBzKjFJT6eO8Qsbpep7kZqk7o/5fQaQ5ywdRkPMxx
QSRZ053BwYbbiWYQlbbDD+hJYeaBwco6dBd9KN28Hhe2EIJEl+kYrsqYbPq2zoe4iNiPe7Vz1bOS
ksUc9E4xdN0REv+5+AvQxbIVrcUWsRPlTU7srKRmYSyh+bdVrJ7/6ObNUNBsxSNjLzgH1V/WukCW
bPoRU5cf0K6M6f327QXGwFk22/MIe07gXnxRoh/X5cHDVNm5K1aFVgC45uDcXhpIHvrl3u0ui8A2
5JZIK+sYeA8rEkoqcOtov03Ivp9M/sfafpVc/Ed9w881hAGt7tOwKDCNnBq7pRsv9vCZ88Vjvl5J
93BGUtZ1mtyp4G8HqSPXZy9b4Xpxuga2F4DROVHb0fKeoMT/TrmdU/LzZHDVGlg9IAOU4J743JQO
hPBMjSVEUgIUrBekRv/RxCh3c0vsbcCfEIT0XxBuRh+PHzVL3ZEQPEW4xuiOgKj7rRQTpnoRNGH4
l0jR+E+VqeAy89jGJ2Rw3M1MgiPHixiQkDztayE6sE2/Oq+ey/FLZwD4roTJlZZy0BHwAnkA5NO9
pSocaAcz71n31PBLtMgVNaQH7ws6J7tyaw2tNxsjnrmH/eu+6Ptep0SZ9DY1/hnUFl8NsJ8N7q4+
AanzfSl0EjpmhZb6iDPnyZ6gTdFvlcuvhEqRMxi9Z+mq10wwxL5GKl0dtanxmzD4DIfOIQ2bhgQt
UzIve0HCEzHfXU5CinYM1xTXdysmwehmwAv8nPtMbLAAuOSXDjdmRK3e2YlgungIH+wspgpwvUyF
h2q6wnaPz5aB7KXYshM78AWPaLHwt7CSYQuqOm+6Q008ieA1ulwhU/gfYFOfXY8XtVPBpKbVv15S
7chonh3EE/OsjJ0kYpa4w1dXPgW0XSMD2vyIaALj26LQXzUK7Lron386SOvprArjjG6OTqS1oMh5
bkhU3xinCcMJYkvKA/P46L1bAkKOrRs9tGPzaclh1tlBi2R2ydd7JKF1fO6KFLvkVdzbgkYQuM11
pvetHHuNjP092A5+aiwGtFGO1f6R28j8XZV+mlOAv0bBigF3eLuJo5+9XB7pJ3pQoralFiuyx+MG
v4dR8kRepZIc3XzxmAX1uAcpGRAA7XHcsogkw+qI8IKt2tEpm47gJz5En/UXO17VrWRVcJ/2oN6s
Ab3PKBW6bygxVQ2sO1zHrjs0GfE1QEF+BEJLKotzMn/CGe2KEVMYCljOTttqSlyJ+Re/muXcToF+
Up1HTqnMAF4Oogv2ffdXBhRm3AKGI52t0DW5jJ2HP/dQ2yjhhVGhnoyHGmaai4eL5FmJUf/HzPAA
1FTprY9HEQNXzRBjxnZIHdUpTIjbeffeLVNk9D+KNyEcggtl6WS0czE8N+FOpBWBRImENnmus2pf
VWQ8ANNA3ek172zhYiKJeBEqcHATLhJ6tabo/hBTPN4nzoEDbXe0ZaCLZ1a/mRfx49TaY6AKdxOg
AbI3Po0KvWwhOSMIn61dJyRJV+nLSLpOkyOneR57RhXEHOZWRT8eUvNaTbhnZiv2v0gh0aL4S6rP
7XR8iHxhns+pP94wWDDb6p1+9tgIb65l6O5m/yoFxUlD3OICP/0x/bHB2Dt48iJ++TL63SHd3eF9
xXDW0ykAbjJXRW812vtQt5HimW4UFB/txJfzlqzA055e7rnslRD2z01RP/lTO4kbRx6oLObvZJ4J
FrWvyn5iEYEOAOgjdt2D1e2bsRiSi2Ysjm3pxK5g+FXWPZyeG6ieEj/9qxqtQJTv7U+IUqNHzKoj
k1wPg4CLJ3kXSiBsWyja6rA5og+xgmLMd2Lm3gwE+DRZogooaLG7Y7J8TQyGutAMgrKXwjbpu6vp
kAiI9ZcrovzF5PEapnWJkd/Ox83cpIIqk/B8El9twijz6PSgfqwBlTXTEBHqnfcmaSnoNC3H8xcb
+uMVkzoMn2jUGxB8krfVjwuU0DgHBU6QY/c429Gumcb3iDslc4bW0A+so1wsoM3nue4JhTN4XI7B
VpFb83iTVnQFcLkNVcQZ81jyPnX+HQvcG7i6Ay+ZV7tSnDQH19Io/jj75lrylzHgdbKA2HGOpevS
B9rNhIN3iHI0wpg5ThlPmX2W29sQ2HnQ2yQlGvTfWaaKC4Gs78Qw564Y9lLlfGxNk4Se6dDooeB/
zKKHeAgW/HW+EFIPhgiVdJO6sPWRk36loce6Slu7vVB64km61GDrkulnK3ZC1P/wbfKL+lbPIZGZ
/Koyw8X+Finp/gHaXHZ4ag1Nh6ISWSYF3dMi/eh2lLEEh9vkZtbNNpOgAr83f9SWus3OkJncrCnO
R6EEiOU/rzgnTmnHRp4aKscSGD5cibwtwWwCfX/vJRptU9wjlaZ+KNnD0CEE+u3wmrV6kss2KE8A
mDpRndsmhB9GoApXhO/BpBxW/td/67ZML/cU7AmnBHH8AdRLBH72opzAzpblcf76bcypcbUFDnRV
ecUzbxhh4hIErd/bGRbgK52q5J8ib3mds/qR7ksoMplBfc44slWMDIDejjrg1bPp5b5gm8GFrxwc
q7KNIgyekjRZF8KrcqR5/crh5YoxKxd2byauPLxwxfyYN/nmP3Y6fKdapWYEJejtOnySPRvzBAfR
qgRfIkTB6tZuh5cPpHO4dsbQnEwmmi938lVZa3AJnOCu7A5ewNeFJDiM4r3vvMmYNCwzRnu0RqYo
XGHcatbtVV+0q4WGm1778SdB19tScfTpWH3dGy5t3SbYD8pyKyx70bd7PqHfShv+HgU3TTNKUCR9
AZKuOSomuMFP8EGiKhx7zcRGgtJKPdrClo78sIMZN1NB9WmvoRAYz8j0BjSIL06Yhxh1tKlKr5ET
O8YqHefzSCtAIXgfPnGuNaa8s0kexhZhuIytlJWtKwIb6felmPUWl0uGzWuF26IoYygTsWVPvr+o
K0HwOF/lcVRLhq3J21i6kVrqPNhLiB4L9HjL7GLbRzc/x9htXpfMM80KwtVl8h2NI7OR8NS2+vbl
qxYZF1drBlJn9juqbuITCz/dzmpzO5zr/KEdoD+zXEARVgeIJtNCAoALFU50DPQJOO7Sm1D6u7Hs
9KdPh+Yp12YgFn4YO3C6/wTknOvXjQnyo2hKN+QU8+XONwBXWAuafN5EcLyJEVHMXpc4rT+I459t
NOHQkGQ+icpHR8ck141uvzlzy8ckWlqx2RgdB4CIRFUj3KdEwPMRwkLG8eFwSbCUIqaO7mnkF7C9
UeeMagy3hcTcqLMe7PV7N20urjVAs5EKSj8CycjbhWQMWCUpIpbuesnRAB6fOqEiJxGc7OeZ6fxh
Mq/A9Tv2MmWwV40pr3wG9zmXZSj1ORvGrzfXAtp2hMo7Kl7lf7unmoVTy1v+OB3CXWV/QtcjpYYq
L5mOwgoq74936+xzw6mb5TVMXlH7zgiDb41+NyiUwRJxRIaZA8DOu4f9NFYH/J6V1zxaCqW8BcV2
iTtabdytNPnfA0pT0ARpKbI8Pfr+yQwBAY2i4oUclo7nopDfgI8QfWnlplTpTDjYEbwEg0dJt2Ov
N5YQRbm6+pXcTTWddtOTBSsSEqCoE29Nrno9QEaAO7NM20e/j6SEAIrKdA/bliGZ/9NMzyzGruNv
YHpeEGXd+O+uWQw3pAII+uXwREN7+ogdbRfxOjw/4DOP/u5zOnbJB3YGxniaFVgN8hwHQWV4Bzqt
io/6Bo0XmvKVFPxSnj1EXqmwSHRNU5/DP0xNvrQbYvRaLMfrGMIoM26p6xQIcmjkGYXd5vhQ9p4a
UCBRjBhFGCwImQVr8C0JwRnyzYfIJoyfsxCiLbF/hjWgS0bZwodp15gHKKkW75ehh9zaQvtwLvmf
YpZpdu/K0lBMDce4KPdR2gWMLe77Q+WwwStfIDj2leHUb6eGr6jvjxjVncAWYzKfZ+Z+xOvwSOiX
cWR98XNp35nisk0Y+ixJ+4VK8ygTnk5t4GGtiYh0XMIKkk3B4aHZ0ydecZ5yAlZXLPUTgeIsoVwp
tWyfKXl88T8q6vxd8wys5Ayok9x4H77sTtWK+CzW4bmvJbv/aMCnNBlxhdoyYqVQCCbSEJCZEvrg
GrNewkmyajNOzQqdNdngz5nxzqIlJFWHpKRjPhyEyPWlngGT3bxAU+CvQOb/EXhmgGOvci9b2fvF
txPvDG4efxt6JDfi0OEM2tVIl1eG/+hg8qM/liDc+hElWxnmPvZErvRErlwu8VUZwu4ed9ELydwt
FT9xriUF6QfccgZF86y6Gd+5r19rnRfQDHj1Oflb+wDqpUzQhGAkgnLHYbhO5XTpI/a9T5ChjTnW
ZGPVJMOqaDy8MqZbkOpPm1a0KWavCVahpxoJoVbbAenvTVy46fK1uf9fMdHod5w7wralC1RRttxk
h41MrkqBmd5iM8xNM8fN2MZ6ZJW8PA2Hb/3MZTfMOAG4EIaJiV9Gp9wPNM4h90ku0XzskSkYyFlq
cULeCPCWINWBFzzvejW7JOxXlqzseilTNuvLzdxc21yBJPjNWk5C5ZX3MRkmA8pEDb5myOdxCGhK
G4K1f35yaBwRGkdDGbwG8rzdw3r/HYGVs4kPeE5uX+/IgEQ9Q5IhSqVSdrFgBbJAD7NtnZCZ56Vg
vT9X4HPiGDe6rB640jRr9YCA1+ZFeB7qhkDrlf/FDL0/zDH+F8I17NoqINVk38m3j18/QYieIJ9V
GofbliULEmaDo27f8XvkUFPIDxIHTmw+V0+OEPZyDGXPvGMLoFzOQ5yBQGxOH5WR50RJVybYBs4A
ooLN4/HFt0zdLRnwIisFZenrOOI63kSKwotypW87F/5+BrbhNJs9w4t1QoP5JrWu1pL+bL5rgB2h
pgWGUYLemrskMBRYYUJUNpN7XwZQGhgGWT37/sjIetASRMVWAnreCmjjfzy7XduUL4+cwi2fY8Pp
Au/A3pAYzKr/uwFc89uW2eVvKK2h2EbJxKj/kepWO/Il76IDZdiEl5pDYFu7lddP8yRMj4ZeymDP
m1WIYnHnhpnmYzLtayk0+pV3JnNOY34dHX8QsxMk0w2QOTdFbjOu2tmaSKQok1nEfXU+E0tigSz1
kEndECAH5dr+yfr/ThLoNNRQvgdMMuvoMQVAGS4lQZ0AEbp35sl4dX6MSrpPo+3oCC6DGx7ccfed
xENFFJg6T8lAI43mQ7G2WOHAaZBorV6Z2gdiV8pEJAnlK3IWKokFtRwM+IQa6pm0gK5Cnx13gvz0
l9QS4+5RomhzsviOjZXIbbqMUEyncRTYwmtk8Kj0/GgS9Bh7F+/Y2ymI39sW67Q6lmaZt2mBuK5Z
XKw72EXrGmjp+adHd5on6CEwQ1QrgVDfS3uybYTwWSTh9AtYyjxANVIKl1atMdYSsXti2GYHZmeY
9/CowSFVAZJP1Jnlle7Lz89TMGklOSLSBsFvQHN8XUuwO7Hc/XWrX9WxU6vwUubD7Ymqe+x/AiGU
IsvCSopfAtWgwGD1UlXaIViPh7237uzLd1IRKY1gnTvVQQ/pfhcyu77tiNQHZZ5XqRV69k1dVgjN
ZDxqWdCoE2niuWJY9/W1cyW268Pog6lOKbPoX6TSx5PDzMs9MkeBMhmUrBq6vnflyLcMXb7P+d5r
wDm0ojuXA5/YzF0XlBpeXa2Rhtvaedx3hWVWYCn19AcfbDYZisd1PbD/yR1E8YbLkWI+TP1M+1TG
dpSCXcBxtcdHoaOfTUb0106YlH5AF31WaNxav/WlQJ1WuZV7r/fbu7TONltwEMgqOel6L8ry67R/
sZGMTjDGXl43iJYgUg8L5+HBlnLjtqMbA26Qjnb8FJgEWp/VxkEK6SVQgML6iATbBZh+os0jOWkK
d+CanvUn0Xt/gJjKOiAQWoFn/lo9OCbfAOG5jbCABlX5Z517kz43ZY07LXXbmiivQUUHNt0vaqxW
R8hyTCdecWfSDeBR7ZwWD9wsPVk/Iu6BpFT0BlGUtoAgVB23zX5l1ZouOiKK6fspWOpgThbF3zQp
1P1+kiua06EkOPPBtC41ogkmrmrO5tDbdlVCEaqeMxdxdWtypjpSWXya8/8w/Xyzg8fQBp1SqlTA
RHC3ufySp8KRCgFIqpwUqpVHdN+0wWyNsqU44Fb4P2x+P7atfI4+ddvtWoqiirHHdyji9ckluyxx
PMjl/JDhN7TVwbhs7wzPcZKdY8ZukkQ1FyPtUCUJQC+4iI+HGZxNm3QojbdkW59jyVZGO+gF/gKK
7kblSpwGtKkvHOxw9YZ7X5RCmrup5HJcfwDeknI5qNLIF7Hg5MKtZ3VDWWI+2FrSaoKaoolQrct1
MUm/tOG2mZakszI5eN65EDgmxv31LhEan9IDX8H3XCtxW7JLp0sZWxdbp3Z/fGvH8+4agTODFiPT
omfIudcIcaiNWO8zRchYthZAqTC0VDtd2KWGI9ee8NdffZItONCjbGwen1prTyrNnXn8NvWQEWFq
7gNTD6cAKMeX0c+8HY1EzJdMOoNz3b/Z4HuUCxYTuvC5wBcythq017eTcWxPlJa9DkyCYHeSAziw
PMYiKWwdvJK2w+Z8ST1Lacn+qVc6RhKIsPQiKFjbAKdkO0C4+lEtUoCTAMVtD/O/cakFY9gKz2Mi
WnAtyI2R9LCcj2FWwqlYNF2kwyPI21oA53cN1xilSXz/avafNC1c3areYytODEyOPzb6wwytwmY2
zCWJRW48JxlVTOAW/xanjmIFVqiOC1ue5ZXOg+7Ra4HfG5ck/Soxbrt/QnRBTqfl1Bu3cnmiWnEP
I+Qife8PE1uh7u4gczdlTEuFhZ6GNzAZCTULDOPkmTS1ZJerQ3TpUSPBd4E/qhvw9TeHnW6QjRrQ
nGvJwsEIKUh6xIEnoCbHzERqiWsIOc5unDMaloXniTqQbihyWz+golOaV/FGebkKyNdBq+yDfP/o
fJ3nc24VIuwEmrIr2M2err8LuX5r+NE6gk0nNwBQzxbSNd6MRVgQh8j09okZ0zTxSJ/PDX/WiI72
DGxo6o312L0YXEAPFrwWNBw4s+4Yv10quenV9mRvm25AiBy3amFQUsemBDxajXXDncjgEpZrEdod
HARacoeDb2X0VQKMV+EFMRq3AkJjJ1NEF2w/T+7x8TsvsxOutGVKQg1yJvIIYVKoVHADzn+MK/kA
qhyD9G+aj6cNW7H3+Dz3ZTx1l9yFlzk0Bw8VfvfAKdXgg8vSRZC+uS7k8IKtXRQapDaFve0PfiTM
WcpQ58gn7DqZ+c5a1jvDEh8oBR+7uM1KRjGYERc7heuXIDybuvHkLotRc/SUzymYch8dRvNL6Ujv
PYzUV2aky1z0Q4atah0NEfb21adaRiTNErDp+W1+LnYbYqNho0FU4m6oo+1oFtbysma5gTmGqhpH
0LEvxMPsaHxUBHLwq2AL356UOJXxN5mboDI2jdQb5h0ll/LjXLmAjyEbMM3rFit6pCPWcYEWK7oY
+l7Rh5ybxsAOGIJVEqftxnou3nlD7cDTMG8rXfUJzQ2MeZyMm7Gr7N6Y24iSPCFdjzJrrs565b9i
ZOaA+IOD8goQ/4xPGcck0HBomcIcaVcyabUdijM1NNpyQ38hwerfqhLAlDqOQ0KMbFOuuiWZvssQ
Chv8wl16Jop9ewoxnUYvwjSZ7R3E93ESqmaEr1Jtu1GFkO+L0UmgkCOqyRADlA6iCVSBj/bs7l/K
eYaT4XopM9DHKknJOjS+HdYbpT/5Zsd8yCB21OJj3ZLCOFkV5cSjLQ0NTbq+ztwxKAcnBPwfbr2K
0VzP5CNZ636xVaqHJGtsFFC741VQMi3A+sH5uLaBuikxjGXiY6BIMHeUSjhS5xhsvaEikI9XBzEE
CCst3K9I7H3ehc+biuAB1sCzDWmTkulc0z5XE2gA0zNVvsxHT8oE1QjVn7Sa/90hAgFenuD7qtEj
Y/5RtYAnN7pU3ZVDizfzAucDk3DaEheWoabwt8tCe2tNKcyxh7XaD/fhEGJWdlB9o/F2P5kO0sDF
Be/XmAz4dKm4kgtYIPkE4hUNtGhmNLQNoZIdtaTxAomUeZxf7fq3vWnnHGBbQ7YNfOMz0M7mdM2L
4lN8ESf/5IvZNIYHlrFg7tLq13K8zpZjtlge7xWSLqHTTZPimb2v7qX96NyaCaOxwxoe0dbkE56P
x+S3JHi5pRoL8EBDuxR6qrV8G1bxBuKg45r8cLJzriW7TYobYUzwSp1a9ZAbqIwnrU8YXXSGy8S/
rlDviFfOBPQzLqRlaqSa3m0sV4SI8gi7LbE10oeScuVRKT5tMtUdQvyOkSWLOFPXgreOnQ2eHzNi
mxhDX7rLOAc6ZIJWadZZ4Dq7+ohvQYPD2pY52wRBCWSJph/3kHDVVNo3jB39x/+VUS0aiuS+rUJB
1wNuDMOX3AdYHeI0GCtS1SoGrYfGAxpL8Ag4kQJlX/hlm4oyv3uii/c2W1Z5z5vyqHJO7zv84axH
+yuKpVzyIIRitDLmcxktU46DtDCofcyXxxaW+tQFFf+xlmx/nZln7qEoGtVcAErpRaOhWV4/JpAn
VF3PJEu44YaFzmKXdYJKu8pHmaG2EuS0JN7KLA/wmIsZj9jHAV8lCtMx+mo4UFOb6VlUYxuuX2oJ
vo8QxcFBaYcbQ7byeaV8/0b5aid7trtLNhlDNenOmNGfaFyE+GLm1bWJC8mdvqgwWXczBLAUUNPx
SsdyUGt3QuyqglC4n42qIK6LafPzK+34xryEV1/bSuMJRhmjMZ/M7oVAVPIeyNNwatTuYHOxorls
9KzRBTTltagdJfuJ2EF7YBMDrBIMrJ+7q7vesLkJntKjha9oLrrEkdBbLJPv5wc05R+dBZ5ul9Vn
ys3PBzAEemPdu6+h9Oo9Up2UHDeR+oPs4Jn2JFWFvAwWWb6sEF8r8QiaqBCuMQjLb2SJq3htJX1h
4c3FBIZjeDwwHX75rIRTEmSxZQEYHhPo/hmVphvWg+xRW8AS4QMO4RV221L3kKSKZU632/cvirv5
v9wafAGdP5SxthNaFP6EX4WgPXNoQoV/8nYia0BYGNOdSt+cq/X5aiAwHk4zJ1d541bDhLXYn2iN
GFmJuPxE0xAglVZwwtd5zCYGHGHeEC2FXsPoy4zUOlMLEOESO96DnjwwdAWzhn+9kYDMJ+8JCoVY
QIBq3qhxzIp5INB47sDVmta/Lv3yGNVQ+rDCNWwI2oG6wqCebypy1k//U7DK3p6qd2F9YkJGL+BZ
LhIkRTpjQmUiysowZWaiM7GNjvgv+KZjJsoOtEcNc64RdDXpY4SLe8MsGiUuByz9IDNw3OaYiO7/
kjRSE2d4RsX0jFuRRE0A0VOcIEJHtrzJ8Qwng8Sr17EaP02/zFye/+TE6UOC3Gh/02CwMMwS7juj
4wwgwNy5N9aELNKUTOz2vI8bT2DNFVsAKxkEtryUdR1HYtpqemg5WBeO9B/SwRGDv2A7HLIDIx8E
iB1l3IIHjkTZMuFHtVGPxSjNykBPeCnJky5VsWwXTDtUHydCnMEmWsUsOpZSRy87BdB8vq04MN6R
GFIJOVRkB0BBLb2vdZnnOILXI5cDZF2ZbHcK8AAfM105TnI+rB8pdFNuMQXWhAsLoGzAt1OFK3j1
YJBbkAaJdeeBRoVgBLevPhB1fMxB+7ji91BWV/YrvILgrVn0PJAt2MaGqswo4f9yz2+Rr3dR+1lf
yHQmNg5SzybnCsbBlGB/tS8jpERhyyA/zfZ1qF6+FpL+kDE7P7vA3kWGFsbLwgWH1Q7DVSYEn4Uz
yfAmR/Sihsp7+VcAOpr03Xq+sTUKmG/GGn1DO7NUudgjTm4DXWpUJ6JQJ1XRRffdPtCKAx55Zlh8
aJImaz7+H3KnyHAgcruqVsTCMn05G7xR7+UiadbIZPS/50YHuClsNFHgt6jyhZI6tg6KUXbHXt+X
IHduGAKE2HcCOg01wH23jj5x7PNT0rieyQ3UI3qHj03rb1svj5Fu35GKz9TfhJZ78h5J6wmE20q8
xaI7WEYuqOrRBSCu6EMCeWxSBYA7tbGoV2O0esoj7EhzvH95C3h8+qM1bSZR77tN3EDNiekzT2ZP
TB4vnecwvF0Qq5Y8QjKT4npCqV01XhsiUB7q/qqMwLty93EkdpnchIoYTOGDoXfllhYXJ4liBXl/
pZXloIf3FHQMoTw6JW7nzcEJcpeMLnlVQfCeIhUri3+wjHDwvmFZ9lfjSFqPH5w5DvKmRH8rbv1X
PT97Z2vIKy+NDOCmcaU+WL8+5EFshaUeTyjPPJ2xQO+MOcwSaBit6kdPghVSWXIqkss8Yb0MENth
BztPG75pEJvepm1u1WkQ4YWU8zRTF56dqoEfVDBl8JUrWYdEViz4DKCN5ES6mrzcDNkKx7MHd1it
q0XF8X3goi0zt22NFMZg0IhUlALzaCNz0D/rnXb09yW02nM2eXCpvJLcME2xTLwB0fpDv8bUcal2
R8/3roT8PyeGdrDASEYqW8VFbTtnLO7FjExpQntqtovlbrAyPtuBhSaJPy4mXlRjlwMSQR+nBCXh
nMzIyit0SBfZki3rr3OdcuagG2+Ea2yBsS7CZ3AcLykFVEOTF05aMn2WqWnREo8qGzFkNXtYI197
WE8EdkWzSzQVne5xhvtVe5/4hh6BNIpuDgaEnudHkT6Jw+S5r8HTF7G0MZTNbUc8EMreDoNjIiaR
kRxtr1bIl82IcB630hnyeJ8fgxpEXkjBsg+woIq6S4O59uYm/4ZmGfhXj+6zLrGk8pECDwjrIwKu
f3BS7s5i0QEYpOsb1uWyxOL2kmFPjNmM1mfm7bmAgofbVfnQkmjKrw2lBUfq/3vbslKH3O7Epbmw
4UrU2NCX+2oUIuoM7Xk6nxsm1IiYaBcM5mFgOv7634cR6K5MnF6pYHNA8vid9cMXaC+EKlpFf6vF
vSHzm5itwZQSFfl2rojLTi7ZZuWhM0UO3rwdzpgUml9Q9mGMz52QchOXrFvi2skY2Z4+zeIJr0O2
huxmCOdD8CAf7UXubB6kMnF5sH6gjh8aq83FRuhleWT2xG6msiRK8jkN/RvT++78y/6rwGol7+T0
cePty3ngTmS3Yqr1vR661JH9Pc9NN/glmLiAqu7SCwpaDaQjhOja25klEp96EOqE0/9wgc12Mssq
yFGVbjdDxDTp2kuLOhERyBl3S7rAqHq3UwVEINGjhOtLD9QfSZrBSQh1Lj6gqyuGlJbrvcKmDnYf
HEzANQPRBuTugpOK2f6SCvZ0J9jmEOOgTu+LVXCnkBE4iBHT/KiLHhKPJPVgU5Dem0rSALVhwTIx
gABaK9aWCDWwHHkCLsNf/Ltd4zXQjqWoaZfWptqnNd27/vWzgIQDIsVACHH4Jf1XujX/f2tOISpN
2yb2BsWDsmOAusJLVtOmNUyKqzHYwUpsEddV+wW+4G1MNN9O/GXiCL5EQTrRrOkNSqXN3SOyKOCA
l6ttO4HyACdZq1BuxZv4NhuJXeQN9MA23yevdP6gQRo8+HOjs7Ak7i6hzE3k9x5HzW+jHf0+AAP1
QpcerDKMn5J+OjfvR7sbS0t9reymxXofhqfH16GrUrsbHHbuw4M1auxEiiQwrI+3RsSO243b14z9
pyt0e6mCGv/8v23pgR75vKtoNXirLz4TbyHv/cNmKnQdb1unclkqtWQQ0/2hpHY+UXpOU0HnyuNh
MF0wBenB1GDBrj27NUkrY+Ah5DOGpQrc1EcyWzIBszmDVe/LLRmnBK/25au+uC+vavGXEABPKwvp
CZGtnO//DS/wo7pHnUi15GUEZynDFvYp6xOOxMSbPNkC+j9OfF5UMHs1EkhukktM7woq2Uc0jV77
r/Wb43iYa3zWWkoMyC/P0g5K/BxlHhi+EvKoalPBzSCs6rcSt03O+xRB1expiR3XyP/mPW2MJrUh
lYRCsPJKw/oco96Z960kY/nTtIcNZmgcFYA51GsnKvEsSzTT+2hVOjXFDFwQe4iX9+SLrVRA8vnu
yRvnMuxsPDdcnYedsYK+o2aq5JU2OBSAND6xEL6gTZ7I29j5WRDdsg55IaliMo24xniXD3P0Fec1
lPQ5qZRyOF0mWzY9j6RuckHRaCh/iAeVNo30gGoUvOjh/mrsHC4EOCMiECTMdmXXltnixdEeUQKA
YqYNv51/Ycw0DtPXORTa2vh5BNCbvoHFO4Wh541LyFDQN9AoOuqSF5UK58swMiKh/M5s0EbfP13+
HxrqVgmNp6ob9/kJIvuyqrNeSaYU2pBTARA8QX3qg8RQpxHh619a0YLICMTs84OTSwjHVJgrPL38
HOKS1lkVj8wSI3QiPEn6a+nhtu9Yrs0GBz8F6XSYSSXKXRIxiLmDLH2ptGEDWj8V41U4XRk8zrff
/80VL61fDY7DlarsueeFhNmxIBmIyLgj6FsUsdehp5hgw0AKLkW/0Gyep/A+BbcEBwvH3QVfORBn
MzG0Rfu0+Q+5Mc3NgkMmsmAQfcw8IDsFpbsbkJbdoZW58oJzHpBLmahuAkmac6RWjlndAjTUZMWr
otZYa0uIyZmB1aleSPgwnVyadDu2WdXUBrI+bplu9sE4d97whSa3bPt9BfVgFRj+EIhS221OjImk
KFNnI+DlGbMaS5MurH+7XjNJPuAxCtBi4RcORgMFc/E6x50pJUT43b+3UJR7Fg7D7XarMff29vBu
EClRAJrCE+QEigOl/ptAR0yNJ18iE2rkO8sKUmajWpsVRNKfzXf4WO2LKfYiZGPJPyllzCc2MSFl
5tkJWGHdq58/LIxr+58Z6l8VuSDahsa9jwEBJWbDFWDHEBbILBiEQIrc+yrlXO9KbXxjQZspuVsJ
rYXGd4ZAwEGI0s2GvK/LgVKtKR+GcsoJ2A3JyGMaXZwl3fGdX8RB6nAz9WAvmmTUw3zi2EYqCont
kaFmBEFEhQ/rzhHnokx077bLXF+l4GGAd15RihqQudnD1kuCGmS92lan2wB7azEp32V0wnEUFEzr
LbLesiRW+rFjqQeU34pIHOdXq25IwEOySbIVxG9QZsvsR708dstVa8utEjZJ8phshbEFQg+5drqy
QaWjxH/9Aimwte4CZKXgordNT0wRjDOERZ2YK3NmKjEklQw+pn46neRlghk7HlGLIwP1ZHp1wfHb
b8jbAdx1gFAXCWM3HUNy0qJZKHgwmKubfjHc70iXGQOXXmkIhCqlPyr0kyJPMZRKQH3ku8oAY82c
xUDLUMcWqc9brlzQ/nAEts/tQdsI4iHUil3Dohuzk7c/YV3QBZPLPEHdFHuCzVaQIfUBZsqh+WUd
DfzzOBfvqS0pKPVaAYzEOcQyQxQnpNN7mhLHOhbS7LJuo0rJ+AYH21ViyDY9TcZ9NoOrRl6gnvjx
ayuP1B71qCa6CZ3OGLmNIHQC2Hj3yZFGPOPxz+kx4BafJDRhbYnS5v2iJw4KcxFLZltGOPHuO3vp
AeCuo4vXaZr7qXKkJt2znRoraQVLEYpraQ2E0CHe6rGbgAGYBV3MHo3lxJeSrE1u2Nvikg6UANhc
Uycr+TnEo2Y82iKPDoucVBJA693Cey05b/Db042SpSsVLpYznWPmq4dQEbe5LxjoUIIBV+ShWATy
VTEWydRoQkRX9VJ8oUvlUjQ0ikWtuE73dsdPzmNDDupycrjjElVwKZKEO7vxn5sO5BQZ0IKRSpTk
KbADAQPwzYwhJcMgERdZ27toDUUFq5n6kKKWj1nKu3IzpdaNlAi07y1s9ekT9WgEPasDstzolZhz
BmXlSkfQPt9nsKoB4VSJJaWzYYyisTkBWEnkR6bFp9p4VgS397L6MzSvUr+qOdazSOd9Si6RFcEt
nYZGrWwGHjbw+LFiy+pzFp1QTfkiebbF3/MzuDXUanaQ0a9TE8QC16ygCnK9AZlxceR5c4EQKNhH
ufvM9TbHN8dzYDD5JNcIaeGFYSkq3+aggyByjPjvBoBhMS4v0EtcC2ydjHAX2goxN29PxXVugbPr
dSvsDTSheJC1H4lcdH0y+bScHW6qXYyWscYzbSUh9IpVCvA5OWDO2YNlykLpbBrF34Z9m8Eviz9s
SPhWGq18DiVZaAEa7qC6yCBcpO3FgOamW8In7lVVNv0qnMMo7ZzOfN2zGWym/W8IiKzPqVmceNuA
Xqkqv4iZ3GZ4raGLM7y+SEVxW2n90gR6zGsR4CWFR30W77OAi1SJldjetrAs4gG2+5UOuOcERNFa
8pmtCbgs+KD35wriIYEwEUZ1g4XuXRwcKwLBJzDFzYgwswXdLBk/acCY9WUsu8p0oiCGX9UIUWTM
SnqLQkUgpMaZROL5Bk8JdkUW2ip3J49WWphUsCCAQmcd+vPJnhVCWKDfH0bo1XTe1ZO0tuQvTiRg
hXV+3YOMdcOyjxuUvcWrsLX3VI79WdIdTbtWX75L9qOcfPbh9uDEmRL9uEu4jW2OoL2HHGCePbcs
x/kMyBIMgFSpMCM2qLCr1QvbAPPPpAOaBlHkvPEs5PSL7uzTnGWdWgPD490zhwEF56dwyszrNJnl
HDMqbQv2neurxRlVPgKE7jIhi8Sa28fsfyeAuHvfG1sux6g18/7WenSpMoa4oOjBBf8rTjslpdDm
ZZZexYBZPTAjsQbytr6GX9FoyPZ2oJ96TOubzycSPFvJ1V3Wu87lP1u+PTLIMKhKoFHTlrjNS1yy
13XqCO7EHJRNfVGGeQwif0YESF3CeCV6o3zEm8WNFy/VDDEvHIRotPYR1eZNbnW6izGnb+hnHjlu
bM2y6JSJi0lcD+nO3WheNd1J5VPlUTUlctqCT5zuqxsx8d7oOZXiM6h9VYI1fvZIfJbalEW1kpmE
WKcIEnOC9esIN4KJnKOaLLITXv6wxtRifqOhJ/BsWl2Qb4ZL3wtolExnzPCyyqh8F64lFQ1JihRg
bhkNx0P/41X8WpaW77xtOOny3k/3f3wzKrNLg1idr4o/hIXswreDhZPgeKcSMgKsj31kbE6yYcKM
2Z7mE6edFy95vCDrYZdKfehh/CTwNphtyYwdQKA7xcTu29XZqAZh9afxsnhXffqdsZnVP80ipe9m
6XrmZiwUAudDvduuqO7uBxXJMbftBfu4dZay7QEjo8tXI0nqMfPn4oazjEuPK3RZj6FQWhMcubTK
DBWGFDOOG+9oUuttzUEySJoOBtsiAmGQTf3DgF4W9SQg6Nvp8Xo3Bs6jlDzYZUz14RejVfiwhkdg
QZQPPYRRTmFBLdhjRVEA2Tr44yiVmJioP8pZxgc1DRzTpPCssnQmdFYgKfgafH96yEFpdH4C0GCy
hP+nKX8gQOBYa4QWUY7nf/u3P/eJ2UPhdaByDwXpAx+w3TpA+1PkE0LxTL5MGgRaoc6ZJfPCbaMd
+rBYxfT54YOebAohQcuBNMfXalcg3LJiyL7Q06QoYyocy/fWvun6Bfq4HY/bl2qPy8MSTSHdi5LN
CjBQWSCy6vu5KCpqnDHEXNlcRZcPMNGhSaxAl2JEfZhO/x4XINGa7bZU75CfzXFHlMXTnwlunmrM
sRYIpxyz/e5wB4kR8vwyoFWPCFaCbRegV0yX4wqeLuzVt2Z05McVPHQPthGskrdPC6blJ1cz5liM
NTBIysyRipYlZYB7q1T/V4/SZW4/thZ7s/AG2AyNlaSTyufkCTLt4KyYyjOOvHT1+W6Io2BJhG4S
4apD3A/OpFtH/ylAAfKmZsbWsN1O16R4EFOEJ1Oiuemwyf2mAaBVTwvtuJIHsBXMf9vAqNO3gyJB
v7BWVDm8LX3PtIOwPP1UxPbM2COEA4mJXngODgjmAVHCWR9mJ+KxIJFlUfsW/ScdTPlVIGY44caD
pbqIGm9HsS+xRXRSdkX8VR4Ss2XeoNOEoq5uqy+pnTKz0yTWLm+62HvU40n9jI1nOn2MROzo2xNK
Y3IL1A1R3VBC9Z2qq+EF3wsi+tg8dNvUVPvln9VFV10tMRrzp7J6qccLZMhOl011X8qz69L5Jo3D
XZleH5wZe95qlCiT5qRy5Nz07I+ybSehoZPfePAM3ppDfEj/8EID5aiSgUrbzmwaJyushLt7Zk9S
bdflq4eSuFGOXHORApz+EUgVrc6kNC5Taj9XrWd2l55F6YXdw6YBaifpTjVgb8NDLOew28dzgb5f
fbGSJ1hrSwB3fS9lHJlhyh+U8uyQpc18XtHv+fKq37k0kMcCr5SVYpOViJgXqnyK8xQnIonqwxvb
x4/LUyuQyJqeq2PVN0G0yp06kXqXXeWHiw496AfXisjZgeqG0+xphWC5uP2on9Mqd28WQyyIzX5g
dYR5/7Uku52Emw/2eKB1bfDOe0mbbme5FgnLDFgtbewmqZ5Y9WV6YSi+wx8vzBDTW1yImTi6PFKF
0CV4dkveZLh+JiLnCS0WN/qDCWduGUQz/fGc3t4lJTeNtRrgFou3dphgnBnAZq4P4LQu6BLLNwub
ETJXX0+uSwxzmMYq8kicimBMd2I/POWE/5TD0PpGR08lEeInRaMs9ytmAG0FuIc4Uplj/gZFVRTO
GoLD47yeTtyUFX6GiRcdfoqrEQ0C/+ODTdwGzcZoHNXuiBWI2JYC4pROzSgMyVOu8a6KorQSNPIR
tBe9n6J5OABNDCMa1VNQMUnpSb3+tZGrv1vgTRZhfxWMEJBFjLOEowNXWk2CO1hfh7lH97AcRt00
fYNn2f3Ma/cdUkNLTjuzEtdVuD9Apykqm6FiiK/v/5zqKJRMb63+BbvybFi2lD91S6BJ4fPrdHf/
8HUB8VRuZrHGslAtti++7Lh6aYW5IqcXTRpRP7Tz/KhPgaX9M9g22jDJKwCxpw/lGmAgF9EK1ESr
W5YyoSGmwM5t5dIfG2IWdu5d7A9Mz65bw0DoKkrKWGw34r2DBPXuvyzylYg/bHDjZe+1366C7dKB
VEnjAuFCwyno4igqj6RRXW6jDTe8ccdyrJl67fb1UmepbaUEgxSFKOQ9FB/bSkhgjaokJQpnKgF9
6pHtXy+WC04I8rxoOoWu6d+j5gN4JtS6Hwqxo5cc/bJfSi2Vqk5rgTb8LDZUTofAJuE70RDFbspN
GxLwmBxK93lqVsHvHQB/Ryh6PYIqj3ll4js2xsHe1ZzkBsbSqh+0IwSekdnO8jTDRwjT9QMLxYtR
xf7eUE89tQ6qkTLXgubwhGq9b9aXxZrYAxoeGHHs/ybDlglWIIQsyfe89nzz5hxMLMKaojP3JVb6
P+CNCzRjGdYUYFQNRpI09js1MxKhusmo+eevZKrIJEsF6qZeFpk7zgc98EiSOpdZnl6cVbF2hMMM
CKbGKAT47rPKF6gsogMyHaj/HtUNop19PYQIhoLvp8zX0YR4D7maC4optxjO+Q74rcMYWIbAdMAf
aNmdSzVjUGygYC5LUzI9+EnkZScfh1h3EoZUdOvCxO2wvRTuSfRJPBIYOo9wYfB7oVqqV+YwTbSa
LY1dmasT+hwEazonMxbpOpH4l/Mb1/5qsgMldyWe0lj22x+3VUAM8zR5TRq4MTcNH47RmHgw23zT
C2JR9MmCQ9Z5iLdqEgWNy3eX66Hkb/I4+puihed6bIKePSRnUQSc/562l9pwBgUFyWXiIbIYEmzF
rVykopwN1aZEFhblx8ASiS1OK7m7tI9y6KiPDBAPTVZQO10DHtyBIeE/D0sKc0LkktDWPD6GYfaK
gMmbTFQQt6hMxb5K/mBu2O6oDhxpjqu6or97S5AA6nxtSPsUQugHBPyLJNCSUkRS8VY1OwVXFO2s
NvaM7Lf1GW1FQ4mPANPdOPu1Wiema9lech8fm7n6/Q3nQyA1yyx+Hgxm1lclBjVVCUYQoevXWDPl
uB/XHRhvSV3wp5Ky1+XpLsfOWPEq9++kMMPFWeGch2OP/k7psqA8pgnQuixvgQzj6IckHo8KwyCx
mkR6uZNEG24Mc8qN3A2/68hI47VBprLSbNzRUljPzPviUnegBvRY4t5BFGei1AKZFNJWcP1IOgeJ
nnrOL+AHaoJrBhVrq8m4NdlmLM55Qvg8yoKoMVWL8/889m4vp9RmGDfH50jm5c3Ti5ZIgT7X2zTA
RP+jkaeMzjTUYb/KBa4CrlTTQcIJAqlXHGdjbdcDVq/Lw0j7y2RYro6qPlZeHeJYE04/Lb94SIQj
QwqpyLSXFuRjhS7LgAqPST+9JtpuBtzhET6k/seOcigRp8DiY8ICDekSFvVdWPSJ1gk1DG7NLKTa
dgOuQDqJcMc7PsSzie2of11mPiYcK0/ZRl5MVcp8hfJADFjbyRuMqE9EkcFfpo6PKQjgnJ056/YD
khTGG880YL+33mMg7nWDx+895FYfD9LGhMqBGgE0fQlNY0b8BMNQYOqickvxoJd4VG2jZ/99C4Av
Toj4A46BJwh6AT+7uKyp7tE48zeOuuGH1/3OEYtDkHy0BkNRRdTia4Y1xRG/7EpzVVDt6WDABLJR
KYsrTb1trfcosyPpxrxrFE+IZYg6s7rDqrxo9Lz6ZcjQ7mTEg2n7WvitDa9I2cGJh1kzchMtE7V2
ujz1q57diRGrJe4G3O+LO6I0YbTnNNYvXsK+NbFlnq3YZYuJzz74YsuU++YLVR2hwNaithKeynF2
AluzLqC+YaP2YoVWU0KfllTHLfInIoLk72vv/4wBpagJRtK3rnw1XZkQ+Si91r69fgjFT6j0NOvs
er5w5WqvueYd8EOI3A8iCQjCHKGnszORW1kFiGLhxIzOZFtOO22KDGQ18njAP9P8JIu5NDlvYgYd
joDtmm0Naf48yzuoTQFMrbvgQgld5iHc04xhmPMAqKmvdRshrCxS0iCf0pf5isg+asFYoSAZfFTI
wOZEz1PnACNIxkKvfA8uRmVNm2cfMPV0b1gBFqh59C2uIo/MHYFUE9k8dtpkqr0BLw8qId0D+qw2
8HpPFM4qNYm9dasRJT+Jdqs/uA/3ccnw/DMji8dAMYlYtdtSWix05C+jX9kvwWG6FABPtUEOu6yM
X98S0B+ha+v8qAxODJHAlFzaVA6Dxr0Bxo9gB9tw1dLhEOTF0a0X/b6xN/2GQvpf2vVh3Q5Vogvh
/Rz7ymHkgEXgaoNJ2MXz6i7rVs/IfkpNny1VxsqUFb+/oa2CwSTrgqX3kKu4Prxm1SB9Mv2rtUsm
7knN5ANVCggiJr2rtRtVuGZNz/dz3OSle5LrIj3rldzHt1ttqKbuQUCW9hqAeMla/ySBf089X9DW
hY5Xaifo7eHTmOB+zM4AHKJMVkmPqR6fGF45IM1/aRjqSr8maECeWbJwy5Wxlef6FND5Zb29mYyy
Uso+a0Yd2Yfo/uyH9prrPYC/ccJQLOqycGB15tSe7xoWVGcZNxteL5DzYvECb0AQJ7CAsAdRAXep
AWe/PYkhGzPzrmnOFGbPcQltoCWPFdSZrKlw/TD4uGks3BZ54sskCJIDecTX1lLyohcGaWL+N24c
ebFRjctYnaja2i5mhyd8lehKEW9A1jWYgP0y3p65cbvOOMPvYBmy1nMIOyMTa6vHGPsH2GCFHAQy
2qCS3KAMjWg0CkwuiPDvgUzVM7BeWL3CmACdYGAko8to6tYU1KZBJOfzm30wbbTZ+AYzRMDzwDG6
DQEC7AsHjVof/lw9V9sePec0ZZtZbRu8dIo2nkrh5ynFjqNLLehl45oEBAbpkHZqzALG8EmYOXGg
zfQRAed2zUF6FnVrP66yAYlRW3jTtkZZrhv+AGlVbRbjwcIhhC3Vp0sgXjMRaP6mVA5N5ccCwQVL
f950PlVsuMNx7/jP7W687UUfnCYQqs1C61aNodjSSNmcf8NE720uOY6E2NIZPqdq36TuORklh9g8
/p0Ijp5WRNb96Sm04k7LsoF8nlTwa94/+x/mikKfMkN5sVl16AEtVXJ6dcl42lhdbIve4zlqxRzt
fqGhmKNHgglIIAIKSp4h5Qbf3W+FsCnRhm+oFqMPuND18ZyDaUhniL6tM3vohszzXScJ2wXoY4AI
z9hHqR2ANxR0uaJZnCXwN9kQrfmfFLHqiouGaIpdS59GMC2xZi5+bR0earHDJaKD0OIaXzAkQu72
UicxQvaYop8ZNPYqj1dA+EO0D91aYGMyuk7ejLlpU3ufrS7+YExNroS/XP2bbKxxUaSGKQ0CnKEa
cvuyFCAS1n9ufyBhT7FOx+IO5D1v3m3R0RAP8Qe3AVRDzxWbSgsbSSSZ2DGeQUa+yMz3KeEV7frm
5DuuFSZItVGK9XNH1TIDK8RboiQUMfKVBePgjjXNFaUQR3xGZIgS7Brzq4M//35Cw52H/55uPpGa
slpVyObWdZCwRzkqCavz1E2FzXNNetQjDpEf+ZkkxxoaevqMNj3eewibW/arLoV2XskykxJOfw/Y
SUwd/3fZdOOJZcUujeh4dyN0gytr567v8ywwZah0xOtex5qu2G03zmkj94EnQ9wqCtYewdxqbY9v
pgw7ZZK70pE5EHV9eEEZbjOCY2OAqj9/B46clkzSpjLomvhNCoTFfX/6EvFBIB6BaowqjiqTIflq
jExPbQAXHzXVkRpdHl7+PKKbvrjvC0Z3WubMxp/rrlkkpEgsi5ii0RWuDeLJlguo3IuBAYnETXx0
6zYkdG593yTs4NrHFWN6vdOyeU7Ro0dCJeoaAPWLEuYUSoybelj6aoo1wIFycZTmWbrnKhskv3jW
d1PgdkvGqX+5i/nCH6NaCaSS8pl5AT6EDVVvnlSoT3uX1A85oYne5RnLdiGkhpLMqyKG8hYEeIyk
NH5N2f0pR66qG4M3nD14fhILQpwYxiBS/lFhZdokdDMlnnLArVEYFJZG9SMeh6WAxyysS43cgc5i
4TmXsqlSm75Rx1/UEwTgNWOlkw0XgxdISzJj127KlYdGIfySHmvzqppWzXCqdmFSomyPawg3HEUJ
B2LqF7Ju0YL9f3+dLq1Kx41LV5nbrDT1I6Z9xDHGO867Ej3/AaXAKAEog2vY3YpltktY7+Py77aJ
l3Azun6imXUHxIxt7W2JOFf2yXU+lxXcW8ZVDCwunSv1vArySZUdEBvxb7nbVxuyaZqFFkzFaddW
18nbCAV8sJEQGE+Q+X81DwwHIRLSJBtQqr408uijdYUX3/6byN5UfB6nwKUPvms72GvKSr5yKC55
ZZUFnDl0twvx+RIqOH4aVK9biIe1redu6ynMmSGPoB0pHCdMkF17h8ZoYHpyms79IIZV78xVSCfd
fKgmB/gzXFFs8bP5VpNBHuiVnb8OA9SURKBSChrMKcmPg96n37vSjQeM4NU5WsqeqKZJrUNWK9NE
5Hq2b9f3jPusCm+uClgSrKkht7TfO4GgvZWvLvKOJKygpT+fq5Fp9DMvKAjVmB0yySNmTe6DHLlD
0XhrUl7VR2aWQhjjvsOqRtPLWjy2YzIS8q25w4OoCo9hyAyCcHkQePsJLnDqFBTYud16+M32Lr0l
dNosjcGVgRQwvGLbufq3xyZRVm4QnJK+sNFJx8NNw41xcAu1TwsvOh0IjdI2dfaltqISJtLQFJum
sXxRS+SGhUusb3Lsx7/6m5DSFIWTpnbI+nq+QyzP/36NWTJxXk9u1ONPQnG9HQXQQO+8TGoBNZLD
WvGN2/m/H1Q1uTPoZ7TXUJ1FJw8JeLFVd9EgdeUicS+SWPLZpXQsqAdYorw6G5oZfapAgHWDnAXX
3js9uCERVQXrDOYAm86miNUwAtZGsYXwl0krJNqzUCDy5nROjyw0YbRRX0IL/5P4urrbjeGQAhg2
xT2xO0yOiijgQvdAv3dcSzgz8sG8HXdIFguboxWPMB3FDJQ/Dwpe1SDSBArcnvkswo55okMwdl7o
UY8KolNgLuPaM7iRe0AQQt+ONY7puZj2aOoN6zPwdTGWe44PRNcemDesV1De98ZPI5Xi8Qd5BcVf
nSQ4tUH8Hd/jCPR/Rotr7UIDwxKmQICyJ565olYRQdzsWT0olMSfwY24zBxP1oZTJ1BzA5zhC+M+
oJdxe+qJe8dxmkKpR8tmpmFIqPW5McWt46A1A378IOOTjSzfSwDP+s3YNJAcmn5jiuGSdqgBk1gY
EpohqhmtUlFEan1u5ckdbOKSfgvOZQpgSLvL7NCmjChohzjpCN+N6tN1NXJgSXDmsyuHx8jFERfP
48tIJNw3ufJz1tkF/Z7BBnklr+BAUzQua75HHTBZoGT0WbJsGRLXdXlOVxsfWAMsNSVmxbWwomXt
b6D3XZnqa5MLqIipvPzCZpX/FV1iugJL3jMpqSb7FX5JV+dtlyWkQyfJoi2IHFysWSUP7ZxZBJ6L
q/QzuFNTpiPc8lyIup/V6nZ2V5yMCSk+evefl9dnLefCjYIwqN3NWzyQp9f3O8itqZ4gBxB7L1SX
CD+4rHkI8PWma3A1Ea2ndeE2FbnY+7jEDGr6EcB5TN1E9vf5yJ18m4oma2MPCIAfLHUBdcm7KTI9
/B7qJc+lb51H3/dg+0b2kdMny/zSY5w4LrgTRdp6IhV/4LXZM0fkYoP3aEJHCsk7fTekeLxElpgN
wq+dQYnSNvbvZjEmKVqMWB3qXPtLz3E5eYzPLyZOSNkq47q0dEJCeczIiYYlpXAjSc9PCmhD0aVI
xZGVYoGOszMl8b+Emtv6jemzCyDzzyfPY05utYMpa5Mc9aeJyoz1OkD1sAsNDhi3udlroL5nN1AF
PrD+qT0yX9QouT8Bw/mk7eMtE1jSdGd9Zr4OwaidD/GXTHU7eEtct0KZtwrPapA8b/JZT9wcf4pq
DUxazNPET6s+KVUZJ3hQouYr0sGbarrPtjGYqB4fLf16//KNupXzAu+BdKQFLNJYQkbcGZoYMtFX
Cm/M4pVtmvHNZycg03Zb08BPWFjfm2FoTjVydwBYxOMTp8npBrwqAe5HzLeUeYeyq7iAtAs9bHHH
cMLXj8JyZTnzsSDVsm8VOxbH3/O4+M5PDJiUFp3+11qF3nxQbj3LgsFq7iDlfgx0FBIMFZpS3Fxn
MCQEqhWeKdEHuDZZBaIYOG9DSe6jTGeGdfPlvftO7VBPoR46HvYnvcdx0xqg86fNc0s6V4cQcApg
GhTpQ+T3iEyBrgvnbk0awD3LU2HmdT5Npb4pmj9AR1xojUm7ZaFhPWejka0tcOvLj66Qz99ZMdrM
8DNT3jZGAFNentSOpzOQzHOQMya4FnmgAFHc5LsKINwPAoI5S1jDOuCPaIrk6k95GMHFK6M3ZVk1
vRrsEkn2vAeoo6IkGY5OSuXmReVDdI/2vYIXb0Af91kQX3EiLHOIbo8yMrRt17IbNiS5Xd28MhZR
jyGZdsV16z3Z3WF+59a78RxT4m9DTiAlDwPtoY/tdPzEQaF8yRjnpNkjjh9PzBeUM/zivohw9hp3
GKWeqgdYyDlMqOkBUODCggNEAMaBQ7hDng2OdwAXTAS/OMfKAgmr/3w1b4GJSAqX2bl/wFBCW8DM
2DCElgUz4Weirfp/1Wh5yUzTwcNZSybIhXZHmpM91nsSKxKK4U1x0ml8Ipa5FqWAqC13UQuO0ahy
jRuVHeSKYG0FcFgyiiY5N7hOvctjioSxTxF1RDQEq9JOF5ETzNcfpHxyXQcFhabSMOV2KYgzRGzr
FTq0ZKOr4aVo4wnZp5clhRhVtUjJeYsXJvSE6WHMM8l5kHeJr36naLiZ5knaY0taatFo+LGWG83G
IeeECVLG63FrW1GYKk2PuHrS3JdKFtw+ZdW18EFKo2eV1rzDcQvsF8ZMGp3nqdyJivH3cP9omZj2
rcb4q42umU2edILzPWpPbpWyVoGNd6LsisxH1uiG4EAjBFuPjGeJzx5XP7kUohRGF646p8jlrbLL
iWQm2uOjU1sScj/PdKjbMCOnMmfhvM650CIDbtnI+Gz9spr5D083m+8+FgRvzlHz6iPrKLEjAb1u
sHwsQMuZXVHKm1rHM3hLxBrBFLgnSgVEWhAQj6JSyix0jI3XrWHSC0O3E+8TS87+mvpJkhbOYadp
Jn6uAC8NZTKHzDP0w1nb4+55io9evKWbLlGCqGWYX40n+agpdkN2mgMqiQkDjOVJlD4HTL5l9mFg
qPR9xLjdzabylYSuKrRzRYXFgOJ7lcjO0rukdln+MF22yjfbcWAdu6p9I5dMUTc9IXPI3PQ1sHWC
emW/irDO4ORLqzkGAdpfdGAA5lUyDQiSn3zsc5TlKCf7B55D1BQJRZBYzlIv1PEWmH+iI6R89TRT
31vcwqpP+EmNvLkr9JL+uzCK9cOhjhRcTAAKYAEo1wT8LSqi3OULsENlZ8TXDBtORzDgNQj11+oI
nTETPULxmJ9phjfhyGaoCvAWPQ9neLArw9qAgryU57Ru0TZ9sURweMmht5OQrdHi1hgisjjGmeig
rBnhk8iNq+QhVGJWihj5ruQA+EGyk5YUyE1CLW+GjdUUrRL+6WDZxhXtHm/1MKfAjD3sg981atqM
UoXEnL5Hf8TxmRx+fB/k0AEeixUW7Vtu69aJehKb2mvcGgDjs1dDLYsU8vQtg8TngPIgLl7TB15r
QLRWVzvkFNgMV/Wks1oGldL4UOF7j22RZVcjAMSBfg7C3qWa0+qayrhfvwEoGctaj2WU14IBv03i
JedCzL6pZOub5EjX7UpEw06hIv2oMumXqG7J04jeOpr38ueJ2WuiK8kTSTYnqQOCqvYk33mXAhJm
nQFYn0s7IfBs3wKatLzRGpW3+85zUC96ZhRwEtb7bUd90poICYAk3si74AS5/ta6AVQIIo5sy/30
ZihrMe3kGf4YZSCZRTn0kbc0l6Jo20vWsD8hSjeNclNuG/OZJqmwYazHi7SuKI/bJzHPnHultTjt
yEuldmZcIl1kAWnaxzIe48L/9t+fJihSWoKj2kRjnI/6Yp9VrOIW3Pd1RG6AmQJKxz5m4P0TLyFH
fJX53CsSvfGuxsZ3Xop4iiDvaPENbkEb0hw5ZDQ/+Zvo3m7KivbkAHs9VpqKdyXegH4Jtnc/v+mY
Gu9fXF6Ut+WYk8uuAk9ORKCsX2R4pq3DIkBL726PVNaEH4vs85YE/CqtbVFDmh0LF3/WlMcyFsVW
sv5NeotFW7ZRukRhDVat8kdDI+MNVGE1LAfVmF7/ft/4uFiGXxeYIb9TVfmDOhfy750PDresh58p
Q78UlDqUeW401TLLUV5lVUcSVEs/7R449m57ZUfnWCrU4ClOjTY/tMJgsAR4loTKjdB1Z/9m2O5b
l/FTUnF1DtpvsNxkNXoBGtuFx1RW4WnLEtPyH8Z469hU+5RkgF8y9DzMAzaFpDfqSip3TgyvaB9G
pRRjgwfxN3//T0sadbyjR5Fck8g8/EDehwuBZfe+ZAhM7qVnuS2YprumLMZJBtMPPBNKS4SssPg3
6npJUabvNd6k2Bx2tKlfHvwhd8162kYxJ/cs9LVaJK0E47Ns459V/tk62Offl7poroJoFlfage1e
i5gsQscsC27Wl1csM006GUjzQ1xLv7Ph+DuzfJf9JTHJFXJjSC/XMKqxG87bDUbcVGsPIzbwEUBG
krUEt5G+BOZx4+elXJD+BFqAT99hzxHMQU2WIE3Zo4s6f6CufkNhr0Y/nmnSuWw6YZUKuUCttsze
yvNBRPA+4oBKHL13lLkwJs35dagkxuM9lN7vOIrGW1IaJAjttIl9PMAB/z6hA72JfDyjUNU5HOdz
d6W2FYxXLdCgq9NvlXv3aR5yLZD7M2T0TBrj0hklCTkD+rfHCLeUPiFR77d3r55Y8GHJPaGm4jSa
Y2rbJLCneki8remxShVnKEzuTkAMdMcR35jzs/BFoBm37OtPFD4IfKH+JHWqHL6cWdfUPPFG8Ina
Xm8kpkKUw64+2JAqFrsm/lWTlTQOLFP53LZM3BPle+TsCXIHBeFnjgVxfsitjEQUOGmCUGoJ0E5H
NaZXi3AiiuHfu5bN1JVtEfd1By6fUGLTKdzVomjBUxPfnTvk9E842CB2udWfowgZxJVwmjFGGtUK
uLhBT9lj/vvi0tGNC8EXRPySFoFn9/2sURu854LA2MWpJwfVGaES4n4XAYXirmS36MmxCiVJ0Mhs
UcZoMCRq2zAe1h+1Cpj5m4mM/80BU/khhtJVZyE8msk6mUN26Ny/6Ag4Ap2dNnURhV+B30fgtMqH
ULGQNjaJ7/+gkMS4o+svTHQf7eB8k3uYkYocUFUSOOHSQgzw2FG8FA8WKbmqeGqGf8RXgjbUr23v
XW3rj6xCxK0QXBFMPd9QROq38ygrNZEMIlyYZj1i1C5dbP8toU+3CNOnQTcZt6n+Kgqz9B5fq16T
Z/PjgUdzwWmrOHM7CJkCs/027bcQXqPdoxzfRdmYTvJlsI9pn4KeaCkwt3/6Tv/GQVhap8kf2/Jf
vJj/w1Ee1k0O0m0O6z9RQAbbLjtc30Uzmt6h9Ch12YFy1NrTz2owJMYh7/HzNsnx4NuPWXNwHXug
t/OxkB4CU9YafPcourteDIHCe+NBikLhdCSIlc29uuCU8WRScmrhTEyvVpk97iH1DkkildMge+bu
AK2K/LnB7k2cnuVszAlqQVM+xtytFA2aS2fH0SiCnI4nVHJp2S26qox/h6IQf2M/twOQW1edOvbi
3FM0vqCK/Dzd+8FxWOnlnjHhWJ/so2BA4rwxyZ0k1gSGZQvlofMnZo2HjOZl0Igg2GpoUMGyXDTu
/33VLARlLmZWkXUn+F0YzXMTwVThArGQj/fySQE6pcDU9d3IQjLExV+c95zAIC9SxMc7R1OCLJlJ
664ET/yWaLL868syJhvTPO0JYttFwHkyyakMDZJrKQ9r+McnqfEMFZ5ws/sqeUaYoSnJcWSD3g69
NO9sADnKS+XEan0c50GYaVb93YL+mRAAm3IPCJC92e6rLszoINnwoheZSEjTw1zVP5zd2kGIwfuX
23/V2Ybcch36eOnJoSP2YqjIW44vUWmky7CcrfVPXBYN5xPtnJic6l0P7QjxFhwLrWCwhdrreSHf
V1FPRoUaxVcgb2x79JI1aBioJFg9YmfQ7eKaOS7xy01V+9q31vxyNZ3k2DtQZNMgnlSW6GKsMHQw
TtX5HPzCaX/XkeLSe4lTm/CPvdqNaYaFEYhLho6q01EUNtD2R3zAy7ml19+EJmuUx1sJDdFowY8R
f6Woybj0ugTMciR1e/irECToScwfT5ejyZsOb1+bTMeb8OYS4uXKPMdaC7pAwyRnUXN/qGu6YhdT
rsSF8e/C1N+GyrAJgN4A1jnO8PnIA8QVf028z0YY1woiE10XzDPrGc7hSXYMdzbeeLfBdCAHm/Db
7NOF0NXFR6Zz54rmlGlsQkiVMgb7FUpncSXicpXcpbJzG6GIrQNTqHwANl2QWoVqEHFh2YPNHUGN
Jh7tN3O7aW4AxRee7m4dOq4yXTRgDprEeXE4FPos4Yc2Vp1kh3jLGV6cZs3HnJiWVbIbO9WR2ZRO
jDnDdZXdVs8dgyKJUz1ZAKR52pcyt2+++uPf5YEPAsRmfVRMZqQh00yEfqh3CfbalRzxQYA9wKOB
yGM2r35hpuaKysuu9yOCJtg4nnztzGkcCkL3JV3P6dspJgq4XFzW+IEMiAjQ1V7VADq4OD5/WD4q
tS/nuk3cfB1S+ZQEbJSt6LaDfOSxDEOutQoYwcrhxhHzIqR3zvMBKzIhf1mG0gMCE77qdLh7+SrR
i0uvxm+KverqyYrjvdB8vYy1bpUh4cwqHP2G+iEuI2gbQj1fFjN/dEaN1m9f6QunLeRxf7Th3UZH
deHRnjlXGC5dDo1Iu/R+3lCyZWiO/c48umCwgqZJVNaMC4ZRb11ZMYm75zF457Uj0uQMWdD7Zkx2
+GGcpitXC/Ajq9KS2q4NKlqr1BiE89eAwYdItgWqIUaa65OD42G4qg2YuPNNdrRwB9GigoXbZORB
DHpDIkHGMPOYDbM0jqbW0WytSzkTSmfp3RzXuAvEPhbcPenXlBMijRoKHVFdbjErlOh12NIY8vYn
PxDXSysDtDmC8HC4JapRXd248dU/jpDgvFlJTDVh3TuIklUXPBnPZbO0jhK8pYjMUScLiWqsAiGK
pMpwH7lEYMaTj5PU9g1+D7HQIK3yxFJTD23tOzDWWr9qnWUu7D2MrXXp0T3ZrqTSW/RMDKDqgntN
BePQEx5QeQCcbSSVJ+cR3MVDcF/CQYH4jOelui77P9VYgN6mCoYnsrokzO1Qc0RjLmPTZJ4VWcW9
zC2ZvHQmfCzUX4w+7KvdIuEmQx1C33HZAqRNQ/I42rxoq3ox67q6fi02IPrSNbxFCbIgldYNyke2
pX1kaGzGGBt6iaTvcI61ta2wfaout1NZu+fKidgGD+UmeUVK30Bpe8EwJh1VbV+aASdptoMBE0H4
QTbg+vrjf5Ela9DRGVQAxgrxGwBPTm+bchESBjiB/vPBAMcC/fFnBizJ1FYdMBGKZuBkvuFKmYx9
v9oFy976q22ue3xRkjkSVyl8jZOuaHHhMmcgJLnzPfByETNwCDr9+zl513y6BqDZeLkZiQLPFSj0
wLQRFT1tVbf4sv0dNbwiNjki1rkRsXhONJzRZ+zlgKZ50SO0vWdItJiDgQfL+vHbxDHbxf6XV/Na
aqdSafocfPxk8O7aHkQGxlMyV4m19FBUkph2Yussv8Zev8s1ZDf2Dky3DMn2M3c/pm//PUP6RbDF
fYIlmeT/3paQx9WoVbfbfhxdllxqLoEIVWqcrHDTtWicXjlblUhlXYecDPdc3XX3vXkOa7xjR1lU
IOXlBn+QnTu0x/pi9JRtZX6IxeXx5/SaUI18CYuQXt7A7twfXxrcGLB1SfVb2AtCUu0hcwZQLYaq
u3XuiFgmWGEgNbk9MCpLGGxn2r+A0lLCJLnw4PPSy0Yp+SrC87XBbNyEsLGVT5F68btiZ/rl7e8t
RbQ5THzwsbYZMaEOLDu32EnAhP47Ekb/E/CuMvqbaTV65IijWNwNm/2n6MmjQ1N2OZhApF5WqMYZ
oc6OnI6Qlstpkaadfi+72B1mRRKbWUMA8N/jXyPwinZf6SoJpfxXL/I06EwdLnWUi5d4X2w27IRo
pYgV56kLztHR+MSOesWhvYig8YopKfpmjbc1JsDi8UuaKOoOng/r3cAy7pAqAOjV5w7qsGinMTrf
Z0kexGUEuvVSTRmLg8tvGOw3Spf7JZiDTJpZO+QKsuN+Vr3DY0J6DOv2X91Vj9M3UMeVYRz58fIn
ME27I0O/Fd7zZK3rkQm+gxzCJuAt2NHSgO5KSot/SrRsclFZOXEfXjX2tLdYu7zWvN6RoDs5vKZ9
f8EjEgE19KBCv2cTg9xucukIGnBBNBPWfcUkW63fSEdvwlvyKS1ZceRz1ny+bPQ2g3Ts3yAIPEHW
YfTnzKmOjBvYKdk0Bhn4qmqIhflJ5nlg6QTOCVtYQDiOQHbjD6kUumzopVHkA4+qmfx70e+dNL+8
UDbUIMD/VJXU20fzQO8VdmCIui2hKIyDrR/X4zmEFBc7TjDswfA0r/gAMexiUmtcJVwftgIy5Vik
/Oey/exzLa9inGZc5g74psNyfR5p2erJettdV95VOFZQopUUBKFDhz3S5bAuJsxZITCt/b1Xt3cp
V4FP20fMMNthkcxKJPPz/koNOU2KySwLT91ykvbR5ysq1PGYvZUFsH7pZkCd+23UQvwglhjqErvz
NoSZACppF+buTFo2HtBtzf52Lw9sFJ/mEyyiKNfQZnWQ46q3RfRGcL7F56DwD84odmI1Q5RHxdVo
gCcNZKSbg/hUmOuCjOPdb7PE/VxMxo4AwQuwf+jVA0L1aPVHM33ESKJmkIItWYls8KJc9XfUk7+j
gWmxGzr298V4fDfPXsKkXMVnhWQdtRTtw5t1G8I2o1JtOb2HCQ3tFzDG+BX1vpztNNIsYgcwmSK2
sgAWx5v3BbmrXNM2Z4unCZK7SjWu9N3r/u+PY6TSDRnf4O1OrBc2Y/OL1B7/QRMFqz0zw9PCmjzd
PlKECdz1wWAsMa/DObdTfb0KSI3DtwrvLSsSblv4rwCFo4goTKUIbVbXi/mFKVGqkLkzb4TA/WVf
w2IhWw06Ibf1c6QV0WVYQzvU4c5GBbPvanOCwr8vIZy4xun34kuAcG+8lOQVIR02bUt3D76VAGiz
6r49NUJ4yULlpP6v4vOYiLX7Sjg0V+w5oCc6LdkukO6ZofhcILpqdwuvBgoziQekh+M2ydgQk6JH
d4g1EdgQcpXykrzhUxqdurvtX/8fX+2V/XmGCawqxiinhABmRTvNlYULn3ed7YzWSeMCivVnsmqW
M13uyLS6XQDtT74KS1VpOVyASzMZns3ULMt0ISdXvj1+K9UgPejOv1tudI885PIuivIBh2O7/7Ry
NnJ0ymIffzytjnZEOJJ3Kcld2Aita/PAr8dbH+jb7VxaRdz3cWuK9cyEolG2siCUr/8pBe5AtkDX
SEfqTF51KyqWP1Qje+oqyFPNbcAEmxhOyeiH5z1OdfUkOTf+O00nUcA1I690wWa3oLEgTecemQXX
ZdL8O3993WSeEaOr6ThIa9KNIfv0k2/SrLUxlVu00yqNzSDUBkr5UpFyt3ccEdBel6VE2sfy3ic6
mhGFu9uzHuTPL2csd6mgLqNBsh1niYijjQCdsCWXkkPNKGPePeHLyAw7jrIoCFohhRjjimcbR4KN
lCVU0pkR9yu6olfcddZBmpvlYQzQlTyWQV0e1x1Pfj59hZXkNusrSxCmnGr8U2cbzErD9HpSUSC2
0AkRSzgirpQ8pSHOwqz+PlBec5a6bO0JCgi/XnKIbQAmTcTgkchZKVbbzyDkdJkZ5abeESppj3uO
ZjZwJGx2JsAPEJnOKqlDN4UEIF1GZG4YMyiD7p5paLmqo/z54PsVMpNP6wxSpz+apflcJvaBSOlC
gNLLU+YVqo4GKrixh9ad5TVLWx4KYeKw7yLPwVB21kiSL25MsCYr/p9SPMqMJ/QH/iHv4xalEsMO
R/CS1axHtreQ9uMPj0GxnGszr/JrDlh6b8G/MMy/qi8nKbAI4coFCzvXgmXgrp8GslKoiDB0sCi7
HFqZCYmWDb4ZUUWiYe+5l97iWSEX8q3wB7qDJua7bATME4Yxxb/lFYf1vMqfweDcBWv08azlADqi
ZmJ3Se6XsN8NfwSYpoG+BhSzxakIe03unDwlA8sX4PYXoUUrzlAbLaNmCMY0vQdj4f7urFkqbhBz
b3Z7TsuyMxl1q34mCXikDK+hLoI6AIAw0/0i7xfu5q3wdxMaGA/DvloQB9l00xgUP6q4Sb4Td4Ie
fIYwEvQxVvzBufVACqbYJXgl5be+9j25GUTm0GK6T1ceUNCQ2AwZ68zCB3Vkp6TVONB1K9a+1/KR
fsFqUHDitUot1kyGQ+TZQNhKl+kOKzYEV6S1S5V/1Gtd8zLKuDnW8NY2pe1AKqDgnl0ardGjJDL+
BUgdD8ZIZ/SxHMABJjY6d7fxb8XZAgTYJCW4+J5Lx736gCudiqdSllhPv/kMSgWp681n8fFiuHR2
rlmw8llMROrt2UEb0ebZbQroK1epLWWNHm2mJa35eBq9VYlgGZpSpV3T9NXHNY0CF7yEV5jROT8T
zHnXrZF0lQjyV7Rk6x+kiUpdMp4fy/2LgVL4RTSmBFYR5JaugzzbOBQwAxa27QLny7y85cx/TXE5
70f0ygD/F5Xo/UWAXJFPjZxUNvVlD+YLXkhc0NWTzeei0yeTzCm2c8JeACHwbrhBlVGko2+UK11/
zyDq9rOpW+eKJ2C7OZnX8SB6HQKZTFV3cod3bLQR846zNhrduLTq8AwOBf4f622Gerr0omKyqNsx
RnUw8zNE46sCaVoHaZhNg5/0RZ/34UXFzm8co9yD4str9YXWbpMWj+yD3rxkh/4Z3qaPWVB7oFn2
04FKBVsSjboTApptguxw8GXAE2EWIUITvsFp9CIEm67TjHDApN3WE3FFUMQFeGBspuHy1w8e9EHr
+dkmKV/racVxn5Nenz66tdFb0VbsbNyvhy+lGtfLM3y0zvSA6P4m/uYX99kLgBedMibBUK8W36oI
KnNutoKmf7+Sh3ajBpJjQVojT2QN6/ia6D9VY8VIhxIjwZhKiRWrJVtDpScIOm2Xo08/DjwPqDos
9zlo2VP+7G57zAm5gsKFWHtEbZbBdKsuGtk+rPKRLFbRYC4752R3trTWYtaFseqM9pAZQSLWR51o
vW9kvf9xuiuM87DWAqYVPNb89HITeN478n+MjkseQsXjE/9xrI0j0JFzD5qpKI0v7uls+f2hq6X2
CvyWY5UMd6yIVuQLUsmV7o72FHghuk6YGNyHPjlAqJPnQXNnl//xQOG0VKPyL9sOoT93bJbA6gVK
XSIr2z1a5Zn8bTdExHiw0tIZlDOFtdYapWzYLDwgSyhh5Xd7YaVlAVF+xYho1J+F9mdSJ82lIG9k
UxQHLDPMKqZCokW0vqtbBFNWWKXoKU0q14FnBYRuq+7GofBHGp7+wAkvi6f2rvO/TReN3fBl9Mej
QVu7qC/FcSjPUlnGnhuju5qPsWV1h5m2aDgmNJXIzo1+RuQkckylBPVRDk3SrSJtTcOhvNni5xlq
/5n/0tNFc/fUPOHt2MG60zqddRgvU3TxqZgceEykpUxw0IX15sclhp5FXY9C4DlauVaE+fp2SA7z
+yJ3QMQWBaAoDlyzcmytjtEve5eD0U3NtdV6dt/pkfoLVXDMX0ElS+ZBz9RBXEhmyPsBTFPT4hng
TQhXkRqWfzgA2BD2tBgMavTuWrdRNd8kEC4I2yjPFB1DuH2auC7rRrbgau5XMImsrKuf/fDmOBIE
szTjDIciharadtxF1DUyAh7yUFsT2b+KoPGCNiQMeaJuWi3prF0yLg6UYk4OqcIhPtnS6NpIV71l
SxaXJLP+igMPOOSyo3RrNXvOfuAd4Smr03TuoIIVss+CUgdfqR1h3pQzmYBWC05M8qU/1M1cggn0
XgiGL4SgBeCo1dFmXBIxJrVJzYwFGYa+fBMd1qGxeXkaNy+ngA8enDLtTC8+spWr1TucwcPKu9ko
i7QHgVvB8X3qoxs2E4ugdHQ6F/+eNHBqy+gKtRCnXyXMHBVJWdwdYGbYzQhEjsm5/BF5fLIY2G4w
kTZN6B+0kYSrzZX5U+7AsTBJtj5X00DuXz3hJGtOxFYYC432QfMGydq4618P5YAfKDNGbo1y74RG
r/9qzR6f190ywzdftzC2Ikxx09k2YthmuTUliYPR7ZRA/qSjNAA2t0u/y6mfz5CxS1edhSDSEnB2
ZQI1sEgN/u0Qe0keoLuvANrm0proQ1oV3Qp3DyPsRJKYtgRHH479Yj1ji8iC/PTvRUygPr+wfGQn
z5hLPTVuZ5eaHP3nnKoGWNw0zvrykxXxh3N2dVp7ugCqJVyfmzQk+OBjeSpAZVhdQ5L8DekbSb1M
gOWHIxF5DnMJGHi+NSSQH1d5KbQ/sqifPR07ng4Sw9zNYveoZk0Ew156tWhdnhwbOLE/gi9a4WmH
qAI3jWuk7FjbdjgpG92GjxAko8JkkGEiD2QQW5JCyNQC2Z6Lf5Ih5+5wOKs/f4gpOHGunXtmiASo
XZ5h4naiuP0hhq4yGS/Vu0rMa4g79vXTnAZp0J3kIKhFqRqqrU2Yl7AAtZlLBJHw0IZ3pDk4PyMs
I825Jd2icPAJzYd/fqL0iY3lXhi/EB81fQRGQeNEILuyq1kHc4A3oN1i4AYTHlKS/KayqRzXeUo3
NIXZmRjduFi2z5RY3lHak6lEy8qBe/pbzj8uwXDq1ATZ7MhC2sCQZx9ZuX8fNxv7fPU3zysldrok
CxTEpQL1p7odW2EIHWL2Uvl5zrfRX4Ef2baRNoSxjh2qIn0iTJ6V3mVF+ksb+go4m/UygPVixc+N
Lku3gtumJPEL7hWcSDy5dnupZRHs2pikUtTZ2FTQjjwaO48ae3RTSeyRHYb5bngKLSCMU46pW55j
X1beJdAKrL+xMXQ2fATKskO7hCQIHlY2NjMirIBAszHVxB4qAplu/8LgyLVMg+NNNt3wQTHeCdrn
pOqMDUNGFYVXufExgSeB/xu7qL+o83+zvmkg6J/QEhtROGapW0uOwSSW0NtjO2uF5wPzHq1AQ6Z7
R/ZnTEigHxYXCMa0rGlAl4j+kTighjsp2D8p3EwtQxlNsOD5zKk9jDUhDjqVXOhAd55HIa4DIKBm
MlW1xFQzsVjTY+r1qq0CHnsWx1i7XsJUBbRLH690OvgAx9UN5TVPKIGRdb8YgP9OHTwoLQOEjawz
Hq4Hn79uXxvo01q6jBHiqnL6Ne2t4uJ92tUJzrR+qOxTdHbdfTb92gpZoPdtxOFnrd86rh06I8WU
kwAd3N+thzkyx7VcMZdihz/9LgmsFI6xeKjiRtzg0ytBDaoUP21SgxiP/YsyuUKR5tdhYh6laEZY
hu2yhXowsfcVxXRIVwmV5PCOfmb+E7ODVLi0p0EmSGUOKzhtPxo8UD4c71UxDt0fvYjkj5cjsLJJ
u1fT/NJE6IHnOnL5FZBQvpiqo5gMtFU0nYnfbFRm9kd3rYPZ3UBESou49wfV+i+IEiwa87AgqZLh
Py6L71vZC/d4L9Haq8hPfDFdnCgLCP3uJWBcjYzNUUWPiCT71m/bvkhI/cEM5xZqgiDD8Nuwd7/J
Wxh/4Ihb8+sB4+YkcM4okdfbW+1BPyj3ZjoF8jPnH+fsnBAFnEKEUxcWCZfB+VK7chcNR0Mg1RRL
RO25PjUQyYSHSwevafGh9f0/jFYBeIm2KYfEaS6Mfs7/4hiWxisVxsBObiAUUBSYpvN9fJ2y4KHv
rZrLBCkYrbtyzBd2FumT4JCkg1QqfmKQvOi2ArSBl83SRCPfSLJ6wsKs0Et7vg52N1UX5ll8L7ce
KnRgD2eB9CQieC+zvG7aSODBsQexofFtTWacd+KvI41PmYh3fzo+Uq0gmrVWSKHV7GPrRREG0AWb
l/Sz7zRugrsx01NfDT+17dkV7YIml2cG4+HqGmoTLe7ow2RJveo9wXEq1W3WvyDD4Urc/ElXIbF6
MoZaxHk6E1Ov5+w1jHDwVQhwEMAzHhtCr+RPKy1K+zPOlQ8yReBWrtWx250P3nVQrl/TXl3/pxQD
/YsXVa08vXwJYjW0p6FfIJEoOpQaWBDaSJoS3D+IEKpnTl70ppxfk2hN7AEvQS0OxT/f9q/Vl/PQ
eHPUWbv2nk91zdvNcwH7wF7t/A1DbPIgxjz+NoAn/zwjE1Ou25It3UBGdICIB8DeWzmBByHKLYj6
WGk8X9G5UdcPe2Tt8vshwsABRYUzPe2vyD1WK2P2vGUISZgInTqpA93oUHywbm/lROYbEGkVxr8M
vYOZ1iDnOz1JlbUFB4nr6cwQxlRBuQYpU69SW1LTj87ZsLoNOESX0l0vaN11dL95AnS1+a3oXr4n
x+AF8XGNk1EfUeJr9bRzJ7Nae1vfsYojTdqNo6rHGBiF5ob2JQPA+VBSnqo4V/I69it6JOHpm43Y
xak05P6y3YQEnshI/I38DtP7Lo/Rox4//OgYjQvaM/vpHK3vyYdhftcIJ4wUadPPgNhQ8S5ebDYZ
BVhznt2F8wuX7iIhNZnAtzLW73NUDH0IR8wtkr6pS90bAnTXLQdPmjHK7EOZ2fQ6RpmQC6+W2CyU
GqqbMhPB+707PjB7adUpKYpBMHnpofS99bPEz7BfBdnghoBmggyF9xIwxVPOIV4dBrm+3ySf2vSz
hxypiZlU8nyeoLw1rcyivi6YN2E3rqU+ANLgYziw4UrHEam7r6tafG8jltGEtuw0tmcnx79bp4UQ
pk/CrtdIDHXeMXLJkUfbX/E+drNIU/1/OD3eV2Ln3leA515Sn/974RoyINJz0tK7lxJpYBNHoDeN
rdKw/9KiJk8Cwb4s9P0of2sMld8xR7B1y8IOIZAymC+NMGyQ4kBHTZoYUowwT3zGIYUDV/h2x8mq
Rtrnu1IoqNcYPCD30S90cPNf+HbmecReF0YXsRhpS/a6Dtve0m9cIW+2P1PaM69DEfPeC7j/lM3g
ezgAwk/Gb+NaOHYwt1T3SrJfyiuBqLAaeuDBE/xVhgofbgG1PsrsOmQs/0bObEOSF4BdRh/tTEqQ
QiKmXtYBdXKrL/uYmS3hQioNflnebKRBlePneD5+dWaXvTQNwulDjhF8r0M/iublzqWWtORDTegM
0xpnuUQp8nj00u8kRLwEWgQ+ex6CkjBTurI706poAwhvWuRIM3Jj2HL6M+T/JQF+CGjBSzDI1dVf
5jMGGxIXOYuNPMyyuwrhWG/5x2B1PK02G/lxH5tR7uasSvf0BVFesynnfQI+fPpfgeA15qD2/17L
wS80R7USexovqm+WvRtkahaDVzsUx2gkRDULBbbKnzQNOmX22s4LpgvOJI1bug9IIw3Vb/e0KujG
TwOd62dsAGO27maa5/x5Vm5T/pTfnhPfUYwPeIVz1TL6adyCyz4bBX1s+ic7/c/fIhnieu4BgzHd
ubrvAk6eawOOILdaWkgi3hqWFwYx+dLJJU6yOWMl1ujgMymww1LxP2kBME2qr+tDsoF/U339evgF
YiSJBmZ7tP2YAhOkQKNrVT88NtixlAfSdLco88bZid+CtLTv7mrSH263T8UP8OVaHf9uJxqfA9xx
ZTD3UyVgko5pH1+LEVdwEr9uaULm37gSaaskgRPepTaiRaM7Un1rFXblaW8zts2lYyRmW2RzGBtQ
3SiQUUUhQpwyxpOBQ0QKgIQPEq/pLwQRZSc2ksRmcNlF+Xz3yO6RIc9Jp9BO01762PbbhT1OJMnT
h4LFM8/gn2RX/6KZsQ6yrRZkcpG+eSNLNti6l181EnHH1o6+BHoBX4WrZNT1CMWPPv2dcSJbSLh4
RlkXu4dihJcqYBgO8bLI+xHTq451+0mzoRBxtro8Fw5a6mp1m6hRyeyRWanWVxGSiM62tqTCIokE
AFKO+n2u9NdrpVqghxYqetUwxm5inMb9ySaQJPT7dIz6oK3oyIhafw7jkMCQnrbCN3ZtOt+5qJ2L
kK9LQTi0JYTZmj8yeKQTQKcgX+bCcuD70uZKstzeApy2xZvs7Wm9cBrRlWrgIJB/NPfli66OxZ4p
ZiTvamHcRkcDgjAHaTVs8js3FHni9OqcJUwkF4aWt2Bl5rC8cav7bSPz9SZnohifys2AE2YucIoi
yPWWA+6PXRdh5N/NaEYRfWS3PYsAuMOf4D+Y1Kpty1FUhLXlcoDOjDAoyWTYr+CBaktVUVeA5oBb
vluhWq5sAOfSctwhGh4mvNN5CqtpgK29dfrCul6NxNuN8f7xQX/0lu8RI63nmjh7HlOKPSRMRUfK
9Uz4GTOdJcLEqBHe06bB7IkaAQbkcIrtHXhRh8vbrY4ZN5q31iW4n74v0D8zJ9vPaV5GHnqyfAjw
YH8kovUVHYQhSuZQIRaKNkYyVcK++N9FfSPaTKcQzcj2ogmzfBY8ZFUrhPYQPs1mEaaAqVCrmRjp
ipzbrPwbPfjBBwhUwDYYW/2HKDsnYcTiYH2UwcmE9YgFU7V3xF6KenrFss/a6WyTVhQ+LLe6q5eP
LQkBhM5WXBn8LD/6Bz2B49KtY3GC/EWlEYAhOyvrOK+kNJUTtYeU2+vSAAjoUmaY8nHU5cQKuRXm
fRsw5XI2e7UuIw3moeBu2Urw+t2Q69BiWsPzQ9BPxROvf8vZ+URpQkKUznCPCe9hvQGA9uPVCfjT
7AWY3iRIRxtMgs6lpAnOPzZK/gxKe5fSBTZoZ380tkDJAzl5DfB9MEb56exE9ho7Rvh4r7h6ewFN
EtnK0p/Z26GI6YqQeyw0wMW3kJSwBxz386FHlf+CLzobhpUPGO2O2o7atxAIi9nQ2WCufEpn9r/N
59LO+ZARv+93+MixaXtZ2GDmiNfngfWfBGQrj0bLdqh4lddl3YIvzGRhpvaQdy87QCOURwR8FnCv
JOsk90wZLm1AtWrDWO39cBrPbVblGXe82yW8cPaej8AQJOZXmQWO0bO/0Uhqnwd7w24AWuzgfoD3
dqCtsVe3Vh/pxXyjPN9RXUMViNrUgerfAQ4/Wg+vk3LWBcso5LBQd5wkXCmc0jELEGNvsPcmkE9p
6PcIU8orUcJxY2E5990/vWRLO76RYdRC5YTXe565KkLRRfjecOIwCWaQIz85cKrrhUapc6IK4BaR
lnym86aVyWjfWo75Jv89Ja3BNhwB2LWI+FNJ43cBUAmWfaITmSf5oLqeG/fxEBRRWACiYa9/Dr6p
ebT3vjWw50UvVTTLnYWD98O2hUq9K4QaIa519l4Oa+4D/DAiUqzG5Wj5YZZlTEiqcMA3QiALsZht
OqmLdejI4ZK2ztW7sJJJNuU2pYsWaCJgD5shxQszZHke3VcDqtC2Ocj9eWQqY2JFRPL0RHHLI+Wv
VKDJL60XemRDgCPD2fh4cVQ4yL3JaNGomRf+DQ/f7swA4bmrw3J9I2AR6JJzKx2rc3dsG5+bzkOl
5nG7m8C3dV8HBUVWzqGu6TlFxKKxs69awZ45QipNHRt2ctFMgiJJCdtQF6IkUAy85X7rUu4NhBiu
nnR+6nKe40eAilHmh5BGWZa2wBFupyYOGpSGdpyRtMmMOFNqt1JIG0lFdpxh+EHF9MG3pyVrfM/I
JJNozl3eYpZH2Q3W4u+INeJqPnPHEMTH8Jc51sTAAK+ZEg1wwrdiktl6LNgcksBI0U/oSOmvAXtc
OUMOlw83sK09+s67pKfLone2Hg6HFZwI1kqHazvqhr/WVy2fVRCoC+XQIdYWoTxKlY5gx+71L72/
vlU3LB5GWEJjuqTXKmp60tT3khJ/CwT1ml5PKODlLUDgj4shZIyUq+3TE7kv2w96ect06VXOQaPd
zIzXD3c70NvkgMdcj7nrdadUm0hY41jVhyi72JZAluyVQA+MVdQUXQ88jxqLuDYUrOecqBY2vTLB
c3Y0ZlBZiUWhDxpcxJ//kdVNg4xH9x5A5XcPDHMSWXeliYPbc0vy9Wge5DS7EtUyN0bkPv7W/M2g
+89/usxaF6NfBmhjusYYs9G/hYKxmD7Usec0VFy/vjTuiW+dST+1nSkF24uNUSPgWZbcb0tB4eqO
vHyQRTrAcKrVlNhvo5wJ9j4PWacjA1zrAdr3FeO5AyUnxJcvZrVMlmcKi2gRkOcjQoSnjV93ljge
meY4XqsS3MJLtvko0cHMTBtzNk6jGaYO9P4rzyy6kvbAJSka85BLiqBG/iCW2pltXKU+gLSC4TZk
gQDbCEriAUkEgIroXAn28XuSQ6OUaEyd1ddcBIvz410thiaUxXWLDRa1pXmuajptLp2vHqcmOGin
6g5EtNZp7boU615aQwhx5CnxUMdjEaW9Vy/mT7gvzMyWIssSIniZbBXiNy0fV3BSMU88CJCc+BjK
0h56I2oFIhxRIH8PALYqpc8T5GAsTrgVTBHf4tbY4D8FA89N8JW1l10+0U9zRa7r9RkwZ6zcmuvP
LzkKTkNDJrer7vYTVgt4emi5WcVpwx/qmwxSLGrBykm6A8wzLnj/4D1saxdBiIHlarx8pdwuphm9
Cz8vV3yWQBvsbtT/uGWKPj7HNUAzyfZ6GPC25HyUmpFGtFWhbsq3pqeIuRobp9PYmCPqShZMl3Ku
VdFLhCdIDJvi0sWEqhv08oQwRmRYlpeCJJnAB4e3doMDDg9Rjs+CzKFGt1psoJ6PpDqULeF9Cmkx
YrdA+hJw9tR9xUv03dmVsQL6+ZGWxjnit3q7OmSBTw1EeYnkJgnPWGwMsChcBRK0zdokB5T7ChR/
fBNsiojCFHA/5l05kO6V7eI75o/MqK0MeqMugfMje2jcKYBusYzpMpPgfT+OtK/JgmqEAbV5lT3n
jF5YlKW96uX8HkdQkH1GCVWnvQJeNNalbomzFjgJ+fLzT4q4nRBD6f0moWx0kNYZ1rkRza84XZE3
fM+PrmcWEw8Y+IpmV1rd4psydMtAxOvsiRFhl6ipkz9NaevGq08zb2Yaas8apVWoiBJeFrCYJcYn
UW11/ReH+7BefjAtxdVfvKwDPwDXpTODUUeGQ083FEZDZXzWeasNiRf0i8WkE2G3fVPDbIRo1Nqw
eIOshSL9RCZBaXHMzYVjHDtcSdMqAOQYlV/pe0p5lJsTApaPKeFC0V08GkZ199iSbHmAyiCxcTP7
7OmAhVoL518GsXbO8kkCKrRK9CKipfv7yN7AkoiSUHVCn4DnsghsfZm8asO46hSf/U2VvjxlX9m1
PNwS5J90/vGnvxYlFlWB3S7n+hJ66xzgusfirT29RQPmyg0xwcyJJscSqf3WXmLMGfVBKu6QMnGa
Nx2k8AaSWfE3Plu+xTksz5LhoGzHv7ttgz47+yrf2LkAH4oPuUvsHuyRpnJbRMP6zuLps0pL3cfT
H4mB5dl26JWNQb9ctllx3NaiMhCLLtNLCUJRU66G5fLOkU+A1bc/qD3qZh/RwFToxdyzSz5QK4EG
AGWLYt4gclxoRYUlR5JjW2HoEXIjU62qqc9tn54+z1hCYU2LASfbwcwcv/I6klHxGoJraTv2pSLi
xi9YUriXn9y/IgSRj2lamK0PhYu5zwCUeRvYAdaqztj0lNZXDP4jIqGfJinRS1ELYUKlqb7/hIUv
z0O5lSHHG7CTYbVaZTklWh6R7e7wbeW9cls8eRiSd2hzELq6UjP8lvjRWXwCEmZhLNNaia6280CF
h0XD9M+4OOumYHHMBRF7OZiySpWOpQ4MH52QHE9/LpgIUzRwXPErIdKwtj9MfaqitAa0Fc6MYeDz
e+Q6fHuLjX6JXaz2RHapOzK/mFTGgWM7D5qFRHMqT6I9KPg1aBmVUJg4J1AsD4CApGizfREZjU8o
rbEF6RTU/HC+VwZGzJJA0apsRj0FVKzp570o2pdS+RBq9ZJrdGb2Dguk9y2aNTyfAQgywr6A9zA8
yFXuHfQsQF2BBBunTAowVM9eMVBiGpp5CgUMyFXy88bPZtFb2Spp/Ydfe9/qFSCX1kWSjLLTU6QY
PzUoUinvGi/9zEwkux9bSuPBnZ09XPfm5GrSXTLMLFnX73mdzhl1Oa/rDzUH12Tr+YeDWMeXYU47
AVjGIN4CpKPhEzHRzgWb7vPAXbgyjZ1rJyh9LnbEc53UYziwBJp4esA3UgzfyB0aa6OcFUgRnPyO
BsCV0nQY5ZDTqWysFCKf1SU8w3svdynIMK9/0XSW8VlQAXsmIB09kkSALcrofx9BCsKf2/J62WG2
+1MMrU/v9KuYhSauIRb0l64lC2db+C8bWr+0fY1ptp+RI3pCc7os8RzhA30nKC31NBMmiWTSEJp6
d+9Ltl9CaWkZwm6rUQWHrb9ZTtmowkSP9RaOMvEgCyEwUFKUb3Ql43BzrWHZDmeUui0NVzMnIq8Z
AgWNTOoWLZMmGmZnVAS0Au7NASOhahlRVt/35lV/KGRYbzbJ7n4KGxNH2dtod7jcKUG2wL7Yyx6/
ljfmoEM/VCNRA+yJtj57g9HaRYE799xFpel0mp97xvxIA+5ojckdLOUBOAqLhUT+/bJPQ6Fi+BCu
2LGoLuv6yj4CSf3WVaDlucsJqaLE3iwpO2COMDPsAIykOB+UpXkkx/nM8sKTCE6Gk/diVd+lsa0n
K+CZBfBdKpSrfZLOMstKYD/UO3R4u2P+0ntaCXsY7a0DmDAKGEJPxRWpIVThdwlxppMzjHQ28XrJ
1ZrURkk8tTXWlL/ayiww8ZZ07CQVgEqN/2OmwyPSx3HaMbndEiBN7Hu3+hs/SB69ISkTDciIuEuX
nAgtIwF+M0yKk+ojSYGPbNu1gwuJlCmoTHcd9GU+RrRhRsCx3ksNaONoZfGbBmUC101Grmdoi3Aj
ippxJkfbgufGH6q8OFTnANNSEDSXUUhR9ey32YvQcex+UfO+vyxOHK60QVMjtkemOvHmYq73By0R
XjjMav2o1ZVxwNFsH/RmuvsfckKwCB6+Iwa0xcrdjab/R1zYoDHvWRyIgXpSehNK5Eg0EIxcX68M
ar4oV9eDVQBeFZrlKzlo5ZpI5l/M3fdxtrVCIWhnwd1q6obgdkhTOvQJcBKT9Qu6ZBxi4YKnJ7I8
LfxIATMpE34A5GASRv88hm+VdTWYZYErfVL+ZDpwPvXm/Kfr5CG9AQ9h2Tj+Njie4HGCF+zXy7z1
dfi1CBM46YgCVERbU7ZRy/DgdIbH2YiIRZ3VPWyUevvlD4cRFZAYpK6O+BkXR2bKgp9RQe6wnOlA
6CWjRnohKOoffKYyN5j0xnJT4WmFiVgUcIJQ5BdfbjYas/Hj/yTATukt7zV1MqmmfuWZ3ejdRola
doMgQLlNaJgXc6NA2Uceswri7ANp4n5ll0DMNMqwmUBpPXH6AA+QdJh06XNUPGNW1jG8Bc88+4I3
NUH1qX246rzc7I8yN2YA/4+VQba6sxjkUDOr9Dd3qi2lQMyzFeN2uDeAwut/v17AvWZFRAp7d5Ng
ZPlxe2SBz25I7cODBFchrIWCTHY5vU6JD8suc6+Ro0lk8jQNUJbHsGTapCpbnjpDrpfGXwKDIqDp
/bcVYGSf7QbeXDrxkHhkXdW+yUoyxeQ7aea/pMxLcdLOAY0HaVad7XXyaLOhM9yMUoG5A0cSCK5n
6D/rbJ9uKxXXD+X2WBsqaGpSTEK1/+Ej5DFSbky6Ici8gSmdSfe3rPrp4LcQJkOdEAG4t6PeRLm9
/tvB616vhOFwVIYvVai1/qhNyn3gJKV8rIf4an1LcgbV28KzHFGZfiZ0qo3oyMft2JHtlfviyNvJ
m2Lq7Xhgj7sg8baWlH5guCmNutdm7Acano0YUSFKwVb4b39vw82Yuu1GQJFG4yVH4nkN4XIwO9pe
hFNRhwWWuzB7T8ybzHePF1DfKcaEBFqTnV+5qBsCc5q8sDomyiketUlmLWjiV+07HM7ATEFV/fE6
/n1ppZWEIULBbsulHIYtclq9/MyPIrhNi/0KLkHiCBA1u9KcUngulF8ImfCO0ITWOAGvAJmHOT1k
GXqg1jMZjDXKvkaXyK0030k/NBgfE/I4y6+KGLP/68UAgqRVMDPYDG7+Tx2n163bg9aNKniUFMgH
nTGpJfK88mT7QgLz72UEoeE6AANhMyZe637iuW4JMz25jPzpefzx6UPwgtUGMfFA1kaGJ1FC86vu
b/ee+h0cZMbjXKBDSqS2pTLEvKPfF4gbedKJv7u9MUoTFpV0RMJId9rSh7ZPYSMOkhPa7khZhNEG
rlU3hiE6WY+PHwHIhZ0xksXHfF2jhsCFmAIBImM/WyAVEbEHVdV5FIEA8LxlA4afHJN2Yw4yC14Z
UDFjYAp/mtKTd0EPFiOk9Wb6zDZGqFcRQtE9482gn00QxkVXbIYuZitIDV/k6k8EwJa3OPDkrLo3
VGJXIGgoxRakD0ahIRIj8wwCf/Rc554qJDparJd8z+L17q5E1zquaOS6/Ge+jKoIEU8i9w6iYTJT
FcdhI9JCFtpz8kvG083mWfRm3y3wM/072uss1XprSGzNAM+r/P1TcMUI9twVMimIPXn56SSIMloL
lW03yVce2xz41MZ+70/rPUMnsNnEga4feBrxhe4kMAhtASfZXk5ueVHF+s88B89FJvm/26oL5DFO
O2THEIi7JVf5h9DwhtNYrZTO/rUy4u1aUehL6GqXOQU6y0Lx3+R9CcYuF5DiBaMpll/gKNQRp5/M
9I8q2ykZ43A7bRbPEmZpN4ar2QOkeO7Vlo+7DHT1rg4Q1RrYnifaf/fIidGiH18HxcVe4Bc9jmbj
+f4U0lcLlN0Zwj3s5Op/Btkgo0VEXymGxWRP+UTGV/YvLhQ+K2B1CqzvrDCxZ5oOoggL8rZBSxZJ
3TqkQTVVt8WHJdB2dvcIIsV0FFGI/aJVev7/0Ubw+LabCTivhM1ynwaQlIp7hH6itE0OPfnOMQS5
m9UxX7LBSPFYyAtUW6fcDSHn4FQyCPwAEZgLqJsx+kqyt1gLQ9MNU8CKbuXotBIhGAG1bzoyUUXF
/BdukNG+L9eut3Ekn2azLkr2cQSj8naE5eKq5eGADaRJQXEpgRhY83hnjrXxPpX8BRqAIZetal7U
X5usJaZJY4y8r4L0bTtRrIqLxUuN8rz8zEtVUmDjV+fKeJRwrfaTBWsg7ChQ5O5a/HochV0uOgtR
1LcXI+UfRJc/zA4EdZ0azEeZegRFG53182gXANboBKiMUcOSYbKyzasWSUIJRje3JjWmB0PJrFOg
h+bBfml4aSq8CYxPOmI8e/fcnrlHNftHZH+f4R1+CeZA6Z4Ygqb7EMAttaI5+G2m701lPixLNFr6
rDH11Q8sUJufbIDOrCEqAEHbDoBFpeStM19QfR4LzCGHMQc+uYnjqV7fdH8D0Z1c01gbGoYtGWp7
ri6VSAN7OunxD34GEzptVJs/sbhlI5LxLgL4AsYB+h1gGrB5B0M04GiUToqbqagh7xuDlsupifZy
pZzjHKBuEZjLeDpxo6M8ZxBPKU1f91FjeOUME6Cekxc2Wr/TBAPT7F5zEVGpS71pYG09Jo5NfC76
h5pwINAxqYcO1hDghv6S6ba/dZP3P97eXH9JSpk4+gCVEsn96s8AP8oNRyKvCBNfrZuxzhiFJysO
E8V8YsjnowLfj/qBk6+fkQHiuZ0u2Vgm2tvwh2ncOcPLFF1kdeNWc+6y6PBOWo5AVzQNBhyinmCs
NQzGg6xC1yjoeJ0uLIXSELyMazazjc0bpLR2MTkXKBHbeJX2+tEnbO46R2z7VlNZbFtfy2/olmCY
m3TXE2+0kFFvBSClXmAh9bNArlyYw8Qb2wiiO6tR1Ih3iHMYBFVv2aZUrq2vdSaex97xMwqSGRRx
soQL06pZ+w/m7mqareZO2xIDIzmH4rpEp2If/hCpsxko8c4/zm4loyUAKwBDV0q/sxfiKB6qNZWL
RPA+5RBgaF6vQZ/1xKO+JPNBPYa9KIM10SrdQgUkefxfujW1G+4wFRhrZ9YYPhz4DTcB9oiOsIgy
JLMb8wOwXpURe+P5W7HV8d0L9QEJP7RDY3tEWJgiwGRR7IeHVXUZVnB4agHzI4utuvlvxX//w1jR
l1K+kf3mLFdOBCZvOF7ATwb3ZSCUx/TMJIc5rOg62HkK/UwmO4e9b/IDOD5+pzy/ZadIBQ5GcTcX
jqo0rJnfnsFFxCpYf/Sr74hso4zQnd7Q0duO7+cX1hjhm3G9VM1CypyIHZT1Tw0oD01KnBA85p59
97TjDfThcz1gGNpLVNVX4T0ZQ2pjiaGHcEvfxPvxvqOnm9jtDPcSBRLu1r67d2xMnyh0LtFJvzeH
sPjIwqSzxax1XI3dJc+vrmg48UJLRHeJcJCXpCcCuNvDEgmCt3As29hM2w43jlds0LlEo1/kvAS8
JyDudRN/si1dVe8grUTJKrwvBbTw3FhQgCSAs5sLmMwt/B1cyt2sQSpNhixq8JVzWQgQhDK11e0f
8DyDwRqSZVIhsky0YJms135PzgmMreORyVgsf6Z1oX3Vh0/xR6xagIr+cFRiNDQCjTB8PQ7XavLQ
IRNrU5U5gjR7C7IaS38o2AwjoP/aX4ianNsh7opmRCneDzw8AV0ZRIV0X61kbSlJsLJ7ZziCvhub
B8AkYHRvTAQLlHMj7FBasKN2HOf12DQKIKY4WrkEsHb1NuXZe6fIawzEKUtwONZVVEU0W7p043MX
HiEBKq56C/eueCrCrBmkvhh3CiBzmUDGJEEUE0GWAVcmNCeUY5HPio3IfpoDQfkF7wqNpn5EEUBu
qvaYX21WRy4SrK5FfSMw/U4rRPlL263DjagTkhvenSbMAkAQ/XOrRbgSSG5zoLUiE2GpqC86Ogvl
JQUKTOdb8WRiIXRzgF0o0gDJYEcPPr+Eukj7MNQzbijmc5IuR4R2kw7vLXvUd9/Hy1lCs8GTNJlf
DmIpgqOmpIeHMW12SgsUXLkyZBdLBV4dFLWQp3oC9NEjfBNHvuKCVNiz64XYwoemWTkFHbSwm4TH
fRtgrZ0kVAAsMNjOwdkaUMSEAGRFVB+t4PEvh6Cwhcuii5CXJ/GyCTiWDVbgJuVYTKMQ7RbMCP3v
Ft99B/XTP3sFq7cHB/GSRdIi8V5mN4tII5Bvdjl/EQr9qz8RyUmEbu1zfiCntjGtCcwA06LsAs88
2VNOLu8pviXI1NYlVyX0HvR8r87IhltV3O8aVb+CvNXOU/d3JVIqAVpvez9DBNTNovsXs/FWLuJd
27T/0adeGe4mMNjzkS4rpM/hwm8DbDVMKxdl9nx/Ubd+Hkz8Q666dQ+RUeSW1+ynyF0tqpL/s7dL
oezIJMr5yDDgsxxwB+B2QV0FntykaW4exhQTF/1wlEj1kd2ItO7xVbDJKvUAbGFuRj7tnGzGCBSI
ysqg0rm7vRYZnfUXlQqPpnOx3obXgClm3CoEKE8r37mxiuCqCdsZ+TOc0uNntLzsfPDJY/wPvIbm
jiTeaNVIfE7Va5sHtAt37uG7lhwu0axxc6r/ryQfaAiYi38HIXpMLLIC9cvwvmnDTzI9qQkRzBfu
wrL1SNX2+6jrEXG2v9XqjNQ4sBSRWgOGq+rM23Kzb4akZEqRypDDaWxk8pVxnseYs8Ea42nnc0sc
vcd14YnykDt/1jD6+Do//+VoxQv/bgT0sPkmW6s8/ytw1Tdi8SbvosbUJq/lAUijg78V+xnCpfF7
Tcr580tGwKfGsUE9+URYUmh7ZBkNQG8DD1zToYl6I7cH8Yz7lXaQiRo/l3wGwnbHh8irffwXU46R
5iTMxdnnL7M/kuglr9TTs2lTR54bgkBcWFsQ7VEvWK4VyJGzP7gxcst5sesdx2KvfFouDkhpkXUt
9iZmigcwfw3IQ0EQnUYX/Y8lzXm7r3kD4+eN9BTp+z9Cr2YN2EeqlV9h1OnIRdDFQuNKkXlvQ9P8
qqkSdY/ANC8wypQCrrAHWWRu6RPJrMsrhlyznZYt7n3txInKCYeCe97aB9xMR2pVCxF24nU3bnsk
TcQkavvgmyJ3rkJ+OccaiXT/C3gEZcgLlvzBh0vQ5RWnM6aIs82NGIa19G5CH6dBKzW9m2xD2HDp
lfP0XiQtDytNXzCW0EDVEV5cajJP4N0aecIIkUfcILZTlWmqpTCYio6eYIETBLsGP8ex1v+UqPH8
oC1k93C4NmGq0D57KtEbqOrd4Wh/lpJ8pkTxeaiI2F4ls4dElPb3UyeGra1EUkMtlf+EfSRAUuP+
jQ3rVE1JQRxeF12P/YYuGwIfTxqFdFcpSzoMKeNyRfrGc61YOgMnkoxc5uEnjrBPMzFQe2EdWE/h
pweZr3tY3KSWjms+vuCXniaHPtMGgfq3vf2aZ8E5QJVuIx63tvmmyNkpw15GWf+oidFUXnNUVjq4
9XmiEx7+wntbZjMR5rgX6kS4T9Kzn31S4V6iT6c4U9FKy48OsiNm1bizeSB6xmQr7gw+zaUfwJeD
/prZw2BhJxpqTqAOLwajgewO98slWStqI2Ijb/EFtHPxTeVkg/hGLIxi5ZxRbHMmV1HKGg/bJAmh
Z6P56ok73yKMzBFIaEe3k94NwVF91bxp2KySUfrNGGe7VA7Vfpru+3rYEGo7VlDUZHaoYNIZ0NAU
sCSf5BV86GfDW7LcfqMc9qPUXEyu0+FjD7KnFPDjh4lFLcnTgflJdJiRXuNjGDWmWQqlMMs1tZzw
LCgWDcz1x5szwjrgDZT4qPDnzuAPedW7cGYmV3ymsSdcwMEfRM4Dr59iKtzsK7lADCEYo37g7aIO
Wd7PsP7rAVZh+WT586ACaD9i0JLLvAuNNaOSxX/wIuGShDsBVq2X4S9GJKT0Ak1efYx36qYfyj2f
sQ4IO07oCAGK1fGvKsam8T4zD9kwPkF2+kGOOfPiQIK6Awvf1yZSFP/4xIB7Eo9AnF2eDDvo/lGQ
koi2BNP2nLpzSXy7eAFi4G7DElS0nMIgdB9sHGQy99KYYe8M4KnYaMemZZ4Xj8bFlB921SAElNxe
Rnw4cjTP8vA/K+4tiCDp++HLpW9Ioe6iKbSzMvgdLlGg3yE+MxmfjUZJEddAsVhaBPrDrI+WsPsT
brDE0lYVZz1fC/VkfbcF7dUdfFunAZNJ9p9w0StgPYeTMTWphUpWCgIh1Y/Paz7LSXcLzyHJlgwC
b9T4p8rrUYz/PkTy0bXm2mWtcMEwNMk+aTYRNfUxqSFSbNoiBWQxYAT55mnP5caVTYjDKwQt09Vy
JFiDnfVQv0jN2CmemnZKqt0kEcXr55HUvUccRpE7uZa12+6cOGAEiJWIK7KkCvS/a5GgqIDHtbvz
JaS7Mr6E44W4+ZcBP60qmVB4CDUzfg12C3fqUMBDLqj11Qg19RPK/waINCHFLtqpfCMLiU/UcFj5
n/XiHdLZUSC/Pt7Usz+H24zPxW7JN89B/94Gvn4uGd5UxsHF+RJF5G/y5PedcQwUup8gW0PP/OBc
zPum4a4un+uALnoaCE8q+ZMC5AGyxD7P3YxMWKMrYZ+EVP1HUL++EaLHBno+CehmAqAJCqGI/9Wl
JfoVtnudrk+GQzZUCQ2d+qnF6ttj27+TOvnwpTC5s1VXd0wrIcivXVfgwgc8tvS7XlEFWr9jygOi
XEoXDFZreasik/Y/mhoSMQ+M8/bm9LuSoL7jLjVgs7L2A87SVP6bPsQvg24hiYMAYFJOIqZH88aV
+ufyk6EIGc/l+NB5mmlI7eNqCOcFM0pfDoTbBnmJvNqdBwWY5B417ac8GhKr4RwNugRXj8CuGiOm
du0ASgWkm5XneMETf7PMGm5owS8SSBTDsOSje177GYYo2LI2mO6v/rVXjW9DMsxq2beWIEiXvAna
RK0v+tFyYv7eLFcN48Vi/yUZRWy4oEvtZUUBEurnOT15SnY1ptakN4MB6Pmz9v45V4Oi9AajJvnf
JkSrU4IS2lCWrs+eKejetjGw4O00cssewh/tbrXB4W29KsTBrQXdRZTr6APlXohZDM8ceT4ND5ms
t39XlM/0MUSfErYNXia5y3OcmKYVBWwYJcuBYvIkxaOjo5goxS3rK8I89EmRtJB6C7LdhOPs5vD8
jKunHiA8kC5vGKrF3ZYc+tRkrpv7CdmbUN6O9mE9joLNxEiVdAOF6iTloKzI6vKhn1dKVfIJyu2J
jfWjSL6j3aNO67TYf6I3rCgoUHe0GGopdhhO9S5W2/9cznvfv7NDDbMFE8/rMwqfD5FoAqx68IGi
WUfCFtKyY3ogXSS8htqQ/PBRI4v082MtozvkwUq0F+QsaeSjxfDe3wfod1rPVos+od0cfyzXAKCb
cy+qlFEic7DDCgY8qxXJdlyp/2D+STH49IXcuuu0JWONsj6lqoKJYxnVmJsJwP+K+/uprIN8yh0k
Lye898zGyfuDV5SqFXTcD649+3DYaOugnhVlmDURbObOmBy79D7L1WG9/WLjJEX3+JKOgcsP912I
9RRQHU7AxELvhpg7C+Yz/Pm7C2dJMeK9asMiTaU2qzbORQeN61tO2l3/YRcI1u82km5Rssj9yBk6
M7x9E490p2RWG22Qw1PRFZIMkwn3yY0cjsaNGYzNvpNrQt6OWBuXkGop5Wg/0agR7j7Xyv+P2nSN
z08kgo1TWUKWaK7BW4jQBBA+mfoF8lo6/siN2ZShDT6QF6DpFRnlFu2z/6by8Y/KDrei2kCwG7zS
nt0YUpBvQTSBCAYRLxNyZC4ogoATB7MPx8a8Vue1OseLMnVbrjKm24EFgrpZAegRKwf02/t9Pm2x
LczXBRY9RMRCa8Z6OCZuwKGWms1/F2l0zxOuhr+6V1NwOUvbBHuGcEozsxD9TJJzm93fXfgLKUza
ufGYrI48X7wXbNu7qVpXDTPYPrihwlDqR9jMfAsw/x70evS5hrtAlaxLDn304xtX/2QrD9NvUPiV
FNlNy6U/KK+4DOjNwFTVlLX4UL/557xxZzyUE8+IuQomADm8WjVWxttK5SbAkJHBjQ+CJPveDnpl
TJTOGQKb+1g1TwaLAYe6VvRpBGaMAZrXYajdLqk3xUaISSJb+cb6PDbTYVVmMAHT8SK1A9qt0ZUh
u5pXobf+yDNomoqUtznUmkvPBdw3AwQTqxG2V31kokAwDngPh+Hsn7DeiYvO67zdrvuQlz5bYLZp
m+9jFd5J+4KM4XEiRZd1bFdSCCp2JNd8Eam5n990Tu3ppUunzMdGItLlAwzigicER3sADEFoxuuZ
b8W8caFTWmAul2u+1itltLWF5zmu/VhVXu0pHxIoStMyfusDyvg6VREYmOSJeoV+RuYO++2mbfQ+
3X3J2Z5oK9iO5qir3Yoqueo4EAfb2Fxz2MDKu0ABlesKMqPEmjmKHaJ9NlFW5YzqJhojjVLsV82D
S7bWO//yv9CoZ/Fx5JD/X/n2zVXtzl5YBAkKv6TdTHRsS0vBzY67TWpvNr+N6QcEN56rK8DAtdKf
P3ADp5dpKlxQK9qBNhSw84Z7sgYtdlKoO8gfMKHsVw8jtE1oaCmg1iP9ZcRCNLZYFhEduL+pwxxy
ff2E22RuKin5ukgGM7pPeXir+w1kV2k5WTVQDa8JEPKV5mFdL4RVMmcGUUi4bZJLj2cGvN6z8LAp
KAne6kA5d05PqfCn+4/J3ud77hytkpkot1kc4Sbw3GnEAVhI/ULhlXyD6ecfCmfxjTI6pQjryj7g
rThjZBvvOgeC68pvtvhHzAph8mM9c7nCX6rdI9ZdgJLXiVEvFtsTKYC7KTVeYiMHgE65q3cT4Pj+
2dt2JusYmCnKMnmKXC2swoWIg3ZpLcP+kd5J1vBmIDOuQy2SdWFD8cPkCpmzW2UXTEqAl/wdY2MK
klzzo7Wa3YDoAb146jOfo/Y4OP6Tn40G4pe0gu1SpbUrASjJy29z5c7NspAb6SwXYE+z94/X3OFY
Mf1hsVXDTbLmGIxTYzsdQop4wGhJnCjQxc+MAOgZorvWLNluK0zyQlJSN8zrOeFhJ4ZKXCm/R/0d
P1xT2ECcEia5tEZQBKSJvc2Z4sOdaQe/lKCYXG1mXlukAo3RBjCIfHYmhGO2hA0sga9DyB9TsRmT
lv4iMc+EWVFR1buxU4F3PCFoQmKAqSfxs2ZFyOPa/+agYLmfQq72Wm5Jel35Q91wtjataC+oO4+h
Lfjms4RoBEqq/q+L7BVorZzIqDLNeGPZWT+yI0bgGE7e1LqkrzLG4UOnKTu/HP/j5opUXcbPgj2x
sWeeLp88IBBGFZCMHEUdhqyIIHxWasx7pyBbbxWPbrk2TCv2YdiSeeWf5KS2ujFDqAusVC2Wd7j/
a/s+v2LyOM2fkTtKnLdKvn5hpdaPD1O7x0MI/BlBV+VaiR2iFYaxMVIofpCOpvaPN7BAyBrX+owx
70lhTxWKdHun9e8w8MEEVI7lTVrl2HFeLelLAjP71Zzfmm8XT/L8NVTRP4Och3OOo/d7t9PZHwSL
VMs0wvxZj6slkyaHyASvQtpkQ7VnzNYOHuUP1PBHxga8YM4Btpq/fXu3k1XFa7fuDH4aa60SA+y2
pgQOXywnDHUzadbMz9kPMHrmzYZXOpVeXZ0Wsajp8iNaMqFLwj/tqZhvLyl91RnCRU2FPIHT15s8
QagTpYEKsyAjZRUAfkqRsnCHVjm16NMUwJJyLqcsL8xFB810AD4wB2Kp4U4aI87CIvvjsatUl720
FW4KV0M5g6lC6KHNyu0W0Vw6WKI0gw8FoWxytJkxhP9AWrk5d9WMEiKxlDq1c9d8YLcPEBXSQ7kI
biOpc3mWYlP7ckYtT5Wu09cIXhByigktLBWox05w6wYwXKk21LBGwmujZa/1ETjyaD+M1VZXv6ps
1wD7ZhvBIdbI5ONSiP1llO0SbrNyzRwczjiExUC/2bujas3+oCU6/miurFLvcym921ueX8zPHm8f
IS8L7pIGW9YSnGY9PTu36hMXkmX/DIdh1ktFYytxYnk8PgmF7jWXrq5fxeD6P6x/3Z+bxCdV1CV/
M58LxVhDeC9OaTj9DJQ36FaLZzL9mOFWvi0C7+yLcpkn3MvAVYpMfyuaSGXOm9i9CFoSzcEJ6bV6
WqfqPSda7+gnGylbp+L9sZP5fSwX48aH1WUN/aseag3NTKeETElJVv6391g4y4ZCo6ek0HoFLMtb
LssxXtllcoq9cTUPVjaOdxzK9QG1QbDAz8zUajWRWAhzMbnmS1cFMQr/WyLjlWZhw++yX9uUllnv
wql4+Cz992s8EZkrkL3BwUNPTcI6lzy8xpSs7pic8OdndiQVZISbGDTmDT92hXjoGZ9oTIaprz83
gTL50mUbm8JRpS8JYqOUOZnwNHJJMKND2XmtexAEXoT9ttAqHqTHM5ZIpqPF35cAChrtcuzXK4FM
GGjB5lsWV/cpl9VufBKjs5nAQAn7gGBdye7pI9QFEh81v6IBx0EzWeZZaIIYmwjgSfjb2VlQul1z
w9ZlnE3bimsgJHYJluaQzYmgEbunLlRYloQCNy9EqeqGYxb4RjGF3FcL8/p5VwIAtPzkvymzjgs9
SQypOVjg9jjR17C4X5hC3uM15MqF197EHTYqBjThj1pz1CApVtlWJZ01q+qPB4xEXtPxZNikkKsl
jw5HZL62PRHeVWMOPK4zbpoETFeSGx8go/3U/mQaMIEuTzymjQlRpTw28yvG70VrKSR3fXvYNpl9
/8C41VwtqtzqUIGde9Tmbv4LQ6K1Xm+DAi/Qqdhxo+XaXNFvuzzOezdfpeoPJsIww/CrFkrFH3tc
TxY4F59UfUMLFFuStaZDE+wFLqfWuV21I++k6BVOf1Rj7Cs4YHyWX8PWo2vvZNx6H492ea9aVBTi
m96DTaHy8HvIHdHhjD0hSx9y1X6P/YGc5/CZ+CqTYEJCXCi8tUto453IzQHJtA0+dAHbjl3woc2Y
1rp8OecI27wCuniaaWOEUnco3TW9nTaGBC4t/LD5lekFhREELeTXQUQkKBpSBfn4kgMaTN7d6Uh0
872Fit7VZegrlnsxCO8GISRrb/5EaeVlJk/uJQ/610PIi4/91sjCBKft11Z1kJ9qlgR340AVjhV+
Z3A6n7Lxo67kqDmZLZe3n5EoOrEKd/slIGlMFoYBGcL6FOgJH1S4fXWSL1JDwp/2GOPxr4Tl8/Am
HbOooAIwGCirFwWRQpAA4D2HxSns8wwOpzAbtYMV0EQnVyN75pA2e0Fh1euKx9oKB41pLdF8ZrS9
+vbvw6Xnva2poI1nkEZ9cgtSZDK81Bjt9DhSoxW5cpi1XIikLTA12UbeIo3EhBIOqQJyoSmF5ET2
ubuorQPtbVH/7a4VlEFtPqdJIYQGPVndIlSQaB5Cmqj9Mt+G/XzvDU3BqzcXbF9xEB1f9xzlBS61
NTjpOeaqWTQwIlDiQKdPMeE/bLpR4BHtVYKNm2dxYOo2YsJLrlDgp8xo9v84PqRlpga3DW8sF4Rp
CHjfW1kany2gnzC+wTGqplzr/OHE86sLFzD5w0NfM8d6dc29ZeN20BAo19l9RknXf8BEdDmC0Hr/
4aGe8c6draQaKjSkUFv+5wrQaGlLpIgKBcS9ggbIYb3kh1NCpvaJsLjyDiz9VQi5sfPMjB+tU3vt
ghtspUJi7IapCGXERAGFcchVBbDqc46qO+xVXzWIgfaO8DbpUw3pqX6zRtse91f4GiMghveJFhvi
YSTVq9Irni23MaWK9BXL5NlMRF8cRsddSFl9wlOUAAWRPc83sMfhHaO47WwlARCzBN/dcBH8cmiX
oo1YdQRJdz+lIBIHHipDBUmEocKHGdl+4Zk538idCDOys82233ZjMfMdug/FuVFpuFdXvNyQsS0S
IjC97u/so3qc2IyloQU+rK8w9VZHVMap1ScdKF8LwtPmeC88faQxlk/9T3BOZc0FtpLiXNQ1ownE
Za05SxbAfQydbR9LXguDgeM03dR5H5Bx+E16rPUaP1iMHf14OxN0WTTO9AAmMZ2u36EirS4KwtJ0
jcHROeOEw0jEDKIQyIM9d1MEJi27UsVMS8SUxEK/7YGVbVoHDBZ7h2yBJdkR4nUgSomp8KB0wSQC
qJo5EqaTMdm2eMXq2RasTRXLxDP5IhUDETfJqnBsSGPGtlyCn1HMqoyJTHFXOokaKC8DFNdEKbwb
gPacf0oMOfxrmpJ7vm/xJHNsngANN49PYEmkCQzq/iRrfau/LVBtrfQKcK4ndPzyTKToQ7poj0sO
pwtaEwXWj198HXjaTZyaSBbARlw5zn0hqeQlbAM5gdkwwoL40LlCQHz9H1jyatdFt2Yv5gLWIW3w
5tXzl+9YUi9DGLOl4d3BMMeMm33OJOCNcRGoTpSiIBbNRYxRM3WRjH2Bwt5irHTyKraQjstlghnf
sVaEpMsBEu4J53SWe5e5U1NBMDmmfzNxQHrlAwyV+9i1ycWkQ3+hak+hZP3efzsg0aM2MV8OL+7Y
+T1ZLUYzyDW2AbJHu7UmcBSVff+nsAMxAtH6XTUZCdUEyThnWhkPSIiKHwdw7Zl48gVlT3b+1ZKX
71FjgQ5X0agC9Bzsy/NRQmmANdVh9Dc3kxqYpws5TP2nOHuqFJTdElO9Lt8HWoKa+PLQL95oZsyQ
bieUva41zHpQDv+NMWRCvybvU8onHtrlMaU185ySGkrLoOMd4uituqYcZ4N8KGQpLqMb5lAN86l4
nvm7+I8MeQqrHUhHn45tE6Qq3SCREb/z12aQDPUw4/AmGA6l5wCjDF4hJmmnfzPbbRP8u/v4Rlnl
NncJFS1YuclrX7BmbLYqzjpunx1IOIZ26oUfqd81kp/gCEKS+exYBew3PWLOoRYuzAjzd90KbTJ7
fve+cEdZfYmjwVeqqU3dduDJ66ZNw9uMvbnJk+luNRHx02Vvvdd9SoyHX58HJ4rxpV4NEX3FiPz+
wvx7yfGbHNo0ErEIBMr1E8ZEUQB1VXX4Ax3fctQbtPwAUdd1u/wdPM4P+NgzPOMuK7MVLY1veLSE
knZ9Kb51NQN/aNGkRiwwHZ+SsaRjt0ix6CALewg7Kz3ffRAetNoeQPTmY8OCqACbAk5B46AOFsFv
FJ9yyg4B9OdoMUAE9KgpBx3iTljh1xu+2RajhywtTGJnLj/GffNHKUwAbkCiT51GsC2dtK6JYMA1
veLeJrJKISrteRpS33N+NoDdqil8GcFRqEqCc1zS5JXGeSTGn969lPXzeXyB8TC8+4VhIRLnkIQu
M7PSuXgmdJccDeT402yBP0srZlngmlvHLJBYxmWAXA2iOVR4rOjRAPi7koVtnnq0sg/jPvbse7HO
cB3njGK8alve7UAjvT5CDSMabQJFYGqIOgUrd55t8i3HDMdrs3lAyIdKkTHWlUR4WOcpThwrAAUU
W1AyPeIGPkzSgHg7ziXsR7qx3GdWGhbIWXXksG1g5IuwGLQFDpDTSbTykpzyK9WBXfFZ6BkfGNbf
0LdeFbTQWkI+9q3xTyIlCb0TYl/fJPAptYjuKWP+8HjApkhqU1saSu7tPcKhKhTmr7cULlWpAw6z
YkWUIYFpAlGjDg4wrqD6u9rTIIvn77R49TacCbJFlT40Fce3xIDsVaCBdxLqMwlF0BKDs3a+zNdV
gCjNT1F9ihgZluNF9LTSxtwVvUlur6V2Do84mgxT/dA0s2Qt26oCnPZt06/jFj/lDxbkVpPHd4xZ
5LrX9MW9sUS6yz4C7jsuEQ4jUxi5oE4HNlRVry0SaAsA3k994Qpsj6ksMaBfRR4f7/E51Y3tLdgH
1oG7dquaKNmmote6sfY9p2wdx7PjKqGlP4Tf/2shTR1CQsgT3ZbbT4wT/SphNUTcoNcysGkSLRE3
wq4hKxFmvNria6Du2zx8uryCWm1Ym9eICVithIXZM0C2OLplTK9Ggdu+qRvYSkBZolqo8ZXCIer4
BrWyrT+wkXDPPbdg52tRDVifM0b+IEcMmZxvtzOqWkUHGtqTwaVKykpzdcBSmAPKfZQa+ZoznLQH
r8woeJkOPfTUf0nchnCg+u34l2ALWP50qtUEOBOKmNF0xqGo4b2gC9j/7n5JBKecc6EChH8WpCFR
wROXgBk/wsq+xAUCwzuTS6BvGkfGNxCciWu5Q9fL/kpvIwjZHVjQJiC/xj/wJfC1BDDEFTrPnzqP
Rtz/g9I5VqUdBvJtBGunN4YVrv48lhjAHzLv3bIFfBwoHaOwdXxCo51o63PtkUfdFjzmrnzzZilH
cHmI2b0lK6WOEAbzlNOsM3XE7lLSFUBPgMj0H7wzgK6nn78b6VWDNSygxKjSJw+zjUpKvShFfV5d
eZtHUBhDX1q1106WBbx4/Z7waZrNAIywxxCsjioq70KKUTnTw2ZiQimum32TZO8VPV9Ad4fi91V9
2wGkLAd4R66sWavMobTti+HPmnS+tBVZoaKZeuzhmfY5cHM6E++4xSpMX21AfQ3Uz7qbPi8DcWim
OWuJhtowV9VDcrhAZ7mvoBbKtjS/KL6eGZ8rIVZp5lYfN4TzCDochJ5cyRy4tIXwMXXWhUX220Lt
3Vb3ht6ycZxrwFZLYBXWWCYVJJ+FRO/sUcu8xULs/rD4mytauUsHffXRJuMxHyDcAzh7N7/EIFMA
K6Bdqr8v4imlclhJowaFgFHGSCgyyt1Q768KLpGqZypN6JQF7Pphj+o2UUiYXt1zsVxPxGkktOEv
njKQB03w7tMBwfxjEd+3ACkLp1zDDJBp7vDu6YrY63NLR+UebsJnUdCb556bQ8arjOaZElAj2E7g
R3l0yf/h6EkQSl7m54I8C+gMZzhKSbKZzuQLCe4TjvUBE9/Qj6WjVJqnTOWToGMPfZKzOBSaSLp+
t26l5X4AhBgbc2Qv2pbRlKz2P+r53fRnPEq4aStcp+qUiikInX6ePJfVkfra6fDv6qsHhu7fJDp7
YYo4dNbG+2UBxuvSJ182XluK3sRkqGNMmv8HUjxm93j8U1Cw9ERR057IuRpdoZbUrEGOd4gCoVHo
hWXSASDPYntKOhPHZOjDYdeNsM4wsfioMu+Jvy6WrJ6InqWv8997MHl+CE9XGC6hp9+KqgRB2xIE
MN/Pfl0JrWMxe5JWSfwkx0o1W6XWjXBrGehi+uMUBINNfRlFFjnD4qA4VemYFLGwsPIh690S/oIJ
D0fsqc6bwkt79iFGVDcYe+3LTt6gCXvBeSXsoTGl3mrcLAbyvwXbElJCdIGvndOoeHsflk10+Eo2
UQrOqstVgUfEo2mZjdC4uHu4BeTEovHh6nrRPOR/dWiuuZETcqs4BwDTKUvTU6iMNyMHf4N4MYkb
a2JPltGU2US+sOuvWz9H+OxOVOSNEwmnBW+i/czG2Kho3lPuJeUpQvg+p/BlkKhd5E0c8bCPGtHD
j6FRSOQEg2dw2cA3wuxt85ZpAYsZzOoRf7uJJhpSy0ulE497nGsTl/U01fBx8eyS2NPGNlcKwpXu
DV7Q+a/Re9P47qjTHmOTQv/7F18s6uYM2eT5PPirflPP2lLteYQlFWDmoBBFgfrpkElcfsyQ5plo
7WKw5kk5Y0kpH2Vkp9EnefaGM8vY7yQ6j8i4iVxiv8OULQIY7Z3NewCDJ0JtSORrvXjJ2mjQuAYI
aOhbbhIyMM+25aUnJTCZcO7T8Ioe+9qx4G+hdODLULn3z1ASlcEk/+aStFKYhXdEhPz6LVUVyv5/
glofleJIzAjL1QOBfBG1yxcMzQJ8WqEiPXp++ZwZSi+to5mSgPPKObkiQ5J9z3PzcZn8lwMjRmLP
Owz8V/lIrCcgbDdiVd2IbwEYHsAowxJTzq4yxWFYM6OzUaeRRdU+xfKz60NELyGRV2uqNSb8Vx5d
b9dmFpqkQ+mJLuH0B6tO/alEWygVHRWJH9vOio2S94GmZQ9A5CUDHdTLy8ahYebpWIxw/+wlXly7
mZLQ2eoEesSR/zShIt1U62hXKVKsJq2SZu4JPtyesffRVpcsSXiH0T1YRFr2reVqkLL8eaR/bD+8
0Ds71MebDFvlRFl0QTsFnByZV6eIVUy3fmbVWRXD7ql4yUzKsuwOSDS7PxenJzUhv4PJSi0YwuLG
+/3cKxnR5GTl+yFTpEyS/ifHHj8ZOubWtEbxa2PycffbmWixldk54K0rWDjU9XayaByLbHzZ+2Yz
urVu4+79DnW/CZw6XiRLqfBH30Gi4P4E26ooZEMt2gf6m5tVHMyc/wRHDkd+093AJ/PEw8Ekjcvj
y2HT+YSeINvnp8r7BRbs11ualt5Q8IgShYsQOTJn02oufEVlJkAC8x5m3Iz0guhaMCVYLr9rrnD0
IdVukkauA4X/7x0QVX/yjbuAgUlgMo2Szvose4yj2yCvFy6jyRahrYEXSc8zgAh17x9cVS8nh+nT
p7+NIG3laFGTw3fck41kytvemcHxPMwru5W9Rvg3hGLWOBliKYSFB+lINKHr3OBSy2udlsEqdnqX
l+11M2+HKUZW3eivSDpB1/PuuDaY0WqoZdAdBkOzGme1uhtNO4uXQIScK02RoxAIfhRGu5Qff+Pp
0iHedFUu4Lo1+DpZPqNEqt6R95kDJndgJeC5Gph8f6BIGsfO4zHz482tGtNQQR44TE9yAChFtWnb
cex15EaF8Ow+5ymzlfg8hxULW75JHu5bKkPDtCzV1yGiZbA8v5tOnSE1bzQEs1L6XBFOmJfFq8mp
zEeQO+Xs5+RuAvoHuXzupitWyubRzBKeN9ssaKk75NYzlgX+BeiJ5ldLsfKUiV4l8h7Fdvgm+63c
kW/2hO5uAblsuWcxLrdp3fNoKiOksTxZKW77mq35nms8GHZ17Jm0bGUwk4w00MKbISjhj2XL5lHU
8rgXqt57uD0YpYGbXVNBqFO0MATya5BO7XUAthz5p1OAQ5jbAyssyu8EBETvap5Bi1eca4BrTixz
upjv8Sp6r+GMfTUA5y9kiyTCN4VP3h1C61zbiYG8demtGUMhRYWiqKN3cJWKxwzK3hACrx/8s9b0
/4hM+Vm2QWUlowKNpy0tiYx7MTfEWf3Ic1AdcB5aSA317BmN/CoDnaAZYm4xo243m9BFNZ6nFlaU
3FaSy4xdhRPM6mhp5oFplI9X+4t8GALWJKTlxuEo1OZAuaLUYPL+TTbQEYFavrZxCem2o2c7shB5
EunpZx7XLmK0WEXHDoxvc64pa/jpC8eIezs0jACxEmGgzPSZnfWOyvjxJD3ftoCh2Mh6BLnkYrHM
pM0Cn4o42wTMls9YUM2oto0NrqxRQsBuUwCmkyBDcFvDxO158JJ36TnY/01JpHQ3MVSBddjFLFzU
ihcQg668LPuaOojBjo7Ujg4L50pTa/MIbB4NdGR78Vl9glXyNfrvovhThWF0XKemEGDZdbwtHjsl
68qfKWvLggOFyilGYt9Be+ucX1UTKM/CuiNC7fGN4yVz27SokXTxOUQsddA8EyZpw9Uzd/kAX4wU
y+0lx8biT6XN8R7+pGjBHc3jk/lYs5WQ1/uw/veRNwtfloL57TlElMp9cwbDmfalrxul0V00qk9D
wQ+oRWv7ESSHfXwQaiN0jTvswvXICvehRmt5cqUubx3BrBnbRlMVovY9H3MA611B1d0bJc3WoIa0
oDAoSwMwv+gvLbEbfEdgw8FfQEMnFr9WCbgTzIc/ZxaY6ejQKWN4K8iSH7kfxuwTQ14iGlKfPC4R
I+SgE4RkXg1VeHtcFHD5MqKccgflt07KjkrCGt8MqmDeDY/1om6YgX4ig6KzM2gBuGYcnmaa78Nz
PAD2c4l9HJYWiKatDEDwdh/9udBywDPowjr1vh5X5kSnuIO/1tZp5WVFWbMCMN57zZX2lJGPWqTA
uMQQoRtCNV/nD8HwzzAFDFoudc/orcKhFNQZpy0i6FOy7ocRM5D3HQfkcHRF8waqZ4bsia3fTuET
hL7uSiwNv/tFhNj2VtM03P8d9iZBRXeyIlKWbqXA/G/9gONdJW6Z4tEym7iNwFbje/KHhRtNlyob
hmBtcXwCJGeiEakxUsihah2ty9R+ejo24H7QVzmZ1bAt3MLLRFc71BRbPLMjTkfuuo0Vtjos5ixg
MxVOQ84lazooh5GwH9HzX8KHIIOuMpFTzUhgdJoUYX4XqUn8pYJ4dxaEiofV2bresbi/XUmmaHRB
e8n2E+bjCtScDuNOgXheG77SJ+iQ7/xms9RgWIPbuT4sPzcXEf5J4+QK62cjdlcMQJIYl+kzcpyZ
fJKykJPOphEsYZVk4hoos83qWCI5nnvGT8P76wHWC5VOpCUgCBCfbL6ZPKbjs7c95MnAkuB7Gfot
cCheT14Hl35paR9bo+bCXDo+Rk2Lo/znaPFjj2eaqqX0hKJiDdtEucJiJVNfIx9/D4KSgKFl4Ftn
RJbvxOQRy5nSxDu5TFXnu7z5zlDGX60Itn7hzG5OpejXIuhDejcJocullHn8IFDD+MwsGhP7uyta
mcg8vbMAD5ZF3s1ZTJuicJfY+XZo8rXk3n0ABDN4cdyx9+hvxfv54e3C9MlnEXNkdqj1NqavASIC
0rYmZhoB3UH1bZGcXd1pC7KuMVSTPUw+yIwo/aKNJnXqnyKMDqNmbtlkRLh44udNMaezgPlqCE7U
1QHME7rrHYb/9jIEoOCFUPjk0nzlH/6/oD+V4JX58YG3tjt+9HFAnluaJbkrWsSKQCNFw8CPUBZ7
DOevYSpTsS3ctKjmr2ZxK+r2b/kAJ4cJxQm0DxZxjivq+YR3F5bmSmAX4LuiKbqisZxGfTgTwmtp
ZzU5m/WJqouln7F9RcWvEzmLFGb0DVchu1NAYku6mUgJnb38YeEzkas9JAgwUoas98d1wINB2SXj
lApN08ITkrvnUuNEZqsA8xOZtgiaVO7hwHfMkde82VhNqcfkk2QRUkemwndXjCpivhu56g0Z39TL
lVT3JriaTT8MG42aOwOwVEqRcZ2ZSCaX1voy5wzhLa44LbCtvxovn1g8dinmlz1wTAX96FBigTvf
9Ry/1AGHj/hHKVhbaqmFDqGXJpJbSDL/Pw8vbwWBFtxk5Kub5RrBXxi43tPMjc8W9JPhDehRgCMd
IX/6UmY98liz+kQ0HsSK4JtPWL7qDJkQP56+d30J4x/vijuE9RHJM6AAvpBHzCUfAvtFQekb7Ibk
MrHlsumJgk76ku0VPFCiTO3+sFsifBY07oz2uXCgbPzLnj2C5xFsrhVaW1Bk1ZFMEdOeAPDY8HhE
AaxssZlYQPTB6yF2sh6jf30J4kWGCOIbeFzqSutdmwwCi+kaERhSPyARrcF6sK3zNsNyS+xTnzC3
eI6vxPNsr26M3pwQU2epmmEB68HG1xGZDrF3wsnfzXaSC83k/qRbKmrpIshAIN3uLQL2u2PO/wS2
gOQnlG8P/OZWbWvE8iqTgBH79kM2Zg9etiOiaqQH4S8PTovX/vBCduCHvVqla+vtcy+NOQnoRGPQ
OwidZZNAVxvADaZ0XxhQ8ibvFQ/zmDxnr1F+kztQ0m4BkrcSo32IBsmnxNcy4xRls+1tn+g80s76
VsGhhSv8pgkVjIOovt48F88i/Ci3PGfjqJQVatftVJBoWPf+JQ4/xTN2gxh21iIxZJk0AxTGzeDd
vu5omLPsdqQ8FXsBMYYiPQL4AXPh6VFHeiwq9zwmg+mgpQnobVxY8lqqBhGtFH11UpRCg4JiVZxn
Czvdji3dSOg5hDo6v7yQJYSKEd0SbIDvTTFyn9qHmhuzhSqtR5J4fMbw7YsHWVErzuZoQccq6VlF
6pz24iw2b6kiI4mXyQycq/j/SQcv72+JZyVdqh1UkcTXHh3O4tSQEayVpyXbgW4parHj22mK8Bwc
gOCxEF/BrwX8fGDbJ4j5s7tgFtW2Bp1yJZs09XmjNcLgzUXWRtgL2BIPxA8uQESunWT8Mf6S/p1a
b2thzdmaa5C+XFDCe7XH3PcGQyPqKqWHB6pp7+Vy22BW3gi8qWH3E6v/iO7AEm9BS+ke8igKAcg+
D5oKe/oRlJVMOO5PFOWymdSmd3Z9BIL4vC144DtabS8X8v3keMI0C/+/1h6lzB05XjqdWggULfjr
1tqj38300FUSm5X0MblHeNIZE/JGO7tBiP7SEvdGcUYsmBs39nqORwwJ8QuPyDhuU9WGUm84zRMl
By0ytRPOgIjm1DThZAUXTxKCO4jRjasjP2PqpyVJ7OAerGuaoD6kYo+B1uNmrJSaLB4gAkN4iP1O
GX5FKdvkSj3iBu2sjc8HxktpDtC7kIZsaA1fLeI5ijolpv37a/rJd3/HE8wOv92Mp73rBLx4tV3s
X1fI1cLaPvF9rOzx1VcsQWcR8NPFSnfTJ9W0heKoQHni3P/edjAQEx6SIYYtI2vwvkab9pM+O8KI
ReElSScpf3Y/vhmmohQ6UI9x9dyV7lib91QFhWuvN05o5UjjsC+eAVWBv4IAykGAyGKsAKAQvWVS
YjCSn72N/6SAohL20FUD/oOme043EddW5Jh1zwcOisGUrZL1LgFw5/WOvtCD5iEAZy5n3+yR4+Y4
+ctDiYiMXb4bLad+4DLO4yH4ZIHX9e7vPbQNK2rkEXuu/EZB1GTp0skk460I6psbVeGVBkpgOfhJ
0PQ8Ifq1/tCgZKp6xhHRypnd1BfzVlHUO7XLFQ9RV/6A1PFMi7SmMVvFZwPBP8OUkC68eP22aTzY
GnJjkSSGINXBwlVswmPin8qnaOah/bXuYdNd5cfETL/5wko3KpXBDyuk9mHrYFe5mPNGk91oQ+4l
cZVsgPvkz73zw1WAmPDWUP5hUt4QpKWT1XPqPydRTGgOPYfRoa1GQNfUo/0kgw0nfmxpm7PzcnDP
14e+TRvIeb2RHAkkmfrm21ic4fV3BBJsXJN19qkEgIrIU4S4SrmRrU0EU76zf9DLBTIP47fHIMqz
H36Q+0QYL4h9bB8EiNcP9sJbOfwjBTcK55YwxH4rV3krOz5jhYzkOkurs+TgTpDnOrXsFELU/1sF
ozGVc8mOgyaZR8zNB/wVPIRN1XcMr1/ydPJizo5iGmjOMLT7Jj9KDMYZEBcdXkOvkd4Jrq3/RWHn
R2xE+PjaQ461Y+EszBPEbnHzi4cuQqNCFH7degwaeP1gGDdaS2EyfZjg1EqVgzTK822gJy+99IdF
7o1LDLfEgxwmFF8vzpbjR0YVqGQmgF7SC893mFlHTf8XZeKhU5iPsLVKNxX9tcZzfIKrKgF1iEew
VTfhbhUcDCuRhc2EZd0hDBIlkp8yqnwV/EWbTrS6Ohx7D/rCTGKy/F69iAn4NBrwG8ltY/Zqdg4R
R3US4BPMSgB6xNpEPqYdVDj08M3G/PCkVK75gPrtLMtSUZzTqcQVgkOOGbS2LlfXeP5PgFtzTwKc
84+7gNjBM2fJHSAtIm7EgrUpW4VehK7e7ECURkPYVds0m8wivdx1LDNnl4PCIkINZ3hUWBdzkVlY
eTKeLvDzuMhnwqWukH2Mn+MTEBBqJID70qkJAFZS7jPbwkV2ZwWkV6cihmp72kcv4bblVT1quHvS
rKi8Cnua4fxV8VmMfvl7eIo91fu5K6vsNcuWdy9R38eBnr9kpujvWAYnxpuUesXEVagSvMyhQE8X
1n5ilCzFZVTrB5lQHW+T2UfvKIDqCT3uXUSvhUt6vxvQlS3c5RbmzDjXnHRrejJWakNwOHE0EI1i
/h7w6p3VTd2WhDsGN2HDNoKNxghd/CMdDqA6LKCFcM8O0LzCrjxNYTvSG2iwPtw5fb7KPCjzX2vC
63iega1JOfm0WgWlsNar/lozukfNwh36QB8v3UceM+EBws57MCLLc+v76/nJjt+WoiW9h9ZA+895
2lceFUVSBMtaUITeJKo0hwRULTLmZxQtsiNn+9RdL3Nm2PdOj/RZy92rx3R6SJLjFEdNoPGUszRu
AyXmhnfCaejJj5OS/npLdnNPF5UFVUvAVX5fmjDIc5uuQDLnRJi50clpV48/Bwl1p4kSv/H/VhkD
IjnXE5UqrCD8L4fiO68FYQ41cODHWMiHH2hAsh7RMmkp0j0etVlDv8ni44kpvrQm3Br7cnCVpMI5
GGcfTQCC7yMGs453Z6wUO4z8IWGr4UMjt5BK7NPhx1NFkXeV7NfGeKj7kKBavt6rqRVJIIK9A5ph
212QyAPO8NjkLyAk73RwicUIbe3J8Pz6T586PpcD+7rEQBnDb+Hay+/Z92qdHbKX32CW3K6r/d0d
Hg3652LSJpYLn6ThMTHMiSdr9uCVJWiI0/CvBwZhqK+WXfCIbKvRwOZ77lrZH1rzZyT3xX/LGAMS
K2gJbXNw7JNASDl/zmprR5onvPcxm9JYnBLInJrUQkiP3zmehhLCTO84Wg3x2hCFIX59sZWCtK9T
6NzqMtI3ArlRx44xSdbTwgEykUcI3NzvbfF4IQQWVOaZUer+q4Gx50+Kp99UPwLcUZj8HYml+Qa/
xTdnZyKtBLIkNQZf54+iJ1nJIWM+RVPOtmlk5F0r1wO4i3fK7u/9lMDe9T3IxHHuGxOzj4t183hz
aEg4tF7u7CiqNX6H220cxIWy5dTw95/04AjgAO89lZosvSNU+UD/I66KDiCC4EGpvHOhmS0FF3yM
YMgtXvwFpMz3bZ8lpwg6pg6zwrbDqMBdylJySCePLmkGoE3PQn5+Z2JrtnPAQnylK2ZLFUFVnOOX
7CjYGCZmjv6kKsN4/d9jP0OrJ0dsTMQRmTtHqNwsm+SFfyuy50oTSKBecvX3vwOrpLK9cxh8jCM2
QYvkVGEXzcPqMixektwAJNEQ5zOyHfpc1Zc9YcTQ4jMdJnRbg0TycfB+cy08ptDJflfO4NYBYhAF
6cFz7b+jeeUgyb9ogTdaGJ1EX+irmfHZ3Jc+IFc3+lzGwwsfYRNEOcnqmKqH8g0OvTUhkUCS5r2g
kBgnWckia0G6pXXaYuyNUTRPihmOKHbnkdZ30/hMBDyQXd52IoZ2EmdrIR+sQgBv0ZbXU1mHfVvM
27DylYuI54Ow3tDd9sNn7MGe1oP5z0QtQxu5N9p7JOMrgIzvwYZ4WmqM+mpixguhA61xJpFwLDq6
dcxWP3QYcCWRZLIQdbafgusjuLYYnguoDjnCOf/3B9P/tPZ9DE2fQT/jculxkTVURLP6a6H+02Q8
fQg4KU7XvERIMLwFkXRUNDvfNT2Sgaa6AnMmZ9L66TmJxLnCejzK/g2MUaCrYC2G8jf4tXEndrzx
Q01O9/6V9pkUvBXDhGjwvWPgwuQiTSosGXyXHlJRGNTfY5xEqIgDLEYTybphzvP6FIU7UjpgbcBo
Xb+Y3qwUz9wKVjJm8CH+nk/71GquwuFx/9ROYfVgQCrAEc5PZTmD7NTvWFs8zL4Thv1hWK9kf3HN
kHz/zlmIhbsIwG3WOUvFkhavp+rMp/0FB/CsFG3Td606yxRN2cLTFn2Gcl6ciAeNwjPVNxTVUksc
AmrUQLGKRG+AMGO4FYt66ZrnEXJethqAjzh/Mkq4TBjP0n7YIn/Xj19Jcyqi2R6fVfbhKhFPn/HN
DFMQahyyaEgfZJIAXqjL3q2acxeVeZr1WlODa7I9YiGEKwmzxL3iOxfZlJ5DKotQ86Dh2yBbx8OT
i+JCYD4rtvKkSrtjyb16uYP9cnYt68CjvLQT4mQ39xnfqD7VIQyTwLG1KUEfqLlYOPr98UoiXpvD
ZtF2DnrIDvmMC5vafOmwGHtECXe2ouI/XxYo7n5jhA5Cb133pdz9lJPovg9RL0RP01SUs90YOAS4
0IkO1YUq1152qTdXWEH0xqa96F6gc32crURUWzhuBqPFxQDzlAmLACYjDGRjLSkjUec/eE5DPN2V
lro3hjQwaPaEr595YdyjqQ9hGXrdmZwSk1t1t/OQpwinN04aF2ejZWeJfCVyZxQDEKohXlIU9TAi
rj/YvHk6ek41aTN2Icj0zX04zD7mDOhrHJsarXh06TwxkalebeKX21zh8C34fh7zGpxMVBeBfTQO
4id4FimsZBqe/qL+PxF0p1CzYA3w/WIB486t6bdb6opzdEd2UASu86WcO6LujnzB5HG4JNWV7zud
XHTLueI+hcc0cJgfBU3T1IWksSAweIInnuaBS5SRgcns3q/0ZFFltMtgB4iOYw/v9v0zF1v9QKG+
zBiPTCyu6veWTwxpJHZynFN1p5C+T1m8enYL+T7yowMVvbhCGsY50QnYhr32yIoJOlya2zz5/lm7
bAx4FlHGJKGzgHUHPuNlJVQLkv4H3EWgG9Gm0v2UKYL+THMlW3009qYs2IOQJki4XbTIEWbGKtcn
O1PjAdwruJLyGdsa7eb6bl5mQSF/Lly4Lpn1wBV+KisNCsTVFcqafJDbL8NT7axLkF43nx6dxoWK
hruvnSOYfRSnVFsSrQ+2+PnD0cmO2S54Uov44Ap/msqagJ9vn82k9HCP0LaUGN0QptnonC+vx7fZ
KTWShV2E4YGXVxdQ+dyOAXMLEDXFO/JCEgOCI6NT37iXZSU5wvEW/HFm5Xg8+xJ7QiQuC4nldR1v
8OcUip+c++1LncuutcvGcRawufqArhXHixocQwtC/SuU2vSuU0PAK3tgPLGlEROIukPuK9eeIgEa
Qs6hchxq0wB3Pw0LyaLhwI605k6nE2aRYUmrnC8NfJqVPiyDd8bMG335Q0h1f02otNshf1VYzkS8
R3mx0sDcY9rrxrFwNJ2174tQyOO6SPud+dStMK/4HFAwlorZ4b3jUW41uodlp/K3L7CcTf5OuIWR
8yCrgCCZ3JYUE5TvmQ36lVCTXDSDw7605hErQ+bETQZmzGvOeo0mAF7UWcAtgxa+Vn0TmAgfifm0
UEpmouNbC+5R4tTmOP6db8wITApxkCNyP+36mauUcMHcjsyjaBGWEht2l+sOuXB2tUg3t6QE1/SF
jyfubxJh9Ua0i05Ejyneo/d+HcohYhLlSPwgsjH+QFQjT3ZXPoz3AYssYIk91654b7HJV6+Lm7ly
JjxlnyqhI7SGP8IqSRUa9+3zucD1PzQ/WYUc2lEfHDUkIFzW4UT9UIASOz37zkyzzEEJeK5xD1dt
4qRbRHwBHndBIfPeRXfH7i0pMGbQr7ym3QME3r2WE9qTkz3qnLWpqH7USWLlLyeOqDeMyY1hceXM
K1BkMSZbPvX6Yl4aWQJGJIdVBvl3i6laEl+eca4xYzbXsNApPRc+sngAz4MZL46SuRmPFU2bdAMn
0xj1VFGis+A1fFFS3cxNNaDtN+vWtVeQnTWEygRymHMKgbqUjlnfJlzZYFalb9D3pEPBgzWDRsQp
qT/OwXuAeVFav6dc8hQQ0EiVo2txxLatMbXhjEEIoSjzc4Uu/CWue0yTBkA/aQQPxIAjHsMABxdS
EOw2v+A9C2ftIq+fuOW2mD2F0RLYZf5zyXs1WTOHMuNJv9h2zRS9DDAMq0U6PaPPU0RSp1DSFwPn
w/evPHdiZwYjV8+W/fpSbQOMJGts/5o7vVugWNw/Z2j3bAUFc/jV4K73VWMHe06xYsgfGIeU+n7a
wgAHY5WsGI1BaImkUaiGak5uATD6wt05NNuJ1tDAcDnfXOqj8xEpoH0onyjGE+PxZc5QkbZ9/m3T
yWrua6ocFO3BNOqWAFtPQ/30jmRtRXwr8rPoCb58Gz3hUdVBJahGPJl8QXunRzXC58XBI0gYLAPD
uaesZYsjSNrjkdf0B7AISesCDUzKrH9q9tGkvDnulNtrp17FvrfoQCmp/v37bmliSxv23R/C/wZ3
ExPwlrz/0aGoZu4iNPtVQmqD/qqvgK6OQjKQOAKUhPm2z9PCsv03Es7Y6tZDgLc5O+Je3j/1TZrU
Fd+RroA7hxV9zeiEy2ZAyq25p6KzrtYLijKOMS5XD3EJc+SDkXAiinRv4RWTX9ajzVHcM9Bf/ctO
slb0LVGyQc+cAr0FQdCKWzv2OXT5gAaOFc6PMz5PAOjpOmiTRQPCyBd3HH0ZQt8K5Sg49kyxNUQ0
wBLyAzghh2pMqwGloUIZcrW1A8OUdqa3z7PxlXUn+CB9DTI2x+5inS2T+IicBpgLQySC7sNV6UuI
v38IyKSmEPgZzWn6vkZ/ODPR9sDqgPNt3DqKnbxiDnjEATwtNbp/RcZrSYlgujsE6EqQjekvmZ78
wwjt5VjVOZztzIrteMinULPk025MMQ73xEMAYZTx8X0j0282grLVyYYHRO/Ik0nG0HMIl8kHS8lZ
1gZHLTB58YaNqxUg1C/GoOcGCA7vLhUYML23FKeWX7xM0eMNiTZ3aTIyFETaRqsyVs2WfcRcwEVA
a14z23ziOPCoPWzA37T1x31RHkfsVLm5TGVWpHtvFF+y46ejJBzpTt5K5WvBvAeh8uPyUWqQkgeT
gHOnw7T6UxTGgmD72uB/2kpEc0gLt9FPKpqL+CaQP/naXlM8H1gTWzHRJ2F4IqGMnH9kioOWGTjf
ibAwBZWrhbdrPcPVtV8vikIAlP63VYn+g3hCqOT9GLmuAGTXOuC0RyyM67rz39AGaDTMiPY6ZU0e
uVOG61W63CN2/VS0wXg+qOP7BvRXOO7s9vF2x9e3fBZBUbDi6fba7MjBrPJ4enUwQUotPde3+92r
8+Y09QmGnIne5AkbpAFWETF5VovOYD7LtsL+EDGB4CO/oJTIsmnhnuSpSx8TJvvhqQm4NFbxPMSD
EM9obkUk884H8DUtxS9kP/GkaZ+VhXiL4gjoRi/BzYxaKvVICZRRFY1oXhf6JJmJtdgswslCn47Y
pE1Yc7XL2xIIp9Tkx0vgRlueJbFbUJIhFdWbL0uWBLdL7cJsG2hDLupyk8Jj813BqnpPw2/aTY7A
ZxLYf47MbWBKtMuiS0aoMbaFec7vSH2oK7/c4u+nO0mgNs4/KFJQxy9qwuZFnGGKi5DD2Ph4LLqa
BOLK8iEMwxgm4p7WucbL76kAoqE4DCQKMAKq2TAwW2iuKKrgUyKbvEdpFHBa/VOvboYRF9A+YNL7
agEucLJUvA3bISEeLUSQWNh9l5ddt2gtqUUS/8REXHQKXB2CrqFQTU01gmaHhizvY5yQNdxYaFDx
11Gc5T4KDcBS8PAEdAR4sJ0ZWsKINE5DPbGVmnKTXepspF4Ae1gOX48XtB6v1cxK+RPYeDehjp8p
l6qTywAPsphwfOkJXKFGYbpLF8VMd/RNNb9rN3t90ATRABH0yoJgzIibeSdJP6ajx6RwzLSze11h
ANnB3kPsXujZbd1SlCm9xh5QXweFCOKCSXyudheesro8/asHelhlP7ARp2tTNoGuGMshNxd5z4E1
4qKHDzvsSX32G76lqJLw0xYRcqujYJlQiczmkipQg+AEIpvdC087rfnD560X+vYnqK3hL9EavBRY
rlAHvXwQviW7N+O3jz7g0U55oaqkA+EzXoTPjtU6OWg2exCnVhvGds3IoFhsKUPtQ7x+qVYhszSO
WkhVdVoJBMTxEsvD1OoMT0N6XUoIXxtPDPLOVh5MdHQEZBqqPX2K11AQH8nWLQLQ07K88TTT/DVv
7j1n+bJlh9mR8H4WmdrjzTqjXvDUMT3snX5R7vr1JCuUWvYgAbwtqDVfs+sz4bvIjLy418MVHT1B
z4PK+Yug4h8KXyofOiw1qleYhQzXFvuj7hJ6YIzY1wHsnFFaTuuqJvvCeaZY1QCFVYf6Xn0oMwg4
I/5uSCyPtHlYDC3s6hopgSTBkWWw/p+FlSCi/cRqHgLs7qZXWKhnXEjchi2eq1WvVsQQn59+sZ5y
HpDWA03RfJntwiGQ7EELkbhfmHdbbQo2sJtlwwy0vDsGk8DweJg75KswHIItYLVMNO/mgvrhUaiH
bNjSZnkEfU+Hnch2ipJnBXoPpVXkHqLziuarKfqh8MxqYcEocEov6JVvrohpIupXt1aLYX3FE1hV
dBc2WCRbTZIerf3tAq8bVUzos6ghCCXcX1WsTN/bfce3glDoYw4JKc6P33kb4OAQXaBisC8+gdVy
dxxDWHPT1Di1OTgm2MnMUCB0yKM75Mwb9GnYxOChPnBB9TJLl1mcBq5BABeulKpGwKLYdIgaBTEx
m1zupTl3eAQEymq09XJYyVgZWwZPMcFKFIPFN3sbfuvx25izn8sDuxP25wqK98/u+7CKVfwVqKkN
A51M1KFSOlSyvoXAxsYqISEzJ+0sYNuMF+ipSbi2Kx5HO0g8OnKgQwftUWHcuS4Yqdi6/L5YyiIN
Ta51hg0lsuaTVnonMrpO+emi2hPh17alAV4wI/Yarv01hIT29/pPVkoi0Lp5fwNoyZ/GvfGmfN3y
3mBD+0eUy4SPweR/LIIekR77V9AvlSibefcreFNcpYLZZRPoa7syZldOYfnDrDruqKFnOdO9lgV0
5hqBu3QOh5l7F4K+100aOJBISUxrh170jBotpfUlDgpsoeYuJmTOrTCtQVunxiJnym5HXhBY8JEz
+zAuule6B/mTkfEkenqQv/LpS/kAwpSDFc6hOaqgt3zIWSzlJZH/L+vwVJ9NZ1EjKOkOmFi1Jmpu
XhUYxWZ3/UbTCbPdSNcGX3hFD4XpFsR+F0HyLhEhsTgQkqv2mml3eFSadspRD+9YaUf1326320bN
U83+7QZFBGHFrpLSaMfub8OEwq3C+eX6B1R0yA6op6yDUmLXaZrB2M6weAhygs+sGhzaxJodOVn1
qkB2nA01Q4/4CIiQuTI1xR3XK4102Nntrt7S0cudRjLNY+4WSqVcIH567j0gRRMZmhPWV1zkpvsB
qM9zsES/nNRP+3k7XC8gWr0wSPz25aiNcBKOwM9neM5tdnKuj1t1u9VJq56tSg0Af93CNUKArC6o
eZ4909yx3dZdpLdsT/ss48EZqcQpexiJz0HfGAZF4dhERZxgS3ELs1u7uOToTi0c8wwcaxur9zR1
jgO2/gsmL9dXTDmbe1Wstvxg51z7+kw47Jm6OvTxDk6z4p28USff/2KErbEncxXbPeyQa6BVFVx4
h8z4JPlYwPBPef62Z1qEomCFHtHkivYdZVTqPVHu4nOA+LYDmuwx8zfateovEQZDTvnRodnSnv0Z
IzlS2dRlv4ycLMetJYFP3Wcd0nD7EtynpdNNkflqA/0Ie7VdFq5KtsSBTNNSZtEpCu6BsBfWgIj4
kZMtDyS7v8OUkg8+X//i5NOKepvmQetBR1pKo2JeVTszOhklvxClsDoQFhOlx5hEeRuc/zMxiSpw
hUry/LozEsHLAua1RbhivkrYfq7s/a+OLHefbfy7osOG5L7HjVCAjI7yBDElDGRyJUUbPLNGWvhE
Z3JNkv3FkoNnd36VJ4kyGLRQxs4ibqB+FlxW4E258zvRgIRVsQ+D35VdD7aQ8dfLUANLHAEZrdXu
7Lye4CSJBebpZ1rC999bHWriPf2gur1McNA351cyicB5rs2OsPDzucdyzqZlPN/9tI3nbmVVBsSE
bn3lWZTdX2SjnXojuQY2efnfkCUDtsfYtgvNFmLonmMcbyHgyCsBUrRe2Le8K7H/KuLcgFqm/y8n
C/4Fnv2VR/1zfHk9dkpp4cyP/5hrEo25ysuJekT7kGQnMv1Ljbj5ZXpdFw7VJEg1Ct/Iel5Ib6jk
eaAkC/HgsBjGBAelJ0mLqR56i+YWfznR/S/5OjzNO43nCGNUoczrwnmVi64emPg24cqvnvyTgvyq
a1esg8Nody1i0BTcWI39iF6lLQS2w/ykTInsd+GQEJfkcxQ0vHO7G0sQGWtxhzm34MRwdBzPkdwC
MZbvn+o10lSMVdkGxGaXJbTp32cRFp1fu8ewNGOMnGHHAC47DF1IMgTJex7buh0LD4kHMoKZJOss
YgEngYI+KDjAozLq+vBDfhnJxFJa/Lbuts2Y/rwAJzKoq6jUIiCCYXZoyjG9IwTgsnV0HNBualZC
01UAAIJ9zyac/wf+zyGM1kDW/PUwWyY15Fe/nfNSlJsADvbBH1BKiul+WLsAct4hG58izi+hia4J
H/Une1YAisbASeuMwZ429WnVi79JzGm903FQoCedzc/fymICt29U3tM8t4xl4x/D3EBN4ewIPpBY
ck6JIr3JC2gPsAPOEVBU3oLmOB/VC01TtOrK2PTsLog361b7q+kzG1bpYvCYQ7mon+unbWjzYln3
UlD8KzKSAKdkv7nLB+EVQPtfMyE6aSWPYaJ0vPGWT6ala9jf6Kt8iRQUQ5HCjl4jh57TmNKiE+cG
2QUdaSJQzgh81IqPoRsZGm76W+UrkAgTegBWM6I2YAv5WgXFQKfs3Gbv8+YvvzO5xNFm4o8eOsZn
L+dDgtCtwg+IeEpyq91j5Dm84cLC5xvmGSWrOPiL8E7y2Hczg4i3w7+s7TUp2HK9bAt10rOhFWBC
7rgdT4tGfpjaGCg5sJg4KE71vlBBpupjWsC+YQ/X8UEDJilvxPUUcJlUGFeuBRf/XdqiCxLSHRto
gwUFYvFahujA2NzhnUYlwXmw95W/HnqzWv0aD4ETU3mkV6Jg4XKVGmbGgDub+b0MBFAltvuspTL1
aqH6wnKC7nnwaUFVva3vhFLERvs9cmJq5n0ld2rqdt24wqmlHDcxPi+DWvQUdY2xUXxRLbbOG+9u
jphV8c/jk0Y7QcMFIpmJHBOHqXvm1xxoovro/vzqt9asv5rQfSZxCmFz4VXd9gPZ0Fa6u+P5fk57
/bkjaaw6E7vLQyZHw/yZl07D1Re6eZ0T7JEx8P31ojtBO4qYxIgsaYSdY/HPiMraADv4ZvR5QE0V
Y3DmWncxYMcYBwWMhKekVWcHIHmxmjdtu7PLL5z47VAXeE/t8doztE6zE7Xo7QRkFeMufnAMxJbT
ULaZ+6fJcCcVwW6g0agqZzUw1voHW98ul6mhPbS8otNkY8kXISEUZwbpbpJYe3kIlApW4RHRKCas
zZzxV4Zr9zbRe+R0r08SKqtYw/Lj7i2Z4xny6P80oZ3YaDjBY+78UgU0KQqOAyQThvNeJPqonsjl
JQvgl+97DbKv9x5KFbQKqdrS8ltrCILZbIfgIzR9jSOdbOfG7Lk2Md0H8LZrF+UKVejcQhb0/AaQ
ED5RVhQZYzs84P4jrYrLjX/UQ1fBX8JjQj+NPfg1aL1s+CVymu9d8ko2RRPFqH6vi8Kba4ThTql5
GyD2mwyUO5mSzXq6XKSd6kADc6GBKs25L7Jv9qyIMOtbpmuYKWSmd9AAdYDhU40RMdWZ8gqy4EgX
j343yDnpHGMnGepoi2X08+GDRPFnFYUrj4WdL9wMuJIc7jiQN4noz4NzBhu/9I/6scxQ07rJnmc9
g72+tUEnMVnkGQ5wlAi+b8Hvxl7DkbDVV9qqd98eJws0Ib09Qy59Jq7CPi2l5F6pEj2Ho2CS0S+6
duF7LVPq0xpmTf4NCD8f5hjuofOI7duMXHk+3y3rwyCiro9dZVAu63aOiUhpsyD+TYbzDz/QQp8W
7b/26IGlR9+3sp6AgSDXYA0sgI07xGMTBpS6P9ZOZutOnBKnfF2FVjNA3maeHUfHoiqPgKUBkBV5
O7DWTm8L2IALE+cA9rGMsHLHn06uG8wB3BF9ovPi4J1qpJf/3cpuvnIDfsHjDSsipxGrajEbsLhC
9YADKy2zucFkBSqOpEjiomVgyqF4vVOQLTCyK5sGiQcO6fsPrBLNzH6lQRg4GJ9B08c0+EeikLmf
np+VRH2WKIZvXl0hySgSsPf27PSiHyNo0r4KOv4FLSI8vNuqeM8ka/MKQV5LNWXYsUI3KdusxzQG
6pxxd97fKVbi72rBQcJNjuCXKqL3XZHB9yOUsm/6fPdw0mRryHVxg6r0pvwBslyGqJQlTm9bJGZU
/91FmE6abBUwSxG/6UKeB5zM32E4AGsPOpwKMafw0zruLp5B5nhZVsdkS77mAr1NC0P0CvaiZyPg
DK2VoOe6dY+Wu4XL2QLpaIUgYipFAeNipMWqMyL7VlLqQ7fMy/sNIfB+XQkoloimbol3yTLeoMf5
FCGQyqbUq4LCXAVWz0Uk/kil01HK26fclKKfn1qJp+U/5qbf25hZey5j3dLqaK8eCBzJhPaqlK9Q
VoPrQLt/Ycp7IrkxDjHuSQl9pPeuFmJ94BNSLWfyeUVFtPDGOWpBUGucuAvsbGsxZPtYKhuQ1ULV
dw14jOgIILzKLl5+mn/Yohensv5MMh7ZqQWv4ANR3p2Rk6zZ4vkioCv7zk0k6cE1JapjuJMo4F+w
I+0/9FRMwKvAjr+QaDXI6SEjPAxOxzPjmmFqUItznqNo6Lm1h1SUL8oUdabbv9yH6nVDyl1qAx9M
0P5GBGVSRvLhkTdF0I6fDbzuUFrgAz2BFYNpvS6oWYDom2ZnfPMEWnERHyqAidp0cphle0fD1VlX
fhmOx5X9qx5N9L6dXHG5K89dIc5FwCrD/iZgaM6W48GX/F1R7qcvSVebGlQ/jLuJ11dNnExSSNFC
xYjof9omA6Bvh/2CcCU54peZVYOkufM2K0+ValrPThJyw8mIBzNF2q3tdisYiXsA1W8kM85L0u/h
+dYxm9OdzJBXxZZtLSbNZsqsD5QtQ1kTkoy0V8KbiweK4gtFhYe9AkNocEToBdubJEZRQ8NLqMgX
WmURXo1aJBDf81mLil8yOfErpWSfVM8yQNByBg4vG7n9fDHCky/Ft5IfLSUu0EokSt5SUOMCuHsY
F3LeMaBfjdJOt3iLH/sBgKOf0r8UaKvoHvyv9Nv+omuiVu0lIJjEs7k3Z9bhM1MA3pmksveUeKqU
Oy20oA6ba/ZvxHNwpEGCsUQ7ZA3fHnoslrH6cYAIqcC3yvj/ucTyyq8YY2xau6vOp2MgsEfpjF6v
WY74Dm654JITw4SDzdIx9LI0FuPj/8dcTUcb89vDAUhWntHhl2jKQlZndIyAi60BPP0ZdTAINt7a
fe3jwzvEPQmuoCEixAtnBSsN0jvuoBb84KGnKmLG9zcM3AYSHh1U9iK8mcqv8JZWDi3S2TXbdNod
2RtFfx04GMVw6P8Ud89yKibTnJ9ojWVe6PNVgZqWbg+FZbGiJjjzT3W7QibgxTasx88/FaNV+ckV
Jt1F4NGlqH/crdOYSOoUM8nqqZF6h62e7YgWNrzkOHd55uJT4bW9N4qjbnxRML3Z9QM+hf5LHGx6
99eOXCU798OxSmss2BQJUL0WOB7kSv22ADt9kEzH2wGzfco+n/Us/vrdJECp5WHYvmoQhgnOQ07d
64jtmeyCmg1bWnc5kKDF8VTEdNtvlB3arS7vfywQshwvD38KnswXSg9IJQNl7iJopy8vM7ashUjY
xeI5suIAgYkwvBTODzsXMk/woMyriGoFuxM3NcWqpjI+nzgNwCf9ZsNZp9QsZhQd4/6Y6J5VlGox
qcVwqLEJECnEavkP+sRrhvCg5Oo+Bob8pxeR75ccSohR1PDcl+e14OIJBXv1Lfb7vVOw+5YQaBZg
43s/ECPK8Czy4/oXV1NJ1h4x5dwJkf3Uo/U0pOjJPU8TEzjYgm0b8Y8JzXKBfYZDuutcVO47nB03
OYJU6XhFArYc+oNAOGkBU6iH1sDi0UyGyAVF0KSpMLL5C8bpzEgl+aauenF84qIhFRY3Hyo2iKYO
q5YlpdQJ2O7vd8yc745gZU8EnVb9gxW9Feu2SO8K2o4MUemAvtLcWkt8Dp0oEy5mvUIXTTdme3sm
SFotzNqNdttqyi2YS2WHYuwJMvwwVIvfY3rVNAeGyR6rgjxEO8cJdBy+O4c2hXzCFdi2wl+dyd84
p6HeYuv0N3H1nMgY0VhcpzYXeKwoU9vtM3+ukeZQ/5QOAyNZyLgD6Y0ItOyg+cnFTjkQ+B4FBMx7
ouvCV/V2vxwhQFPz0iZP8hR/fdAgNYXTaM6xLcD1PX5fLS71UwDL+UE1PO/E3GTzGYSKp6tpVo8F
MuJhlqt2mYf9mrsmKUQ99zeFjAJDZA45NbV4Aud7FJuGRnjlg3AfK05pBh9Wyt7Blvhhg9YkOsIn
AMbXzyygvdsOQ80zgMOXcxVKtlM7a9pkBPvGFjpOG8d3uEQRC3l3/gAaO4qA2Ec+iCL4IPZ6gBxd
Fs9+0h/rbMdNyd6esYCNh3uVH2She1DGF9p34f7lWDRll3bi+6YQJhalmQBCuMqxZbykfQ1nwwf2
5vhZc/7AzBVwOvCuawmW3zR5yROuiIgi+JsMQLGFNRypdGnUs/MVDbjIc1q7VVGC2vsXdzP7CT/D
4JJjU4X/WX7GCWlLOZ5e1hlW6Tq0pLgdL+W017/+I5KF9vIN3vRC52zikndGwWuPFmu3nr9lR7Ie
OtkUy2vuPqSFBpF9zhlEAz3/wB8CIMwENzT+XleR9TC0Zq6r0ngDSWEP5yvXscyLLC+qWfI7l5M9
B94cfOSmI92fmEWJ+7wvsz5zlZujC+oQb9nSh7ZtFW/gggW0sQ6ZJxpgm9nzrr89ijfvc5w85aTZ
1v8iKdltMXnJ9W/FemtY17/C0eW9X6OR/bWorC8ag67R7wd+jQ69UC2UKTl6Dv8sdVoClDZ3ysG3
iHYjF87HTTgBJnOudsDw4Bo97jHzTB9RTwXwoMSDnxwP/k8AgAkIoimO8mwUxaSmMGka8bFWCGy3
1AyuFmChg7gXwIZuVU2VR/YMLLgyVbB2PF6SYEtm08YrIvHoKQkr8sOKwh+zTlw2HD35Szm4gCeL
aD4mzZCDS658JIN82d6lKfruqHZLmC6ElPEanzONpYTJv6lYER1c/u4Cap0pNqRkDOcdRI2chV/g
yiOUCOp9hbc9WiLHzn0tITiKXg6XwNkJf4EI+uCcopVkn6EoIjubvQ254JoA3GnwW/maYjqxt/p4
P58U5fR3/csUEsWzxw25nU63DJ7QVRmdttz0dMbB6OGoBUmtnqiad9jgL2tvnpAyY49UlwNKOeWK
Tq0dldZ94Z7lHh37jNJEHUEyFO5ooe9IBy6dkLFI2iz0Hg7g1VAsR7e0Y0qvBRQjxhG1YpjkWgxb
h0Ti+iaa1Svj2p8VZBcNcNBmPsZgjCxUyHbCTxSl1ZkB2NvcXCQEd6EV2dfUmcLm0GZSB6Vr9xgy
9500ScxXJ9QGJPLQjzleLrVJSsz0XUfXpmcfr1qPjg7L+WPV0dz11+cCxsYxG4DAfnMkVUjHtVKf
gLYW6a5nd3Ea2csY1oV2UGGYjQ0r1LuaOosAgf991thqhgdfTQx/AA9pX0K+/nZXxDekGu3Xy6ir
iqmjHdliTmqgRGEqqR4FC7zz1QZh9jdXjqP2vFFhYMng6GLtb1fb24yOmCtKDXoWAaL/vlO5USHR
wsWGPkzer+8ApmcjOjbn4X2qjrG+wF2hdH/+ym6nuc3hOGzGLQ3w9Wxx/zai9b1o/aPdhklb02Tu
aPrym3M4YyFMeA/qQDtwvyMHquXU3MYIc0D6TaGq+nWDdu2MkluxmVNTo45ijggPekzHSSNr+He8
R0LGnGz6hTciQfwdgV6HLSPJ8xeTLFJVQDtjg2aV7Hy2kbd3pASzxDrIqPcmM3+vlAK1W0YVKhdx
cdL3AOmoDy/1QdfuOPbwuXuiWZPohEj16wxCLMgUWJsUgtOsP8Anl4jbResFcvJJOWz76tblw5iI
93adjo9qMS1FSXE+5Ony//lYQOny2d/NPWjujiSlrT3/Dh56wV5Qvouxpzqu6mmNdjcAsEn83eqV
bZ7py5cPlGDpJRK/zhDWCKoZmt6nvj6Ko14EnvxNDpUYkWu46dZxw56sr2710cBTnNkfieUQrLPt
vEvh2i9pBktELFIeP6tpUcScuoVCWkrkVP7oiQlNj+80vOHTJcJrAcex0VhzNHa2hiP9evLysPKy
7DFO6QmX0MDIw/X5SvLbCIYXGywW3qgQGAwDd5RkEyRLYxiQdYLeaXrCdMnTelJjxHfAEvxvp8Po
ZTPil1lNDPUilBEX+yItpxql6+9XxbLvjP7jNoh5KYfw4ipjqmt1KYmZzePLQg4mGElMHngmPO0z
krOnxyXK33EWDa9QuGGjNpWd6AhBACS/vrGdjPWV5/KShK/mc4CedkBr+ojl3mlmYkoKuZ0RekeF
SIZjyHwwPZGMzB2KRB5HaSnquETFnnlA4MDF9f9c5CwgJBCFd+7ujwMnEPOPRogpSL70/avC5bdN
caD3k+b8+F83aFwgGVl3TNUUiv4XUxF8QjO5iZz+a5/T6jjqzws2OBxKJzcp/7rBDwyG38QcIce9
9h9XG1LVexVhsZDmZkqQAN0ItHdyrFFeP9HTtW/F2pebAqBLG1YOc1N5seGVklRjKxq3L3juEpNk
GSarw52SJF7rNtcU0AC7EspamDkG10fckUuCzWuIKH0UDoTVmkCqvfbHQm+qI08jqSmt2fik6YOc
0jnpNbmJe/pQtK/TiH7Z1vqepoZSEmTaO12J1oTU2UPXOlNV0rpbDQm/bEr5KcBbvuqCGOxSID7k
XsXguRzIV9vYBcmKPCbN0URYsWlxVkZoGu2lZcgEY2su3neFj490kOcDXG61bxqGzuYh+MMJQ+y3
8vmAcWHBx+Kq+Jq/bXAPBIs4OQkREemIfT30Zm4D204dEzyO9AhFhckl4U9kyJ2boeT7PA3quVqJ
AYVvKu82zX4O982ne7kvl+iGOl2hDeX0/VUVTxGwPiZcTHkrU/tL6Bd9jYpaLN5c1AVdDzCWxxq0
w7ukLeK6NJUHrvG8z82q8pr7iJF71NcoAgrE04/xHQpl/QRcNn46fRMAoLXlbDQw0f9lPEmOt6AU
9crdc84ZCRKv+kxWsQGdkNrK2rnZyi47HWwmAOOF3HPhDmC/KSEV1eeQdb8opLakwX+6M1ZHZG51
rmsQR/vxK9/5b/548cgTXeib6ZEthSzRw+iHOS69g4UoeykbArOxCst9yRyzzDmmiYWnLOaL+1nd
Zwd16OdQRbmxqwvVN5HNfRh+0reCnmHz24g5hhdQ98cCsk3yE6K02F0mj3+1hHnntb8f674sCosO
Ru0ZHekx6Ccwtg6SazR5byXiFjc/vrrn7Fzeira07s/H/8CAw77KeCPChOzbIuPBjUO7DV0oa0Vs
ZWeN5FysBWSEAHXmq8PPmt8FFvUSbd6YBl9hQAUG5kQsTFzaduZBc8E62ocnPx7Y7P8FQ3nY4ntQ
M83eAhhSpNTQNf908+ENTNH42hr6D4VkkIGBsTXr+JgDjN7COsPyvT6gl530xU7bFZIcaSX+Knjv
LWhCzwQw+nx4fQL5XFC+I6aBGRVlv+S/hAlDdl9Orl3Hd5vdCrlSD3FOteilJS//Z34yDYHvZelD
VB2eeX0lSymkqi3OSz9P8xQ4JpLdLosNaulcqcyfuXpT6UOgog2lCYz50KGkYWt11IMYrE21k8UI
zw9OdTTwvIzo1eg8xP8keJCewC1yMW2sRGmWSRQYVEm/lIUu8jcNGZtpUAGMknlglp7ZyJWsM9Yz
ZZ1DfWrRfySCgZAM7EMJzrsNQpKWjWUYQ8YIGL8rtttt2zUt/7N9VXJ3/0TQDywKhsNMm2dKrt9Z
tl2+nS8SwjecIXyRFxHipN0qtKWQYPbPWJu/pUzCgpePyjM3EfjzFoEYqc2g290sZcPTZ29SrfNd
yL6PKH5zbx7lWDjUct9mKSwX8gmJfSgVSRKAhMk6dS1ABMldwefINZ0hN6o4EnxSbp+2pZ9wHeR2
/bM914zUyuK/GKoJjmhYAOwjEA+IYFdUgxd12cayDJd6E+N7qVBxelOddR9eb+M1VouFIW2U6Q76
SMasCVW+sygSQRCvan1QZXWxb51Rz9J/6hm/8Df65/g2VGvQeeEqs/YT8zwspI+lpYGTdowUyxpT
EJ2LTDs/YmRbqvS9WSE1fwuCAX9a+6EqjnA9rYJSRSqbT5c/BPLcEEna4mh9HdxvkN7xTxShG/1k
b8UoPKfDdG4oVDbGQWevxX6bLLtgmSrHlYJkeEKR6XoqJ85ppjSyZxuDYYBAFzmovZ0hOp179eOV
XSRksvf/31rhsSFL5X3Ksjmf1WEasfB04YQtfkD8nsp/2OtwNFgJ8mi4p7ksXs0SsRgW+4qNoouy
6U6qhdPxTzMff4an0etWr/9EJXSFHeknpmmznxAP77TmQ/P4CzLTQkISMeHMmXysD2IeYw7sPNy1
Cr9RCWAcVCTxPbQBopANvRUZcL669jrv7Zw3Hib8vvpib5qKJW0H1JhH1gfhClVaIpcNuuJ1sb4M
SGgAph4wStg5pfSDHyX/TRbyoHlrtmvsz4775FrPVTverfSFspPG0TJGItpZAvIcJFBs4zGnwzqb
9M5883B96yvw4TZnK1vJ2OzW006ZD+o3UEwuF5VNYiwJ/JmeNAfh4feWg1A7WtSlGhCXdt5zjBbt
TUVRqvZrWuuRKxWHXwvwDa0oOovJQn9s0F/rvuirEz8+BMzUT4LLiJvqONsGiaWhEz8NsEKBiVph
jhR6vBRQ3AQM2sbwNU6cPs26sMt6K3XGou3Kk5lwCWtpwjoATCk+HaiH6HS4fP64eWbYdjsQ7HpP
JEpf/NVneoGFCMbSLv1tfniCbyyhE2mlOUUtE7yxWZn1yULagj4hvHUqleFd73c88vWmx8CAhGjd
OewHZ41NfQqeZy2Y0xcTUB/Eyzj/fuTY6u4HqbaMAKhcUhC2diI5rbGzDxyyITSLqW6+puqg6wol
+vbVkQyISj7yAnIeN6lEoOxQwIY6mQfCP3jLu1xoZWs46sn7pHKDxc+HE5gH5JyCUGrtAa8+Ju7l
kxhTCD2DDbpssjV7XtfW/CjAX2qU04iNVTQMDFhsy4g/GdQyMi39avGjVsbwASIai/yCQ157ORbC
1U1k9Souy0sUZLnL24Qp30EoPicNCrKBCJ4/a3/1YTta0FNZWvD6MvKDteVi4y0UDIVMtFkMroMW
5Xr1Z/aHQtoJZRaO/5g0srkUJ/Oajj1Ot0Iwk2w7o7kRd6N1ssIlU4CInW6YRIF2tdGGD643aWLK
/PxgbJZKayTixIy/dRpE2ShtUV8qF648g1QQVgWUEjxpLBjsqcLcw4JzPHewhvBtc75pESiDBZuP
NvC9zKy3+Rn60Y1r7Bmr4LuZlDki0kOkBeZuy+DAq+J+UBpNkI1pzs+8nYgOsMbZzStrjVVadXsH
Yioew7lfxX/O1BAbi/l6VJUu7UfMmlyZFuaz9UOTNDJpy+8tUUQ7igDs2g3++Mm6z3igLDt9/cxe
QG5d0hD/tcxBIP/Ppuz18bdKXY2JUJAgZvoO2WrY3LsDnqzjAWWmWWTHUhrr9IK/qUQ51DQlQ0PR
ORRwDvagU5HQEqQyg6V1ReeTF7aLly7LZBhoWFst1//DTdoRllghNSzZmpZ1Ppb/Byv9Z567OeMG
flZPqFSOyKnLh9u4Q4vpUfJh2XWwwZQr2Uqn1RT65T+VcGWTW4ETnuMkuqyhUc0xaMx3nMH0mu1r
7WiFz7aOeRb1yd0muQZct5arpgmkRaYHoD0gbg8jaDboPYUqhsWynPQQdZ98pDdWHwT9+5a1vgX5
F7TlH6kevhUF9GJTCZ1yKteyuW/WgX+MdbgVN7sC9EPO6NjQ25awm52B4rU4coTL0GRxUiDk6bmA
5nc2Pux6FAhseDIxGCK9nX4oG+DV38Cny6qOyP/pm9NKldPIoMeO/l2gVmAOuvaxD+3uJAIZilLA
EMbpwZ9BcDOrJe0GXpIzmN/kjh98F1Dd/msLj7982Lligr32GpiBQKq+QbxlQcRdeG/BxG/NqOk8
eUkoRQlx3rvW2uYyJOUvK639ZXWK7nO4mMdOi4QsviYEhf5JZI2ReEwZeZGlYQz0xoRa5bgiOQf5
CzAMErdcvTXui3cF/KIXm9mLWaJMuopzmwo1F3SBbEfk0tX+guxHP/pki/UTGE5Dy0bVz50oF//e
H2s3oKV9h9s6st6+0f503R0dngey3w2TFv08OPzLgvPTGMZHDa4r/Oajg1vM+pL7wP6/qXJy+55W
pkShjV6elMayUPuPngC6P9HMEDDfRsV6YMF4iR+kxuJPk9ZTjngEf005OYQt0iUo+PL8+e+aInJX
a4o2vaGaAo4Q3LE4iPRtGZ+GbxpXcS7HFwK95fMVfI/IzTBE5FHBZvL9ujTZXV0uIgVp5AqphoHL
AYEyF0+9dqiTrp42BD9cY0sjO/Qawbf4iTT3wxwFdCiDMfCbyKyiA1tL79HdKVm2Vg6Vfc6b2kCq
hi5z4Rwp/sctpDZzDCBJtVo1BYxbQLQzpCoHq8ODx/OgiHLbTzTH4JAW77HRb4IPv7i21FyhdajT
D5cMxhXUfkL2v5bXjFuj6D98qSqNiiV32uHOl4NZgzgOiolp8qj9IEc0jHcYESC3Msry64dfSH6U
HEcCSUzXDnXJboReULMluejFBaW7J58qooS+Kqh/eZU9IKERzULapUV7dNqfukHX3v0PxzqXJQGM
91WlYRGMCk1WLqMOIhn6Bb0ALJrNkDpF9uRAbLTVQjMzAun83rWKtp4cQjyafe50NuLSBgGAHBrO
hV5kJQiSeiLmXV2/eCS74UtAmv6TQUMzhWx23uJom3XELCfVw1KAb+7n8o1YNsX9faVBn0M7q5Xm
DkDnqqcnyrWfilVzJgDyPQv32YFcduz4W97X13+q3XgJ3oGBXh4nRGU1LAjxK9UwoITzJ3TjVZhi
0KIk7oSAn0fFWdv/156KFhp6EFiSChs5eTiXfQ2T0TPB3Uy7Ln/jN8THll0+hrvgnVrJZHCTVdza
P5vD1DMb7vbIsWoczIE5JhbiJwpjWao1W9uXOfe3kN5IIUApHvmT3oKANbFxaSsH7R6dRcuz/5sE
ir5ypUpgZHNi2SwAHMxn0hAWdIVfC+l7dorScg3BrrWIQUc29dljh1R4LioDHrntiUigw3EFIcBJ
MR8k2ILjLY9EOP0O+ql6pSCiqCNUb71xgXyrgE8WlUTfy7pOWrI8xut/PfkE65ZJ82xz7/fDasWL
IFllexYt1ytsoccl/LgApE4tzOdTCreTTF6wQxFKT7IRdRCRSzVw3N0Ug6hHcMyOM89A53Jf/+6l
XT6hlsh1bREiKdWtdtZ4dwBu9vgM/m1E1cZL6oyF1dJHnZMcByRp8V5TcjAOj4Eb6LfOJeNb8ZN/
ZUugfbd8tAWZHP95ejYcoVsTk8h/mnAUVhuHjyddRXu+W2hTfvf6OHvIk1fFKGuvbqhGJf3szHxd
5nJBeety2PhxR1cV4wPEqaoZjtUXPszmgcVsNTeSGAbe3Xaeut+EcX24GNq0xwQkWG/vG6p27Wmn
CkW1k8SHnJ3Oe1hScWt9M/JGfcq8X9dgOiF6UAIxBrpOMfk0oiOOEuYiyqgH/lAfouYcwGPBF7/+
2DmLXqnHAhTZd+KL1R2dED0NiLFnqYu+eQEFs2MXdsFoY9P1Z/IA4h+ooI0XaOkLFglQs+g55n2H
wLnXI5JIO1hc/sN1b64vyHdbtCCd70Xpxo8rDf1WjAYlTTqRkNJjTvsPbAnTFwp3Oj69ClnE9wMu
BwQzB1tbsCuFEtwIr6jdyyNgt/BhcNhlYp0y4Ns/0fnW4WBr5YYoX8sl20EUV3EGr+5YvCbECmH9
XPo7TRP2Qqkb5OCZv3mfm3ehSG+CvBxuMfcy+iDcTTuL51HDM3yP+GvC1cnWFjye2gbh3GOrg4du
p/6Uj+CQupDeHgDz9lQKTJvCKXObJqwGlg8h8AM5SE7Ce5mD0dbB6MuB40JFXg50lK0ZyaXNoat6
b/0ZzNeQa7rPTey+NELZPcE2qVi2Jhw3YkKBFGlexeiqa1Cf3IzEcI63bde3qvbX7sQa30DHkaor
qn+Dq80/O9bvNU3fskCEEKLsynZO6WIxbxRup7kWYiB57nMWzQWfp7jU73PcYdIWbqH0kDpZYVtj
+AGX1cjKklRjGNYrJ7/9Xg71CQCaLSjQc0Pl9WAwiVCdxujwAR9V5V3pWCdxOsMaIQB77nMHkVTE
l1Ya0yz1OXuqeKi0uCl7PTz4mVvKQSRnDx2tExB+8BnKnnV3AsALpC2alHGKlDxVMxyymAeUCZhY
6SOm1vDr+6SIo5OnngLqGfjHhyLrUTREHgPgr/uZ/laAYxOTqRrE3Ra3sGmYxh0v5k0entItLfLt
PCzRofERjHsO4wS0XJrhfledrdREFzse1krDW4WYskJKmR87SUdK+38FCBlDt79QtlO+tbo025DZ
GPxyuBB4DOOnYf/usYs9cErLa6ytCFXqo4xKcRKVEGLCYmrCi9u7Waot5CHADcoZisy8dDoWsIq/
cwe2PqQFH3NpoOmnfmojRb6CcPqPs2Omni/qM8wyoavmknEN2aqXkOD3H4XAD2zFhREaaqgoVUIA
o3qmLIogLlmTYGvNz9n5XqYlWOEchPieh8uoTKg5yFxjgnpnv53YmbqJIy0bXoJSBwXZGgEsvuXX
+6z+K48kntnNh9NQTfLk1Gj8eUt1v7PVdcgQxsFOu+biOrb1IWubLsV8uYcBxVTfPZ9s8BEmQIwP
eEbAULJqF15UPb02Ndtzkc0RS+BjiKVNSql/gFRNXPmHQeAy2dFhMRpXFRfgZ70+R3bojQ3xb5k8
P06GCTvBOL4fSGzBlw2fMTOQjH8qGip0uhMjhFY3e3IfJqMvzLEqbeLJAKitJUcLAlEUWMj0/LaT
3cjMGRRrok+fqGPmdH7XexkVLSY7XV4tYX9GBMAjk/TM7INNtiPlUxXklkV10PE3yeBEP0wHLVfZ
n7qP9rCvnItg2/ti2KEUw4EQXkZMYQxAHfcWWK61bWyTp9so8MmkwB25AI438y286iwE7wP/54cX
LJ3wICl95kp+osJ3FFeLgTRwP0eh274ovmAJ4yOS5lP0J4sUt+zoypD9+gOy3eaeVoFRkF7qiXFp
9w2dl06paJtL6BdzWxRuuwygzVGOF1/t6F3sJUdC4DNLSzJyawYD91VUm9PhMC77hbHcr+6ApUq+
CJb4dL7RbfnlUqZ0guLNij0fkVdbffmKbox8QWJe5P7Lyrp+HgiOhr+YjjK/WHr2PjF+2I2lp8rL
Hem/T1j3yJF2rL8OuvPyeNJX2sljqnyGFAaT8wQyf1BIb1TuyJYtVBaajiDQfDg8RKWgRi7xY8UW
jSEyupZkyV+YBoszKfncl2GZsqkMtl0AU0ZeV4I8KmERTszDtaKUUSpVGs+Oksgfszi4PaiJHRdc
E4AbSWjrqiSWxMN/jOSx4uRkWOdOrCn3pGRAtQAzxr7lHTKMyFeulDNJE60852/Lde3LDZuWoFi2
UhwigTnFgMQerN85OsUaP4Ii/muLDJYawtbgGpihqUZPaLTO0kfiiYGjuMGno3+ad2iEE3n1iyJU
nthcLK1T4QRltmd9+cM4WpEBT0GFft6b5jrhzuBdQzT/m/ywAwvsvINH1BtkiTrR2yaI3lm0o+fO
hRm5O7+oGeOHX58X3uzJaxUNL1XTuDWOfpJmc7rz92oJz+qNaTImzgxPVdPhB1z2gTxGpqSltYH4
vALYP+ETvxzigfve4hjvHuljuK7R89EyHm+CaObiW2lAvNuCC4K8FA6LbdMzDancMx8jjsq+S5WK
GmDr6aQnV0HxHB8AWnaSFGqFvIJeLodkzdkG/wnpx4Ir+o7boRGd7z/L7VuaqejYAC0cSB7Xh9fB
JGc0DSPNbqtREvHJ8yvB9xAi4C7kYLWRT/rI6mQ0mGNV4+5COKajOv/zFjMm1FmsN8kxGJ+m0RUf
3NEdxb0LPUx363yYc9dw9p/GxgFpvivWBZo20+78xLwt6PA8tUQR7nYyLB8gO637TqAy9g3aE7Wr
XP8U/sXXulwxiER9YcKWlx/z9CeRA7lepEJonHQQT9GP5UmBxsC3YhlO2Zbi41l/BBCY8Liref4K
h8+9sdL2uKjpAFIEQf8TyBpyMZznQI/SDXb4Rpy3ntG/h8Z3VOCoxoAu5/GMsU/EI5Rp0BltPsGI
ncDRX9hxShowp1Xw/8REL+rY6Ar2HL5BXYZJ2Iu6ZtDdO2SMiywGGqQKo/27timExnNxqow2lZcn
Cq0RhH1v8u53OVXpFWAuuVPJ7MNg+DOtdPB6Tvj2GEgvUBbI+zLXUXGK12sZOx5c9e33nFisGmjH
vRjX/1Lam6qrHdT0mCAUSIk7HSHlg1PhY//NUT9nI/Hba77uAitntuxqH6PM/i5LhnRmD/QaeqTE
NDiOxsKpr3Qsz0M1We+2oa7kTFj9AA1F998wU+dGgpmiMW3/S76/JioNY5xMd1pKeSPcfzKeapMf
TJgBU9/tpAt/XTaaoxucY5jIXr978Lo1ZwoA5sgrMSC1l/7ke3J513hJWKs8M6jMP7eoeIq0qTv1
/vH7OMeMKiOHsC3U7L4WIoS3MtQ8kxUSTm3azme7xfJtP0WaaBuQFhEIVZDwe+b1wa5TZC9thnD/
E3e0oeiQ5Rw7h/UNHAMT7uokaLJ2B48SHYjFw8G3wuLCaVmTa4ehfRoiHNYHYUftxl45BcxCWHSD
Z7R78ukPV3tX8lPZ9jYCJ5zy4WvN8HGXkhODsfAqXLQPqzRem+/HN0V2JySBQX2SDrxHavRRiPuF
BJmaEzHzlwJsU7HvetM8Fu00weZzi2BJ3dy0q2/IjF8GRzTAH1C7+/aOLrSm8Hgxl5EstPytBtOU
2IoqAtxFeOe4IboZ3/GnN6ihHOOSADZwMZbIgGPUiIxPHJLsxBwneq3QVMXAuyGqQnNKE+uEDCNl
vby2pfh9kuJLWyFqVGp3FDMfi9YrOE41Tjoy9KuHm50MxE+t2OhH4Cwn0AWwjLedh0JSVMR9P7Ru
TE7QYBpI0kF8VGC3BXW73srOfhuwS/0xzcyE8DoHAL9wI1UN90blqbytEDS+gHmluwL9tozkZN5M
J6xDoZu+X+oaZd9aMYHu1nSZZro7MiWKdPcNvNR/OrR3dJA9VIyMtBZU7VfYrKPvMetBURaEQUkJ
CyNG3+/eVADCj6PdYw8Gg1gF6QlrZK1wCDWeQGfSV2wzjDtVrdsy4Bb36HJprtWk57SeJMImDDZs
BXPpy0wx/vy3xpGtbGrlX09DM4eowZdF3nMiBN8hHqTYewqUHDnwAhWfXUhaXOFQyTOqEGRdACRt
ui1iP/welIcJR+MbxPqL9DJFemXl5ZzY3URINVzBa0tzO8pZThttMGGNG7NpUlLa5VLz5DRtnij/
y9lJ5hycEerVGS6cQvbtz4/CMB+TmAEubZT3RdLfJEK0zC4yourxf+iEzxvHtSXL7cm+swyWNCv0
ynqN2iHDuBlLAExRz3RazDknTvQymaIvb0DcS3OE0TwqUQWrgd6DZhUhvdtDeeE3MvX4nCpZ0dy6
qJ2VPFGL4pstWZVcZRfVu1huD6IIOrgLiuvuPGR59oO5GtWfy6BQBxWrjLCnTc2pve10eoH3jXmL
RWj4UF9h3gk1yWuXooeIkgjMmLvusi0WcE6Y6CQOMOT4K97oQHW2JIHF8+iH6BhW5XP7LF6p4R4m
GjkS67+16+nk3ehJ+BTTu22FPoMWqAEtDSelWkydigK8lCz5thEX4uohW/9Bb3qMzl+rIcM8AFXf
1O43axJp0H9KWfW7hxfVYedBkeAXH/55V6TkvwQgwXmolPGB2yKiOrYTxtlceTktv8DyAGTJmOhO
TDWCoDTxplkTiXiJXmRUAKYDHh/WXRcIyrC5/D03P2zLQRF4x2GA1Jlt26s3sOJnN4nInkQP2VwV
djO7G7vTnLZPI0dw3Kwcqeu4wup8BK1hymIP+BX5D3KJXD6zHWvxqjMhhz3fomjv+8BT40i0mbi+
ZvtY+5c/Yuc+NxJhgWeAJF5gafe4lfBa35k6Ty/dfkNZ+dGa6Mmmgsoy3pOFJBoJJcNKimrl9Oig
XtZ+QUMEMct0//1FKUui6jEJjhPzsHZZgi4k7aIVqknOsXgGMhK9CT5LVrg2i1kd1e9FxuYt0mbf
uOQZ8c6qyDm32QYs89Cy229Du9R5b5dSl/9nYz3Pp11YQk1xIc/nhwxtGewjKXZNpIgENS3fVyyh
fk0vhNorEcrFFHuKp40h/3/b7+oyyMUrSyn7q1uZMrK4BN2/547GCL7py1+4fFXnc+MiOahRW6G0
SJ3F88RX+Lqu28x+3LIKED0ytFLsjKBxhbkfyEYZ5Ze1y9kZpAcUd8dLQhnMtm4R9guvCFslZmAW
5vheS+3IOqumSAHtqQ0MdjvGRw9xPQzT6lKLxrb7EDDlkWyXacICapU2OWS5bRxzm+bcT59x2Mev
rVMn3Oq6N2gcjVZ06bhlaKrO2I1tCAqlN5TmzCAjJ2lVFYYDotnWEHgXbMn27wzAnfQ0wGgb6Zdk
MJzWpJwF5Dj4LzeoGC3UdRqUHuJU92bOPhyYc46wkWO+OOTRVi/S0sjT0R7sk1HNfrsZa7kG4lVc
bA7uxZ5WAwFAr7bEpS7kCwHAqxOujl9fpvH4mKop3K+Zkm0zkhlQM4hdOdsaFdNBdS0HnuZhWcYN
YIuNRg2o+bl9B9f5Dl6wif4VR2fcYSbuhWqz4kOBuTcm/UzrdH6fWBLGjks2EZoHUa89fidSwlaD
UjrDzllQ1ukeusIzq+mAsSX1pTeSvnh9I68PoAtnBgndhbEb5uh/XsTrLJcHbWf1TY/ctv0+KpZO
agTFEJcQPmVjm8ktMOodyI9rvmfs+l3KptdivZ2bFmWDM8zveNz6MwwOf+/Dma8mZHUo4ggGOOW7
toWKPp6rUulVtWajsLU8YfQVoLe1QqWA3ULvE2DDV3xSmhVTVqi3WHDd5PDS50elL8Xofvg2HKuQ
TS0osVbgO8cbo3UY1ly6VNay8VYo59N2ViloIbkEV/Q2rOle7QQm99dY63jBgcIGnnvJbKDFucOK
WJxbWl/lV/sGyRxUFcwCm9SdE8chv2UL3eDP2xX0UMpTYDIJpJR6L2g67Qx8iJF7/JuQS60m67Bi
Xx4T3wOpx4iUAp+vjwdcKqX4qsdSg/3H53NDRDE/7c0IeWVxtqjnHilInKvSIPabVLTGDqno6ca3
knTQI1FMTnHL6GthJx9O+WL0Qc6JpOgdzPxMzgBkGFZnFi1Cjv3158tWL/AWupkZnLvreo9Llv8M
EYl+/t3NBOiezhKQsBMBgHOrZAsicBYL8g9kzy5RnzzN9ESsJELmzNuWZAL/2uPwntPacoN6uzMP
HrdIoR/iQJvRSYjQyu8Pkg1pOpHm4+9xpZb2Ia6/sYJlEcCv2Fw1Ybkmv+yRQjgX48wo89E2X88H
ljbIbit5K32bRVYp9jfk8HdrjSW7LJnhzGvebIeqcDEpgDOKl6+KT6oCqiS7rmzcTMiEJwq0kXPB
v3CPfD89QJ1zRZZ/s/BLL3a/SmNPiIsPZjMEeK9+waggaE8cnAx2JA9GcGVFVqcLvUTd7DNBeWjz
38lsRi+MvgjbRSoDquEA0t45Rc0vcb9KbEUgadmvY+N8NdXhy565eXxXLjNrUaaZN5dop26d+wee
06yT0x9bOBwA7elZ55ZsRJQeRaS2UrrUHDQYCzs+gbuyNRPEXAe3KIXTjOudQj7kbRFC23W1yg68
qoAafbi5TkdofnxfLBilIwXuwDLBSfFESDwqoUN1gQ8VXjXZChjSqwlHKg6RMiWtrHqgZwstTJGm
j6olIs6mHXLzIZRP3JsXlMS+XrzBLg5iyOXRu6th4cba/SDQFobj/IoAwZyLOWx9qm0AgPTCrkN8
zlbQ4672QBDhbkh91t7h3hBBUpZRYUJ3eTD7lQE33iEBXvlhVzNaFJlxoX9Bq9TDLErfawrFCvrR
moOXghhrEfptry0SCNW9S7hEES+C+J1vdWLHHRfDhwZgnOOq8GdzEdjzX8PlnZNxNCihx0/BU4HJ
VKy5k2ld3Wu0Z6mwdeaCAbY1XRZaIB03iBobBTAiqDJP4w+dwAYDtSL2WZmngKAy3HtbiypgeWq0
ODdr3Mho/ATjSZnH20YVezkaLABgIxgbMWag/WjPVkNU9FKBDM6H9d3VTc4+Y6vfChbzno8ZV+Ox
gz2hBOuXp2vLJYYthIT6z8VhoCe2p3OT2DFhbvmjE0ePmmoWLpNTadVPC1516Mq1lEHiKwrmtjQ1
fTDLLc83mS/Wwr7wMNpoXap26ws1iR3V7v4SLe2wnTaM+k4/EVbZJ/y/iXNiBcFz9Iodp4+xdmIC
7O4Kg4c1rqzIdTyB04xgdqiJxqtzXgfwmxA9+cx9c0ah58a8/1CLZQHXqTedV1DY/n9hKgc8+pzC
4i1+dJihIG3fTph7wqnDmCt/RBaK7Z9S04QK7/cxoiA8tVNxZUceRDC6aLpq5/xvBCUtec/LRhfe
utlaMxJW3YXpxGJOlydI69VjPC7cyu0gR7elRoK2zyMQ0ds3PQq+MCuKzcodhyRiU7A0A51q+keQ
K2KmToVKP5bqQErxYRHiX2renf9FW6V9IBi8NJ/o4M7q38mB7vojg+fYhc+HXu60oa42nUNytP+D
uJ6HRdKEI/th6Yqj8JlghNcjR5mWJB/aSYiE/KmEF6IfgB1MCSIw1Rh/QB+8oilC2bHjuHJ2Usio
yLKvdUy5HeNWI3tLOVQ102k1kCFjvFQHbx7i5LFdiWClBj0C+p3k1PewZnGp4azT67fRwDSpMUzY
BBVs/AnlLEr1rcPtTO8rDpIdTSGZv1CwPdUd8dT1t0bjeQckI3qcRqMsPjPTdjrowVEwuH4lWLUF
nBFkyGnSVGFmBt3M/GyugR0TZYbFnU273Y1LjdTbsXBNV1pR9h1P0ohYGwk6YnkvjhrXSc3K+qew
vqYg4Y15X7j5shXynF3BqN0pGblBtolVuowT3cOE4M3xQbfI2X/dhc6A56PA8WY4ayWkXFo7cGDc
TS6HqDvGtMsEc4MMBdoSO/UAs3W8sdbDK2xC3boh/T51NQPs3rxcjrmMzTAo/J+uMsEYAA6XTACT
aWOz4rEFk8EurlI0xiyrN3SlrBwxSOQRAtmhlns5Po2Ojihk/poFOjgiZk23VmizSmMOmZOCu7yp
PUpxhr15YfdAiwpYZ08xeu9Bj/YbGQTJjxPi9ezv1Rpbh20BS5xugdy1HkdiZt6Fao+lkUs5cGdc
vyUa3VwBqn2jwh9rT8sPxcCU+S56pmESv9VcWEdEnbKmPGVdMPKxlZlSZsfuvN98iStjDz2Oa6rw
H7oxCtfuNLLwWJyt8BJadQKwo/Dlx87FyjAEIT+bWogJF6pFSizW5+/h5uAhPunzZTV2t4ydL3vj
IFNx0PEELmRY8y9HoAJF/45/t67sEn9x3kK1ql0HOD9bgI/Mwmti2UF+HPhQ/mfPr7E+pgjEdwxS
Qn3r6iaOBuDX7I5OySB4SYyGf8/So0Rr5EsCQ42BjeRGjZFGNCmgrm574/paRuWLd8FrDCRVen+B
ARPFKJzI00lwzBYXkdMXMDEQAGu7wVg0ddoCUFI4BWCU152ZHjAPIWKIhNOmdPmcHTczGA5FzlH0
cJEDEuO7HzFWKYaq/9GmgeO4PjvrhjcZmHRRYBKvgnGSYUnSZRctKLjqOeS1Dn3r+MuwmVhwspt2
e9zSnKwrueDZWfX+tnivTX2mQyawh847YMieZM9mH90ytP3R4yZ/0vRAgI7/Ajh5LRWko7IUkMHp
MUMceHjYO28w0RlRYOnKOhsJP8lmpiH8qPIDIyaAPjoOzrDoapUb+Z6gDpZyMn+1x/vP0hSdwOtT
POaWL2iXxTimna0IbmcCXkkEqHw9RGbqpihXlaAwneyMlvHyimoWiH7ubTu8rWPRrZ2yUd4MrZem
pygx6yy0oMzVubo/NY+qB2ZAHESLJwA2CfdZaDxxIA8lg6y2AHMOZnRvlJLDmNsSYzh4rAkhzpBm
GG48/Bnlhet1JzP+b6YDnw2LdZaFx+rTPeaXh1as66ooso27GCKvI+A2/P1BPrIGU+OdTVfux7/f
6GyYaQ7rGTo3oKpj2EOir2LOZ5IKWAGTvu4OXNq5dyjzm63GIlvOxFrTa6nIWbqTccVysoLDYPKW
wb0VcOqbWdBlCKqsM04kc+ocLDx3mIYbCBLHNrMsxMHALRKDRuY4tegLVKUH7nYNKetnTjkwONQc
ngx+C0P4Uyu/dVK/EttGY3SaJ2rb42sgEY+YWqfCtkbK2CW3IfYh/AfIMesQ+yX8LCbhPDZbgxTm
KE4M1jjVb4fMVfg4+3fj0oQ0E2jOLQCzlF96CPRMEtE4mi3CGnRxaK4Rv2gm88eyZcz11uM7DiZO
iTgJRNTqMLXWZCyQ4dq+0p+dAo0rhowvecfI+nFXb2vHZF1b0/7lURcWUfibFDJbT5VYSjXatJ3b
qbVc1huPolwPwKMlIb0TjSOi6xNbk2FQr58xmHMdaH60c4d7L2b9qMK6giFEhT6/X5xFaT7ghKzj
3lUd3XLv2G2rwFAycXnoH+XV3iJ54lufsp14gmcRE49YDvmTynZCNT2eENiGYkKZLnkBKsqmwxmt
1IjR84KPug3ADUNbeiVZaKBgaOTPIvd/lX2aXqPFNA5en9eNuua9hr8gpkLWMUcm2u0NK85RJM2Z
2ld4Yv6SJi9nMiyKZNGim13Qhud8l8rb8J8+D/0Cq6Plm00iIzbFk69GaxVef77b3WuPK/F5rW5C
NvA5AhWt+qvXmD+EkWd8SaGkKIMru/zlAq4OyCKY23AOcMzs0QSZlVpjnhXEJR/4dkXV4HZO9zfg
jxDFymmRirswDRLmcWMJwSSV9j1krbDutCXHzdjhRTQtXfWlp0r6peBK5ZB9H65iW9/KoJjoQOuZ
eTmrbfltUzU30KmgMMc21irB8plaR5oItpMrJ/lfrB4wGBJgzPLCDlYwgTUxphNsmnGcxuA09+ee
VI6hbk/ZtXIKkW96qcz0zM7jctFzCN6T86SlACpQ787hpOoIikNRW/wDb5qBG1wcBpEu9cZHQbCO
BJnLbfNTOVRWsI+jaAq1rnuFhy5YRZ2zZDTzvrsSCk0QdYDcTVTc5zdS0SyVPiZPq+i/RTlUCZtw
1+zZ/vUHUtN/MrsaGVwHNzYkS+mAPji6Xzb0klxegZO6vByQ+wL8m2sG619GPL30zGGigPX2bzCC
JUOovNCytGvpMgjtkC7S2/U7DWFJfJFoS2cR1WoN/jsdZ9nZSamVeclfeWKCXxtne8Pfgbt4owoU
KB3AOZ0SjaJtgVF4kZ+DB3jU9rln5bMO8o2S08CJma0eP9j56XgKgql/uBQXEL5IRnWTUHMEyLU5
uqA25jcv5aMiypUGfrFFAFarbmvShRuQVXir3V8z0JKYtQJ4Ha9A1GFuRugdJfT2LQnHRccDaB5a
LIO8v273yffZkDvIJiesL+e00JwC1z1arJFq0C7eF8yl9bRQEmB98EA9yRhi7zyN2vhiQOUhBUxq
rZYJeiCWbwRNXxW9I+aczZQA6ZrVViildUCP4CllOXIRXReIph4bJG6EbUedSPOLpGifiMp7jK41
LbvTVSrEpLfGn35773TmM1BstDymS1nGt9lQKuAzmSjVBJWWsAFRXlSyd20xem4w2qfBLlOQwIyu
e9HMpf0hHAihrZ4O5fugEr9S1e7aLys0OUz2ZBGEforkGFKVI/PXboqLj0/pgxDfdR1WMsuecemz
MDK91Ve83/X9CcsLIFSUH763gY3N+WgUa/TPBPcf7xBiEE8+sXFLVEpnDcOmJIqGAm0mDBdMDm7a
fYTAftd2NipF4vBimHHxbZLUFd8i0ft5Y7w27mvq7qiTO+ETpziHwh4kli4qCArhXVkcOmpkm0Hj
6vRsa9v+kkPnEyIS7NsWpkZIfgyhK1IY5RpseouNyq1hG8odu5KLEi+SrqkcBlPHNeb3CNbmRVqY
Wc7HCq0jhBOWuhgNN73DdhDBricKOAZiiAIk7pMZ2C6+Lh49c6RT0GyIpu23AD/ImIfisf7Vtk4R
D8Ra6jtGhRtPPJN8RGMF3P9WtaheHEE86sWnwxExCFVa7tatxT3k6v6y4AMVChxv1ok0vfuwC05T
qgX9cmW+RoVfvJGubca7PIp0xF2bbR6rtBiNZ5p5oA0PaJSLvjhovn/oJEeNPdmm35iliOJGYbDZ
bmLUgvQcNhZH++xDWHzPIoHhxjvt2pOTJFhndiYJp80AxJ3TK1vwmBs3OxrK9wRhPYYhimlvbiQn
piGk/B32MXu2qAdzL0Qbm0OKcz5GjyHOs8JiVH8z+hW+msInJ9GtWBvrjr4LaUEQO636ll37To5U
cDsImB68LeZ9yeLQb0+ImctlNFz4Sf8c+mb6EWGNpfd+E0IChgzNvDsJjGyX2LpBmBbfkKNKfZCg
r/xeV9UAWdATlpzsuRLq22KdM3HvFoWGxREtCzjMywtgIypcP8vFxvEEkBs8N8LTQPOGxCXO84Rv
nxApoUDJQR3GRQNWiWokzM5caEC9rMpAtqCyHCEyIj+tQYcXNanwmkdFcdvXyC8Vltfk0IKWWOJK
zxQH6yrcXwY+16dn/lwI8FhfVn3f9ovSQAk/igpChlBGEnXC+M7zO2iwz/JryKfJQMw37yk1t+pw
jdxsbHneNsvYd6WZS8v3mAMM7SQJixdh1XJtnJ5UtiLAGddeYSAIYidz3S6z4U1R+3PMT+sWGyFL
DoJ1eZKAKUnRbAd73OnWLmkKm1/pflr5/qzmgBXmAVP0XBB0GVjaTccdxHqyl3QWcV40UtSj9v3f
uOPo9JPOVnLUEQvgwMlntKOvl2okOyw9JR57qVXI1TT5SUT19XjW3fYE3q26AgoqIIjiXxqp52UR
pe791zJ1AH8JyS0wJHXzlYwMs+VKPPkjwDj8aaEterckwToIbb66Hxs6flfxI7ikefamWvadQJlB
pMmrvW3YxzZhxhi+RimNOQfqTwTQyxEJx/DYZVK74atCV94Fv5+7Uxv5wwTR6yDUb9uVWp3Ti8R+
6mHkSPkIspuqq/0t2bCannF8YBF+wOd8a8U+Cs+PHJhqZz9cGBf0ErFbSKsABYF/BN/Ma6J93W6Q
KTvGMeKTOw9u1gdy7SvQJQ3wkHYh36V3jJB2dHapePmyqB0PmrUUWmVDqDt5c63GHSoNhGrSCE5n
ySFxRVeWqYExlcbuvZ0/3MVtpFOJoH7H7Lj71bJizcbEVYdxvvtgHxXwH+xG3NFgQ3Zmx9Jteakt
86tk2XfgN4UuypPDmqzIFx2hNFsGQewJGTmWCgext6h1u/hIhCZIMo1jc/S9ujSfArVKQYYkYM70
ZB8qRVMqqJ8pVoy1/6oXBzUxHC1FZNFy/Ey+JJQ7xu7CVqIgfUZ8KDTSqfPo3el2ygVyNlVTSnxZ
e1trIpe3ZkNsswOy9p5TDcLFtupn7KznqNfu3Wn2bpwYgKZnEE8q/PziXmS/KNhboPP6rG1ZWyab
Ip2jvOSKhfwGuO6rWMp56Z8wL9r3QQp4oPNk4l3b1d4U/e7BAYlHrl5lfOmKSZ7XumLEhaDPDljB
3RX/okOnon3GVV5HWWLjkYOLBxiTwDHzOO3Ylx/laECbByFUD66pqzkEJybVBd3SgTYR7B36hpr+
Q43ed13ToCEaxVr83g2JpP+TBdNoJUNNmvjQFTBouNLwfsNrJVa2TPT94yBMN3MbaYfUbLGotzE1
tmqUv4Nh5gXU0OlwbGWg3C/n5cHoK+HPrpaSRem1X4zZ52yYpiFtjNGxZNf4sSg1XsgeWOPvg+fW
AZ03o02GprL1xZoODN7Z5cC+Kp7ZQhqaxL973VIMZ2fDZ3a7ScBfSokdS5LBQVa36VabT1INE/Ze
mqsCr69L7F/leQ5Ob1ckEf6HqTHHfrVxuHYfy5Rgxm+yO2rsyM1rC0KRHZaCJ+9wHItHbunBZgmw
EWBjxXClqxlTtw04HiWMMLxtvpLcQE2PCpRqBIynMwsGPhchw3eoFo3xOAsIO/4hZBbBpSjgerfv
T5M7TSTOYNTlH/N3fBP43cL6Ec2aWxCeS1iJgjmIMyALMSOjE5Rj4E6Ff8PAYhz+ZvE1vTpBLw8k
EOSZV0VVeUaYMCiwST2tdo+7Y0OpmqY/JgtxfInWblaV5RNgLo+mzdbVh0RDsDxyGfRF3zPmSd1T
LxcNnuwGMykEJojRG7fk1EkUY0vYHjs4hZRgeP3h1Oft6aiDZPb2Gv7WTztfFLe6m2aQddGXLArE
WzmByhMjr+A3R+bsoKM4Q+ADtU9qX8+i9IHSVK6JArJwdd8IJelJDrn/49nkjUaxd4smLy/j8VUs
L3I1p24GOpQzwEYf+ohpFfzsoPBz48rzpD442OtYQkKkwF7zpeKQE0CgFSrRVYv86zX1EFktjlaN
y2b3zXN4DdU1EtOg3AbW/Ji0A9+uit6MaSB0JqGAOHVJyVBM+wYG+k+5i5V3LHBGvKPJ7BZG7P6n
rlgjCaSmIya0HdvMI+mQ639+zNqf4T2Cr3IAkDZ0f3GIhErDmvPSyf3ldV1v/Lrs8RWFAyN6CpnK
QOYkI3+/jkRRleQFQiLh4uDCzV5fZqssewgibnls0Twuy5jUMsBL5fIv1FarHQ5aIFWE+nbOoyxk
27OWerVbfxrGLG0W0InsHUR3TQpbegO56Vvt53NYLGguzDiYwXCdRa+eeNIYEvNaYAwOt0k1Js1x
A1f+jTaRoMo16oD4siJQpGFo/sLUq2mzXBQlCX0U3RuyAeC7h3fvCdwcK68QbSrYXFE+JfE3yrfV
a4FNkVSZ5QJH4hHwgMrI4H01LZWS5mFmDqNmTLoX2EJd5zddzB5jpkzAs8eKaTSfDbNRAO5MoqsH
gR49goT4GeshJDAA8rMJm6cfbe8eJZHjUUVpr/0biuwR/DO4zORaVFG8GMEIBz5QTELO5CRjS9iZ
ktOdRqovIkxe7nutj4ms5ZDWgeOTi2q2o6jInViSF5z7/SmT5vHmDjlowJ2B0jKhUSdEWA4X/Ca4
/NZMcs9bLRvhITZPWdemA26mbc7qmGmwUVZsBbfV16RIRnfILaxXEOTp62LJSBgWodw0a6Bma/3G
JR7MllFGSbJwsJFnD/DGLBf0pj3uPpCMUSuc3qkt0HYmhVAIDJmwec7M/cdEWVHGFHJQgEgrJMbR
mwq3Lg7AeS8bzEc/k/cyibiFKHqAZ9PRrL8gdYtuXiNhg5bd/SkN3cSNn/d2bL5jGbXQHDbl+o15
Lccbw5NtVY0OJSVerxsxAWER3as4cH2K2Y7HLhnV0/HzPPU9/QJ/CTMbhemNdtV7hQ1zEokiAaJc
pSwBBmKJsX1kGqzGm6X3lKhyi72nL1IhyrrjxuCP6RlzcdcWdAZxABMTyFrkUsj6KL3iFbHiPMCZ
9X3zx2x3XLeMu5nbc2HilmZnU8r3gw/oU4evP1dgA4uUeGGK65uGvBC5ps8DN8kDcS8QdOnOsJio
X9/VUHNlrLb9bbrlWwsRvnuf8anrVo+jj3Ts2oJ2cYzAA2z3cCqq2qqSwpPSCad+2tMgOiUaoNvT
wREecUSAzR3gbLJb5OXylSQmT4NMVklf1CHJ1jQ3ukItRARYN8caadRy6NiZ2ucCVpckoweoeJ3w
UWS/jOpl4VhV+iIUC6//PIiEydIylieF7jBPEPtCekJcgbf5p4Om8XCcjmRa4lt8fSEQrf+rPhKm
I+RDnoUxNpDg26WaEXV/ktkrjm3RnyPCVUvJryPOKIhnfmZODHT+38oLJlqAy3oBPyP2xXXS5GdH
SW0O0J3IKfQJQJT2VovuOUN1XWoVp/hSoovg4ZTW7R3Jy85GwrDZEeCnFZ3ImLTLpF4SUm0RDQc2
fIpoOswSrMh+x2gEjHpNOQgYVs81ncEvftdo8o03c3fh64iHmBDYe3DmjJWgEVkfpX9gHE0MX6ea
kHp6qp7mPah9HOR+A7+AE2QdPd9G7J7vZcxyaMvRxZ6jASsWYOP0mS+2QYqD0yBr9M4uM2/u6Vp2
MNYKFbAOJjI6i9vMKumAShEn/gJonC+pCpL13AMaO6BMEDW87hOxUsOsuV7M+gnEASuyNoPH2hKU
MGr8Ucwf35VQayGScw33rk1RyKXUIM6gXug/D2E69/0FkE34yvJtqDgSAY3utjRiCpZGLoAs5zmW
tv7LPPCmAN/fqyBQSXLMYu5FhP5kCRmrQkU3WetZQRzyGTdgvutrKeDJ/RpAjP08sk/2FXuAGER6
FQUdKJMw8elndAxwOto69dd8d02WBs29QM5WM1ot8JYQbaA0VgYLpBanH7QTGDfpwTnW6AK2fL8k
HT4PyutCgGJkpgpnpjGEsCaAaoCnzeEgdunLDQXzLyBU13qXSJldVSjCkUJXb3B4o/vGVX93IabZ
i54BSR90GgRGTeDjX2Y+g/TjPoqEi9OwysoL/Vrug5YCAOytJ17cMxC8P2rHuaFwfEt1p/87t1iy
5cBWL+t/nkk8mPZGulkzbAyhlrWYTP9hYLaIoBriS+6Ax+hkFtal4RFbfBbi1lgB/vzYn3L0TfwT
eDsTmFcMDliFupcQcNLJQ9LGcNjQmSH5t0u5nsTgjuaM4G4ZcFYUlhdf3rFeSGEV65/nDu65jKlk
9cJpzbWDNMCau6hCG8g1Tyr2ilAB5AXZaW2hlRcgQB9cW7gMbFbV6HgWbuNfKRiHKyIzSZx1xQfg
PkR4VGucEY80Vm83+9tN7EiJH/1sQzFisZccuFwAlKpSKWrIJaywp6TEq3kbXNyHyO4wnoirRrne
mxo/FjVllsW9Zemo1zNWpDj+k5CG4IqJNfPyXP6qWCRiHrfHoeO/Ws8566SmFIpIWJEyoOpzK6lx
q5ekeipHK/PY/7rIs/wm6qyKR0bYK96ceJOhG12wbDUEoBMoVpM8yhU5Cz085tdBJYc7fp8G9U0O
Cv/503JhBP+SFXphLBPY9OTxBpK2rnBGFM+qcmxDbJnJ7v29qCM5bfRhU1o/wM/tN5YW1Q2a/sJg
2/H3uZGkdROlhHoUIawm6pV51gTOTwgQWpRnnOpBITVZcb1Degho2WZojquVXxalMn4f4LdLrB2s
y/CgBNeIdVKXzSqHjltpAhttH1AA4++iaH2J2Y3eRCP7ngFN/73unHV4CEvzqEeQbMXa+SEPIUGe
4AEjqxw/MwpF6DbxB1C8egnGn1TXEuL+xUYC4hQ6hPqXkWwQZkAFoUDZy8hcgNYH3B4HaaEtRamh
rA6HqEytoYw4Ldj+gmsxqdwzWMov28BaxwN4t8aVimzTY0aL4SblvXXHMyphUjGzIBbPqdPT9s5j
Ns8p3Hs9dvkUXjZCvVavNes14kTBsyPygacaP4GOwoJ0Q+wv/jzhHTN0vvtQyHwYcY/67WiaG5dk
X7RHkWPP+3NuZUWVh/y5bsNuR3LsHVij2yJdIuSdwrbitFhZDmE+s6f7LytpTjEwjdPUzwcVrfzR
7hfsw7ZMaR25F/O9fVhawAz76kv4GX/FBlNzapXNn2dKuEzq6oQ3U+0C/u8S++rTm9mUnlv3B4eF
7Eagmjfcsd8m8w+FWJazNlFeWa7OAdaq3mNNGXSYjXXUXvOioge6fdTfQHnYYw2oCga9S/DGPqYL
vh/iVT3WnnbjkuBViEpa9d/50bPC5ici7HKurJWLNZItSw6TvcGHzJZm8jkJ5H47VUfiE/y/gk7G
eej4H691AibYdA+Fe2hR0szTV9dg0/TTmvxtYTAVzk5bvKBSoisuxq+wT+3t2DSIJ9XK6gDVY+V0
a+BZEnfJsc1SrOKjcM5xe4n1nmUG3PTDHdllHE92GJncXkREkImbc7LsyFcTR+feiXCWuP5faeXt
MP348qBno9PJviTbywVGXRtNrwsrQwSb9WTtyEbpLYQVYNdylmN9TQf5Q+h/RW7UfDFrNZrFilsn
SvLhC5J5UZTh1SCawQGvByDfuUJXhTa/Kahp6fmlBLei50w2x9rB/ZxDCEJ+viNWIu+3K+hqI9k1
C6Hp4cRCjMhDRRYyp7/x18BSJi9WxhZgK33qZb5cXdY3LS0TMwzs5C68RC7SGcOmdUH92QcoCL5H
OT2e13SlJoZlCqGI+Z4yraVzx20iFgv/6U4y+SgQvo//RykUuQrb49rVap2JC/Tqluo/aAMMiHue
SVeOJnT8rT+QR1dsKN58xdukjNp/1vDEMYZuSOfMW4KE7zUmIfTeIu9T9mrRxPvJNTYRmBlvQt0D
dDqGqur8322zbobadzab3SJqisUC+/ZqaVSdf7nGuwKDL+293A1NWTe9qTjzPsOY37BCy0EGrbbH
bfpnj3Cwuig8BlPriimt24rU/eUE2WdwAYvCz0HEFAD2m4xkV4lKksPyRSprNCywXQeP89Agzl5o
2Qz5RYAihGmMC1DfzIdw58L1S3TkhDkAhkBhYs68rFPGnoFXjdHXONChNOsiq/UPAtxaP7BclrUA
Phw+e6PJdy2BqnHI5VEPpjTI5mFa1vkRgvi3QfRyR5zQSfuK7ttAye8Xc/nwSo/U0XmyvDI8uVVa
kQV7p9pbFqsFfH2kEeEAvTLJErN6rmFbP9Z4dFmUvXt+JAJ8YTeMcojDEb9XlinJC4G01DeCsur8
qr6DwIDPyr0ofVNJwANUib0SQ6TwGcO2a256YJwh2nIjB6AzagtWnHJxCRG32kLI/mLzIS3RPuW6
cWEdQQvcjg3p/EUHSWI66EYonZIQhWremo/ljgmlBPY0sMYA/KFCn8+MhFEu2SUk2fr41Pq5qVXM
dSJ1oc/aOmmpSkYCLOW9LNfKT4bGHUS4XAy7HWTlMMZDer5if291xa5Rj3+DBaFv1qikwJ5LbFQ4
b7a3+1sYw6gpc3qMdSn0Orsj7xGTU2yTxAGa9MsUW7gAeL4aQzXZJosvCUN6rSXUO8d866Qi22jW
+qXgEPqKlm7KuwKIGmKgc9PpLKpLUHn0dGTd2lPdZsx7LN/I2lzGnzmYKZQKwuLyRn7JryE/On85
eptNImuq/W/KZysFFaWYg6zmxU4vEGXEdIC2TRTc3nhdd7FEFYo9Axbxnq8/Y+Gs1+Fr4HdElSjG
3eT+mVeE+FUOo2EaEEalrI/XX1JLAjwaVS9eQTuU23OnRhvaZ+yQLhkhfC7OHWWL+dSFBHm+mMTb
A1VgoDpmQRWxQ2sbCBo0gIAL/LifIWijf1Lv5q7PHs7PIO5hMD9NyKVIE4DAlNgi9YoV4CcznKCm
1Xx57GDMelrrDbBTfmVjcSFlUJU/GRPHvvfD3/L0cTHc+5/XTfFmcWWzxtz8ZupHjeVKbHMHk1mZ
Dqwe0d2Glq0GQgraBl01rfbXnjRpVXhodc1MKPZIxmglicE5TXnqCm5RwYna6i8Xtw+PWy8Umd0C
El+VhSKoVMcgNQQs5LCjkVCFbYaPXATlzn4RkKViTqlaIuMvB3oLhPl7ca7ccvod4W7n9cwxmOpC
9Z8Q00EBJ715MDORvU3g8XjtmY4x5SRHfNkzLecNe+lpDA7IQ6yoSI29w5t1en8zmkAZVEceLW6L
aodmHF1cSutzTTAD/mXUiODwaj7aZB5Ptxo72s0fKyU4FfgTc7GAVaLmahcXtuIqtTnff3UAIBmi
9g0cUXfLCPFhC+E9AZk6Y4AoTL6N+yPkTjJS16Ol7dTrcoddumzmr14FyL6X/KXrJs6WFKLdB/Gx
xIkrfXhBPg/inlxcrNxszDd6qddHGaPU7mlyTn0lV55L9e22mRz0Z9hpS9zu5GGZYyrPjsvxhgQz
Z2yoISSQqgfL3uYirJpr5wIl7Il6cUymWgky2jkA3HXCr0bdxk/Kai2rtlAmO8YnU0hxIttUBjIM
DPo81Ix7RwrnIEe6vfidTI85wV/c1Xqu09pcrL4UtKp8CzlvcNZGLn53XpRIzOnbQrcs+78ixaWq
k5oRR+/zJikyrX0KJRsMV/+ISEINThbfsHdg/+cwkvt4cQ1IE0kVZ01zGSmDWSmsZ6irnGxnLDYb
JWj7nt7lbumJFBvHjlIA4NKwN9qpYaXl1Akbj0PkgVu+oD7121FGtAi5VPJkh0ni0sDuTMgFi3HO
IIf4cRKYYvE7TqCUb5yV7VQLzgXUujW55V9HJgMpMrB663kTZtnvUpC0FLDaJOXoTYqQNKay/OcT
R2jfBcZYXGVpgAIOflyIx29VfCUVkbX5QAVdv9DD0hbIAK4Z3qrodCzSlZm2XBSjUKr7p6nzoum1
pZob+6s8946SWZ1kFNWIXNIqfAADtNTHefnRE02yQ4SMd/i6c6UaG6zqYY0PuodMMP+OjSZuvCQp
VAvcz9TZNU1tatG2HTaQDI94Mjdc7fWTaCC3o89c8xe72kBF5EVoGj6iNFdK0aKXsaaKK5OHHa9l
yGgFf663/PsJvGiKMNMIX4sasv/f9EKZzbSZaRsMGE04yWgNWCF1rrxSW4O7UjYg7qXs6TEWZXo6
eohR+txOrpSx9AZ7SbsTB8XVEqlI4Rpivj43OfiZ7/E6kt45+KbuyWM8M0UX4BcIPa20Ap/W3ZJn
JAfzNXbNrD2Hg18IdzEy63Zl6qaluNqV5T73P285m4Jo1vtshYUI1ACx5nEC6y9uRPcSh208nhGg
7ZkCw6tBbLIVtoMwjVAez1eoIS4ItxD0MYATaBrjpaebiZIoTRkxPBSau1K2Gq3Vv5yZ4WKzUo28
QfXLGCMuxwEjN8R/Tnku6QA/bQNIo5pBBbdfaVlCzYx8U1UGXT3PQIG926828VxFA25ykLL9ZOMu
G+hKV0mv9v6/utcAg0If/mk0sitcIV4QtMLt7wII7hMoz4zcta+Drucc3BQlSNIIflZMx3gKxsiy
cYJDO/vjdJfXE99eIkaSY5G2XvQ4Z4kqcUJdv59mp4J+EnC9dtAvJYpPrj+AnQqHfaiKHfIFo3CZ
movEqoquJS/Z1X5NeIh9S6z/UnSacyzqEW/RUWvznZsLMtOdJup49BePWdvjgUT/dbDm/JGiN8FY
sF4hPGehvn9SS4dUMcQTIsZOV8XiSvsB5gSlzsvFIBCMe9eowW/IByHEMfR8UHak3v/Cbsg/Gu8m
qZjYXyN0rLl8aMmEfiwQ6XbKe2QmbZzDFUVxfAIrDnb6xq8wtxHEyKBwM6D9URJrXWgpfqrPhGI1
ydWE0vCQxqqOEoBmHqx53IpqNLhAzatKXx/zJykS9ufhNt71fPsSBmAio1F9bYjoYf8YUY9WQgr2
8wCmB9mneldHgW6s79PA+kvT8ZqVv+06GD+oihYOPoH7CK0q2L7rQ7jhAwiD5Srk30cEpVdraf4b
XAKiAKv+TCommVGoDdYY+Ty90hV0F5jqvsQMAl2F18D5zxHMYCWHrf8ROkFbGyFlX38Bh9BrHDgU
Eo9NysaYu30IS7X27fDfGkT+owFujqDF+yfOar5gGhJbXlUROvGjUAZuFXWlepV4VyF9ujWhWmFV
LjncAv+dxaWJQtMFP1djjNOb8/wGSWm2SzI+sbs8jZnZGBm/PfgVvUMYOI9N3JBMOStBrHeAdrJt
RsmrHQFgTnPVb2Dsa5rmEpy/1VOyPr0lSRyHHW1BgLcHN/d7lFzaOJiOgIzKNon9wG30G0p4aNTi
sMcCGf4hWkLX4vX+VvCMb6iuhPKApg3InyT4+o1k4JjUZvjc+gwU7t7x0ZKTS6UEJFEtBeS/a/b1
MLZXxQ9QHNWNdytKttDV0GtisRGlNh3fVjvNVKjEDxbvLXaewxjDkd5+cZmBGCX8QmBHGbibbidN
uOY7g4gxG0d9Vz08U0NvH2UUtGjzd6ybxZhNsgDiM4i3EwRYxqtK0kozRiZz0gAkGvHPyR9+wyNO
bKapS9Q07zp7o2ApyjtIxMUdHm7w1pLF/2qCdWiKDWCZlgS0Oe80OjBIizFg1X/Ppq3GawwvE4of
jVpG76GmoofW6pY006yY51be31Gdg8Pb8hFfNGcL7vK6QfBELyxBiOSXZnNZduY9sJ53O3Lw8dZy
DNNMdP0912nq6qtBhpdX2WoTs+YxY9JQbs5GDcNy4QYjC1rYedCGeBj75zn1RcfStsxu1ALQPquP
rx+M1Jk/7WsSHGARKYXdkSrOZeYgnBBaqLUm6lTsdT4H1MRW2oWS2aP4+ATKHLSV77c+TlelUuo4
WnDwW/OszvYACqBkURGxXB6po7ZV5P5IyVCTUmem2N0jnHrK7zHNtbtkftOReXE87bgPWRMUye71
JLX15GDjxcHgbM9QwkvWvbh3NEulCIRLlscPJDzr6zpBEMlxxkWJIIqc/ChxlDQKPiABSsYLbGCK
ufuL5u7W8In0ZOJ2qBHBVx/cdEbm1dVLGup1wcJ7cgVzdFrBXB+3yQMk+7/GrRn0S7kIbcPZA6kg
nks8vpWzqK7/v+4gcjvLr3/BXbinvs8JoP4/ytpXPvc4GLXDl7ao2f0TRvtrnZfO6F4pN3Xc1EVs
lRmKFrquyL43QbaJRsPIagHBHSeZzWxOgcMHVazxqvGeIBlhokMqSQOIQj3Km3VK58iESGqiIbjj
XX1AAIfrQDjIIrb+hHnrbb3aXf3aCmPEAt7OqhYgGQM5VS6m6qrzTnO8aWrgrvgNQ4svp6uWGUZO
b4/ZsjxfzLvb3oQmXgXnTxVzKpwDd63QpHUFlcYx2s4aaQ9XfdLOv5nMN4EbK6/kQiZLrqG1qcwf
eltHo7Nu61KpIKaSw5lxJ1UFvrZN/cGBkfTbF9KxwtWAsf4knvOaIjxC+tP6ALItOmxGMtZwz0fd
zT3Ki8v9LY4GUKEedIRg0ZNd2CJpk4uaMsWCmiNfw+Otl2/cizPlela5te52mUBeP1UvX7pfSscn
P8GNG5Cd1L10t9V2h7bnK+3C3CTHjuNF/U6038XegwD7QKWIUQXONGCCOqxPCVaLt7IrAmz7PRFF
gXby99tFNH6kXTTBwX8FdS9C2e/nCEAAlnaS82EmI8AlcCcGE5M7pqzTfrpq/CszNn60sgWZHzY9
FssDeX2+Ss20rGnbGoim325tlc3ewu339WMRe2c4IJHzb5iKn8rMcBC9ubEtRGDbuBPx36o0/KY4
2vIlckJd32Z2piAlk7l5AuQMbIZr4tKq+RhMqTdJ6griMMMCLVBH9TjcrqddvNt22qJy+3t09k6E
RaSRRTGPgRp2q0V0YauUsrNPbpPHqyUHMZSsP/HO8hrtVrw8ZN2JhGxQGrhaZn3dgQVVrmA0yfeU
DL9T8U9eeZ6Nt8IVi6UmobMH3NqflCXuOiXn7sbBN5r5zblve+874LDsNh+YCyLSUKfKYvnokmeA
weoJaQJG+lj+c9tTAntr8zERw7aD5QVDMCHrbtYgr7Rv2DKKjtz9xlqGY/I/kqzcfjAZr9iRtWJh
jUUBRjlQDgyyntVGsvui4o7WpMf/5kFkeC+2B3uVDZDhnjkVS8qseo3aC55qTRrt/xi2m0WrVsoO
EFJFATrKxXFJMCKRVOT806NjcdonvhgakVO3/Gn4OFPzFLk9RT1xrzlMxWOzDPHTzfWKhIO+CTs2
oGqP5i+jCjW894eB4UuteZyNbVIFnurAPZgBXn7OkUEujG4WAx3s2S2+zbww+Ew4CoL9GmFhs2sX
XV2CbfoFsr8JHanh+MeNlYw6vxSxKQQAhjFSxAeFko9MMR0UTQheEna+oRyWvTwHz2N94OZvYBMy
6mDibYAM96hmmu6xddHzN/+y3ionX/9msc3SKodK0+CCcGBjKE6jqHE2vx2df/hfN2nyXne1xEeH
t93/EMD1naEK5EySQg1fdAFVHxwX91VDYoYGAJBy+JSWiD+VSM583hOKs++2vdSNyHZFdQq2bFM9
yOv50zX1UUVmBVyHIpRDrY6LBwyVUfVNsSUu34l5IN7n5VDliLxtQBoRWWzVOx77iXOyP6qY5Qjy
GhTpp6wBdTPpjpxD3O7VLfhVyj2ZMZEpU67X2NeQj/cnBYEA0OzVD29RQd/PYhkitcnwI1c8DCP0
pOpzSGsUthL/k4TdCBVVMM3hXkuBpyMDzhtieR8CIFRlO1NOKOIYcKAxCFp4TG5T9YS8rkJSamvV
rOLwu+uR7wdEBDlvudCnyyAmVSYoqqGwKR2f9dXLNAS3nYrarMVSQvXOjmSuK1WXCwN6H0u4ckqq
M0yiJeGpCRLe9U5bZIbHfW6OyinX9pcS2GnkfcTiNBh316Lv5JwJftNHDpEwGvUuiQtStVS5u/Jo
roJV+VKR3BAn8QOGCNtqJjCx+uOWC/FYejHlL4j3FWi+uRPKgGp2iME0EgSIxheIUiIN7kN9MlgZ
d9ATHIy4JR5lYQPnAGeb8Cxu22blGDzz01UFyJ/LiIfZKL9aMI/71Tx9lJEWBDxSLx08DRV4bG8z
GrhKxz6mhR9P76TAbPOfz1grBZnCfxmbhUt1oOYvVFhD1IL7RavynfOogpJCZln6jLEkSNr1D5s7
K6vk4S0RNfFrsVZ3GNimnDHw3DkJkT18xRXAxYhYXH1eGHWzUhruM+GhqzZzdl9vjpdJrrykTXSQ
rRAsUGhZDFkYAyrDPGHrbNpoA7UjOqIXb9Gwz1HS2N/9LfAN0RUbKVnuieo8cHsULZKQudnz0wa7
T6svb0XJkym/UWPuiY2tUeAJN28ysRrLxrx5YZoS+sKEUcfPD4KJNm98dluDqZHqRbNf8psFg81J
8ZU2ZCWLtZc001AtgDQm6/lKU1O0EnIdrkha6eayBUkzc7uIeh3W3BtD+Hrm4LsYaFl+oUZfonmE
cQp3QZ9NuMqJcyyVFAh8exXUB6t/GOnZFtwCkv4zkxYStwRm7zIpDPRFdA1E7GEslyO21wtDj56Z
gVAocz2bA1pt3Wh0IxOmv/ncEaYElQly95c6TjtCZk4MSYsCP2szN8k/KUunISv44ZN6FdC4wdS3
qFCuxJGegVn15ii8dUMriqEXAIk5b/AKVIBbMhBu1/JGJPH1pQ/twaZTDoctV1W5XJ6FjuX+MlA6
BEwiX6ORGla0zVrvS0VXs4c2Cl2LAuIlln2a/3ZCMQICT402o9RPr1jwLMd+wJymV55j/DGzH9wo
9AfAfVhsCOLbUhQ8ifr8Y6CSZHjkFk/zQ4vIlEN7nn4DwF4K/xKm0rVZAOdA4fu5Ubuf5Y7asRci
IRxYNttW4si6wIpQZCLM4Fu4gRr1aPfuS/CdQwrKcjrrEJs6sSTOsKHwDcsuCPJH8metqWg5IytB
7zveDD+ghJw5FuFDaCfgOnEFFJcIKyiyIi4sX+Lxxh6OOlpoR/G6GlWzO74l0f8jSNo8mHoa81H6
T3aCaDVeDOaqM7PZ6FH5BuMZg/4HAt8DApKqbX7Vx2k9Iyn81Q/ZbbnCasmGwM3KSLA5fKbZjzcz
vSQdtiRtaKAl6pjDiuDOHPLkn1lYmzdjOV8UL1d7+gLUPPWduq+fLMN/y88bjICng5vvG6fFG4WV
AZ1xNo7yMPaJLWN8+RUnlR8nl5OnPVr3NOtdmoX77y6iSmbXeQTor+fyhryj3DJYcJyAmZvsbgMY
F3u/7XEtYT8QXp852zotUR6izW/SFKhvNwrQnM+f51zt4huJ31VSjk31vXbrJ8cW7BE7XbBFxhA7
AeroUI/89/GIK0qfSsYLubekaOC0LGEvJbyJiz0dJKp9L6KwXVdeoa15IuOJqlr8s32kXf+3qDyG
cu7tJWUlgFyxWnGqa7o9Wg/vsV4Cj7DVqx0GqKdaDVZIjGPMYDl4lUlvvcce7sFxBCrhFim9CZda
ZGDzqai4hQ8Br4kQRwOYNfIH0PJBlbPXwk9tfScTvUmy/3iQKWosM4E24aLK+gpCbMRLVtijTxR9
rQU3c6+527asUpaDY2S1TIfnAYk6Q7gitQNKvurpec9BqnABkkrX0kZM+nu3Z3G7/W9nJxfMwESv
O0cyFucfxSxF8n+m/3dCb05Mx0qrQSvZsXQ8RFzR1NvIlnnRcntuHWDXDClIdYYFBFlmlWp4yaAa
yHCtKV2/3S8NnVr8YwRbBeHnFGmpEO85sRjjYp1xeoiFLqx07yMCl/rf0sSudeAojhyaWL1YKnP0
RFwU/3efsqqaUSD57Jr02AH3B6ACOBtkvL7rlEatjgneF5iuBpSec2ihRAG3TBgcevbgMhEyZUIZ
IdBJXxkqbH7Y8hZW9cjDW4N+Sy5RXmGvdODLbcFp7n/vQYME8urOHky+l++YPKfee7OE6Lxy8yB+
gVq42xG90ZLEBYV5eHlg5v6oNQNv0sXT0o37wwjZE3h3zcWpX/GO3jJ8cjdWqd2fo63B+cRTbl/M
6Za29zA/9mb595Gv4QLTlVGxzRXO3Lc9PBqBKANgqCHWap18q3SV3BzJBonRhRw8+zjVQSVx0RkR
yHjqqZmfjoI0zp70ph3Ih1RNyzzYhmJiuutKQHdxXCZ3GTegB15jugrXWi9M/OryrtgsHt5BkW5l
qBeM6R2iDJ1D8M8G3AZMsI1gIvBO3Dg0SOhQPgD7fwZ4t7bPZASWFw59i8GRV3bHtaMUtdwyx/Uc
kFSs6iRXQYB5PY/G3aYBRvwX1v/3BoaDgzGY5qEsMcbbGCvRgIlmbUuPMQEMvrplfzjCq8VtgoFq
UeEmEaT7NYMtoX0KiNjCXwvBA28dyN46Umffup0GyjqE+UcW5dR6QoVei6Ik5Bt5MvBXINS02VN8
J8kPiUsfrxOlkeQAe3gAv4wtIws7VfulKxrjqq4ybJqwkoy5+chLObKjsbS7Hv4DD2qCejQUuHGZ
ki09NUSk5/ytKB8EOLfhL41m48Dxyi5Sl40fP1QAgf5hU7xbFdoreb1L3gMqMoPLwuXRY245Tm52
W4XLq/TJc/A/SsOhnfIlvkRNKlWq9SewxoLRkEso+SO7HJU/wvvpaunrMsYtaH2ZiJFNvFSSTD1L
471xzOeRgBgtDhwMkQr3GZ7MGWeu+Mg6E/DbB3J75opZ3H59CpkVLvNpEV54Pq7ePfu6dL5UpIMS
SZlYCrAYYTjXPf1zxfoZYkp2l4fQV3RP/vDB1zIri//t3Yi2SHwfuUTshq3UQ2DHaKAJ+i8YUBif
1NdzbeNFhMKEWXfwrOEiPDsVi5tqDEpAql0gUY6CvfFdbEQpWpdGpgADV2k6y06TnvyXNMp6OwTb
eyLPgXtv1h/LyvIsoXZCeGahT8S+ShoAFPXYZ3XC64alrWCf0AOQ7k5QQJhEJA6NrtUnVKtZA6/R
IsxesSby3xchR3Lr0QT7P6/Qw1L4tkThqYRvUgphGT+miH3gXQcKVnYsUewPmNkXh4MZrybKUOnJ
tVk/ES3BHcZd3dsiORxVe69zFUmdtoYXQNx5EFPdSvFI9Y8H0/jIy5iPtlbz4obH5P5QV1d8XSTz
3b9IYOmJP278ChgmhDK6uq+LYWpni0/yy9PvNRcZnFt6j5yq2iUhSaiui5W+zMEe1beAORC5wxOb
pTAERn+IJi3AWVZ/+YI2eqxZwZhXSOisdC00OXQgNr1zY/TVmPovNho497nGV1gIPcghnQ17H3tc
iPWS+qb+/xqnEnGEBrpLSDm3txaXtzIonvNtbV417Vb6akA7CzPnmVydb8QaSHwFMw3BPSjIu+SJ
Z5hzJfsb9aMyszrQYLAm8Z6P1nS6WH665RCh7Yod5OwGgfAZI5xLjQg80vwrjtJgK4asYGabkxbD
Uk7jRAICliUSuPj4R+Gg3KvoOOjB6Vy+7Q5hdF4/2vXqRQgglwlynEzzu+OWUokoJjT5u0hIB2Dc
TGWxcChJDP+iExGfgq+C0ENDwmRxbosDN3uwsjZo45mbC1urolQ9f2T6pi7600sI9U2iMDnwpSJW
Lh1+36967/R7Qn30iGlwqR6YTDCAz+V4s56vtR8Dy+wY4GSrsisuCzsufTeM7KpF07DyfVty4RSE
l75yueRyVv903KcPmRNXTG4YYC8m4D+15vKEf4y0r9/c8phGu4Cnp9HaudekbEJz8t2eBV2dKj5L
JKbXufmxPEKGKM9urR1huWycqN/TSH0XqJIgtMSOGxtfh4hLBuFrp6DKJ/DZuelrxF4mMsfF0hEf
u3h80JzxX5GwwRVn96SbPlzloz73Wc5kliAQEp6TTlFI8NJEnf+k/2D5qFbHOCUcnQSXLPqhh9jk
MLJo9kQKC1EruqqtEbeYVv95TlkgfSeXIZVTJlHty8bie/VVYnU/hOx+BXmSLxsq507zzEMARP6f
Jk3ZWTArGNqSlJfgOMV/BrCtqL6g7GzHWaoZ+yPVeBMQ8FvsUfFYvjb8TC0S7EawGFeAd4imcmth
9X9+wyAhq24E4YxDIZtwHnKO6Rh3Bl+bi+012+j7AM/joz313Ui/I3gRYr9x791l/7ULbWGLaIxf
XRE08W8T3XM/HXsFH1MvRQWOp4Kf/2KiVyJnoVsJGrZC0Zw7NL11eGM3RaOe6EbFAnvnP4B9vm4E
I6u/JH8UFfHNV6QqVoCp2YXzhk9KdEYvOHeVIx+SIQNvA4Paxv9jk3trsl40kgbRan5WN0JJJx1E
VMXsPEujcsPJWfLoR4NW+WUXVW5Vy3BDXG47k6rrlLnDDJQviwld1TxTNf8a+lVkHtyr6DlfT5rd
vE0nD2HdTa+9240AUgK7i0deoFx/mTNNm1OUGXujO1Ycw31Ifuw0h+7o2VaLSMPKeg/trqNiPt+U
WtBhtss37yuqvwNiO/wf8+aNabk83Th15qc8SQutdhwv0UnU7+KkAXhYdT+E691w/9zTiSYOlbqp
m5rnWCssnB+xi0Lc7Q2R4yGRerdUqaWPaVUChQZ591yPfy1HhwYvSdkV/JbdHs48TG4iHsGj6dBO
ldd6yzy6BbRqFr6LaaXVXHWGFat5gmDvQTVJDJFGPMiMlSwToLvEJfGkvtUic2qo76FkLYUoA691
O3CQnNrhaI4VDkjp7okL09y0xnUt1Ul7l0DpS6z0rv2Nq//qepfO1eUjus4MO1AaQ+Kf1e9R4IN6
7ryTJIWqiOtiBpiRmbB+d5I5c/XQGx52UcF2EKOglbygZy/I4i+Fk1IeH+TrXrRU78Zrl2okiiIS
QWaCQT1irXgztrCtM1EvNbIrHJdHtD0Ut32ZaN7U2UfDUtiUV4jfkLRpM+djch2xsGNoRqweL2Zh
dBtH5DQ6mJPxrUQVogffqu+SeB7xbgamsEQxgRogQkR/nfWUc7jwMQYH+Qtuhuxgl3JsOZAZoOl/
ygfX++gX4v8ouh+4qpxijPvz6mkbGE9zJx6iv1G2JMSPZrmsSU75ag07VeboAqrwOrQH/5zTL3b1
whgavxspkr2hF5yTEs6a51ursJzZwdouA6B7Zpm6z7/sefXj0ZAGj7LoozhnOymQ/btgQ9/2qUUK
p0/1PgjO231QO2fAMP+nN/yOZSwR59v8zvN/gbXhgb0+4JG2Fr4CzS9awqhd83a82nNUnevRxEpz
MAyGtej9kkeA4ZR2ewZgj5Eeo+45b+sb3u0r9/BGp8n0Qhfozf6lF5tzbkqKLS0CTzlZ4leqeY6Q
1TLmwSYMkCo8S263OpUE7+3Yr+57KrdIDsAGNrowP4dPcQfpovO2X9kLVGeWQVpJgsn0TvA24GfV
IR/L9cKI84NSUBOH0i7FgdyKIbzz+aWw6L8xp/6xqnaqvm4vKrlG3rxptEa3O0Kd+0Q91F1ct+uh
8I1xSnNc7rqVzAY5jaTBg3VK5XcjsAhE1BYKsdhbMAyxWOPEE6ni9E7fm72lTYOUHqqeWDE6y9gd
hip/EHsIq/fTR9sI1Jpmb905nIUxYpOknKswJzWDZJ0aZxgDUroxYKP9UjoLgeHkWtnsHbmgKdP+
ji735CBUC8fultErZbmR/HpxQB94vu7fh535lZRW9ukX7oRPhIfdpdH+6HLKTNWo4OUUfFxosZwZ
Zj9p6jCKHZtYRpPqoEWK5WecSZBWD13Fogtt0PpVdnmgAb11QfgC6/fS2qpPFswWcnM7aPD7CTK+
bK64WQffBXCH8DjKdjEqY7s33pjrC9QGNFRpSIbpZWzyJSal72VU4dCPKUigBgxSAoCO/8TOnXjN
s/Sez23l9CsxCYkug8VLj+6Wb1IUldJmARSEYz7W+Z5cCOYtuKPVIrLOGaGqM0+Sq2C9U6GSlOiD
z2xv1Yup4Tn8W8WGJR/Ek+jYlXMkFP48M7aCW9BCJ5NkXFnREABFPdaD/RRCGHwobVEwNwfaItj/
/yWMWWBrjDsG0RFhj0oC8qztak8dS4NUxWna3KTC71QtvHOKJIyDSCsIdqa2xS9EAPFDM6nT9kjQ
5lMTxAc8ZasEFf/qyzd6OmuzVqqWdbD9++gf0nmzvGZ4OIFrCyIKEOJeEwNKMRdX8I9EsIGZqjTn
I+tz3LKUcwV/7C2DY58Zk5PXIVetRWMIHp7yCEIgjs9K9tuU87Jd3cioyIwgPl62eCp2gswhO5Gq
Gl1PmWVax84EtqXLuxubrwJJ/0aosiOIEydWeNXARtxZXzav22JI1TmnIzM95HOtcUqqXzvEiw4W
pSiM92OyBy8vFJp2kXHqXSD2lwGniUf9dejgbWYaKAa6Z0/Tr3G6NQbFtL6omTK6vXTLIIxHr2tW
su0IPir05h5dTIkORnk8KwoP7n1Z+0wS4tVVc7KaAFiHtBfGNnCrxNwvo9CufTkcHsD9+K2QQVrO
xzoFT+2jYdtJVi2PxW/LkoZfUHJ5/GeaaYP4AMmylHTwQmUEXMh61putddyK3DcqoMvUdlt6clHH
O2JNtIrXa2iHXKQuYipXA+fbZZjqCmeZPuI5pEaTXKTYEqMZnXrzdffpQ4/2s1b2r1Q+VjjKnelC
Yrqn4JB8g/TAtiKok1ivvBYsORnaMML1nwSVC4NeVc0UrGNLMyggYjp6h1m04uHQI4qxzmB1H0fI
JFw07004eR3rEftiUqKFJLfnadeMqbweTZC87JSYHLu5bBnYWn/S/MpKvhxj3EZuBF424ltcFnNi
x2SuULPiWX42UFcj6l9nLfhNQaZhEnxz+OkR/CzDQAvwst4GSmwfoVHmkR7d7s6x9Ek8TtDFKLLj
bH+aF+EK/w6OWYY627MIRvDCj0i/cVfiN7XRXcFbj64Lq/AQEGe4mbADddMYjgyB8zKn8FBxJoQb
NQS/Tt50N0ZcosuY7qq856KXP5Gmj/gZnMf1B6RTX7MaNUY5nF3bci1eLcZstADdzisk9TrdfpwP
KdB71DlUdWwrfEL+S/u+V/iq1pWPuuaHqv3ACnBFoXPwFvhhrapt3r9J2hfNzxY2ddUkakiGrFac
K8JPhQAu0bU62PS34EdkpSZX2ZdCVcf960NgDLo/y0fQ0thv079RngNX68QKFcBP7S4yLmnIEY0w
qOKyJsqn13zrL548DLzjo3oGEqwmPhNwL37j/IrXgRQjt0FfBljrAemx7uIs5v8E3rhINBKjWT4c
a1Lp55Hvya5IKAcVsKxFIujeIkFExlfr6PJcR7oyqDpEiTkRKXbZD0oXuzvoKNh1LBT+v2v1cZtp
o+YWOUc/m/b+jNwvTpTaeDN5aEYm9im5TLhtZ4hdgr48amYTYP6J+c8sGmRW8xdu46HJOm5dnvIt
7p6lMzSDiDNS99B/p9OG7gmFFR1mavZ+L8+AxPPp9Vow8EvvIV3SUY5AA/Xqw+7nDCAtypmBWNg1
P0iwUcTyS5dKQxi9vvt/He3ZYT0qTdzTFk+NbkaVUPjVAkjOsSiCGwoRESOIF5NcP7l1AahX1sKl
dp2mx37xQ9Gj2prURErlGS1LmKswYYYVvkOP+hpSFlaH9AGhtFPl0QuNVBvjF0vLKaXH99tM1nyY
22vdIFfEykifA+s46VB/bD+0whzxtZ7bhB+MXe412VeUgLkEDRoEIM+7EA8Gu38qyfZYMEUNnHfE
no5aPjsNKrDakM6E8Dwa6ylGfwdK213UcKgIl11zVCVdK6EA5+UcyPWU3ItRAlNWQOb/2hZyS7IX
yQIs/R9kQzwVlES7r82QqNQXtepwSiu+5YldYCl8CILgTRFDR+RN7E1oylMsvrH0ACc9cLj35Jsx
AXFxU8lSWpnlcA04M0uG1hqcuK1+pCU3Y9gWdf5mm7OOFatUaSfH+m0A1Dgf7afBHpnJ9SX4fuXI
EU2GxQEzlW4fTcKjo5rVOQYqWzktaaGm1ZmeyLix4llUfMaQNsMxm768U2vrzTRTN0rILGXPoyIz
dTWqyQs54AwRprhYik6IEZT6KhA9k0JJcZg23t+OqoMU0qPSsFpyGmNBRQatrTcccHd4iWpm3u7t
cjOba2qZ9WqjSzOUILQ4lut7sE0NnKBW86C0hQF/KI7w3mx5jXrgVsDT0JlyTeBt/AmchNX8IOYl
x7bRCTLZxkQrBvy8aJ5c2KjAQvYzHMgCsh8Yg3sPnwyHNaRsuuMWwHRFlR37QBkDHBE2+D2kb9lX
Ol4j3a2EyZVRQ1sKgow09PqBOx3qxRSBKVwvAeSMxyhOzV1KDOGs8ozDskL6DHM3oSDSe3w8rgKP
6SaujQ3MYF+/PuNQ+vyOIXQzW7Xa04OvkGSlxfcGCP8+91auqDNJLFJdMm5JH5JJREwhqcCo1A+j
g4Lt3LaLC3Xhjob5PR0Hz04uAorF2243/OFV3i+8G3otKZbOtibfkkFrk48CUJTUWW9S5apL1OUu
sHjUoHYR952tPaJJwlzN/AsUMKkPKUPaa/6JxpIB3NKHjcz5arc/jDS/3WMyDknQcbOg1PCpvboI
eF1IXdvIvtRKW2tt1+j4TqBgRLFt5YXcP41JH9nZKngFYagt27M23p/d3ZB9p0WKmujtlBjfzt40
bQ00yJoQxSbfJZyvqtP8dpeWHU8yJGrYDqvVD+cWkWHbW2IokMLLo6+J6LilTNANxLaSHEhFFCdS
+6iJ9ctEywq9ktzsb/O+ThL+SImnhRtO6Wls/WewJfBIJQwIvrOtMSUsvvJkzdfr/2Rbe6DA72HZ
u7os4PwpFJrxk5/C/SGbg7OxDHxETF1rx1Hb2s9/TaFtBgfwNvS7DRQNvGQEi2rMkkuvpFlYB71x
SXpXZfWii7IMNJsoRSg2xtvR1i8sGPH40jutdCMVGJeRxNK1ffJlg28OlMwDxZb9BTzi27HaKC4t
B9TbgEfkec82bV6sYRfiKI6YN/fbrnQQSRYO+kfQ7t6RV0iJhAMS/f3uC69BjuTqt5VmnXPy2Lz1
oQqjzsGHo2XoHzHTzhnUnPXzruuFrERnAr5keurLYpYnS3lZZ5mq7Vf4E7AR8wgDhpqsCZgnBSoe
IrMqFMkHS+cgdItn8MBZBqMaQdaZJWZn/LfwQqj5R5lqozeYmYyDgdTZRjnveQmOfulFItxlmq2k
Xn/ggv29Jg6kONbpyHDkPVldVz0DHsxLy0gKklYuxZRMqluc01ytA7j3nf17uf6KiVWgUWcaiR7e
bPT0IGjuCHXjrp2fQJ1tpJbaVsH1rw/gvOXQEImGr1/mpVfoiuOeQ4ceQwvRAs66SURoAF79N9/A
1CnXnL3s6bhNYFj+NPWct/n0H2AEedprPeb43mvAYZbq/ocQfGKVCGKUsgN+N9LVqlm0HO6F9P+I
95RbB3SMB3nf0+dczrWjhWO8FLl2G1jyiS0ZqcV3d2uMJffCMLPrgszrKFYkmjLhD3hGqltx2en7
lZ2JCn5aKvOfQ5Qk/va0j+f3qLe2Ryng4+k89Iu/bY7DLmi85RIyHN3qyoghgYKF20s5PIEZlD3w
t99KI9oV96vL4m7mJxsJQjPS5HRq3o8YtZak5kaR98lSuhAwuHKpACsrOjX6OmxTAAdOylXl6BSx
/t5TDmhMtXpU+oeLlArajZvOB/RsgWBaHNp2/kdz/XldyIjKwInKTCcvPFI8yMr6cJ6WQ2UHi4aM
W60XYZyM/oFw8KLlo0AH5wmCfb7p5BBIGlIkEDFweEqjP7ckJPIqSUIwrXndx1w665TmlVC7LfPB
A0pGtw/LfXbnWIDQWglWD7LJ4mn9cKZwXjORRda9a6W8XCwwonkTPbf2c9EFsjJh97IZt//KD7bZ
loKQSJ7YLVip2XmanGjyyjkcw8647kj99e6/Tjw8ragDp8CT3FO048HoPrBXAdwMWbcotLonaNoq
cREiIrC4iE3M7oXmK9mYm0nSW7MOAcact/ZO//BoWw61exq1AantS4nhz1RBmN2oy2e95PjsYyZa
BwvE2XVeDoOEAWZ/k/65S/3eXTFEVZYnP2z600AktYE7gMls2ZEpZQlfaq74JLFcfM7Z77oQf5Xp
WNvlKbTI8vZuKF/2xwfshVTVpyCM7XA4xQn/ij3vl6/8tkKxBhE3qqiZwSjaCmyYjYEHBhI8e395
n6PbjgC7W+mMBwCUuVsgKGxZRteM6MxVNDhQj6ArClw5LXVVVhQjDYb7qzsyvq90PT0uubVZ8HJK
BP0oQG2QhMswLX/R/JrHi1BcJLboi/O4sgzGMJaX4DIhK8/pE67scbq97goQUZ0A2wdJXVECEMUw
m6HqWHiYa/ZXoS0NdsiFIK3pEwShjtWBIYTTyLmskA39gtkttboFT1w+BzttSV5OBJejVyxr0l1c
ptxVnzIIRSopI8tADR/wx2+p+tnN9RWEXWT/N+M4qH8DaXnn/MqH5Q0IDvB9ajfoS2MOyvXX/A77
73hQnVgpHMAaIQvtHBpOhnvpXZ/+GeJghj4iBBITKg+oTLkFaEqDQC4sQ63Uq8EsMSk6kUA3VZXH
LH3b1djNaVPi+4+Uq6FBfJiZlRswnq7kdl3BznP0aKe4AxFcJ+O07DjtpgiprahdFkpiUnnj/F6a
oTUK/up/5AYql+gKTfjs1uelDQDJtADSIC/HcQQqQedUW9Z2IlltxUxGUdw89asx/Tf8yy2J+6AV
VIImlsh3R168R3vGigNrPnCnUDAKtmc8NqeVPTgVLCW6FIxrMbBbPPkdbRsTVEFGMOhbaG27by5u
9ZR9kZNvMGp3ejchdRDuNvkUs74Dsk01zh44rB28Vp5WJo/PWen8ILkM0mmXbh7sKwZuMGVLJm1Z
rRWG6BZ8RhNRGRhZe/bLwfyOI99Z6UtUFkKPQc6Kp7RkK22OmsAt9H/eul+e1PRYvmBDaOyLOb0r
jUb1gjeB6dtW29bF57o5XZlstPUEDn9FAFbBHgPDa2803t76/c3nZFzJ7JADw0Vf6TW06NqXhRT1
R23/PZgA8EtaUC6VwEvv8hQolaiiPjW6yaXnGNO4f/EHFotNuita6bKgj7ag7cix7VLYyhbCMe7z
TRu1cjfytAC+52UT3Z5f3m279Zc1dMi2ye9NQ05ya5zsPlYIUGouhAKvnM8lGy+C/IgBzQRZvuiB
cvxPUo1knuYZ4TZNX4fJ7/gisrGTXhWWYcJh1FCnDFq3eMBH7f4EluVFsesTbp/4V3yzlA9jxT2b
wN+RKJgHi3U6i1Hi9QeLE7uVxQXJ1BbWV/T54wLshjAZ8uA6i5wh8Bz+w4pcF4oMrKAgdUHOG+GC
y1kIHrVOyYx/uncRGcXBV9NF7GQggVWWVGM1UJCMim9jRkcGn4SgXsIbR4xKzixGj/B/uy7ML1rT
5MCkXVC3tYJuI7prAO2JJkKdyJztfIUimmcq2/vWqMK2tJu4Df9QtkTGa/3cdhw63NVxJA9AkWNc
6uFzfAcSFIX0+fn4D7ntf20zNnb/YNmScL7JvsBsSJ78pMPdq3B9soYDjDRsew9VsWowQQGBQW8c
T863sFso8BXOurB5T1PFw7lGNxGOwuafnsXt/l+5EFkP3HHC3QaV1Q1EobNrgSeqh6HUWrbYr5ah
y03WKXZzzap6z5NPT+PMIiyA77fN1ioLAG4AOUgSfaXjH6Evz4k/nco+2sLGiEQr7AxLLD0FnOcS
FnOZNGe16tmLzeq88YBHuWgigWRH7HFuPEW3EVUoYoWdoFGaksp9DxFxkXCw3WvDxNePJD/Rooyp
9zCim9rukZLg8O3gskwi7Une0ngQjCyT3iffsb/IwsjLu0fw+eMcPE0jbN2NjIX9XRx9fUAB/e8k
W8NfSZDdmgjMcteO+CAHF8HiiTtXqhNgQIQMe2t8BdU+sN/LQp4Ivl3aK/k88iMeONREDPWcgbW7
p+DZU644adKhYCLVeOhfUQzLY/Jdb2EiRPuHg9N4cXAXwxYiB+vlVUnorbTm2BZYMEEquAP/wRGL
egOzbQMl3o5Go1OKdvUx3Mi2TbQzYEHUeXIu6vQsym1udgKXabVzUmW/OFHUs3nWxm9WiJKTkKOV
EFiZ2cveDMP4eo3jc4IT8vE/4KZJfvJUfC0ZNiTSRyy0dNPdo4cR3rxXtsE3pOaVwJgYw4UB0Jke
qr0NvcLaUb1nrK50g919OJ83FB+1Z25iMyk2wNC7AKF3qPVbepKqqkawm+zPz7iXIkgNFLprz9RS
HLh4din4LlA0+EBCZvU14XrlcM1bYaAIMuUU6+SPM3tn5aeNxySCa3sUx27GwWqK+CruCux440eM
2AbRiEVm9pzWUUMe609Ea2esdQR5cY4spO1dtYID8i64GavTz8cFNA+JC7qLOq5XsSd6mowXRZ2e
VFPXwveA3HvM3eMEPUo/cDN5kwAahLIVrm5AqDoduQ5myxMeJvk6QXabbq3W9uEIFMv4W5lHdloL
AVbcPjfoQrcWgyef2YCNx/182487PdbHBx1G38EvQP6DjxFtPRXF28Pa8ZPMEUC5DG8hh5O6fpQ8
EFZK9aBFeCnPZk7uS/FzUe6X0yQWU8HEGmdOm//rpebd4gBKT7AQi38eiLctDJZri7KQxXc/4jtI
CvumkRLNKGmJQL5ceB9ff72BVCACtXrk5D0YiLrfJ6dUrOjAJnbFz7riNW0RYNf1YJFGmvtdaY/i
1PQo3zeSzlC5g8oRMvlIA2dFpK0w92L9/zQQ82U4XWamKCvjv1TPDzfyyLootCpWujCBPW777lAb
JWvXLE/7PSvW85l1F7jxGbfc+p7IkwsAINForvzW2U7sL1QrZkHQ2R2t5tgZzPZeD+/Q6ZovlC1F
Y41qu92KJHhC4HGuXNb1wrtve3WTuKuxLp5bD5PFPCY5hTL/3hjQBbrA2YVoF93JYZ7u2zDC1svm
pL6UMF/hc8GMa3Vh2d0I4ajriUMcKUbCW5dDclT243pzbUg3FuYSvY6/uR5gzc2QgVy3Qxx+KD5p
BrSG5I+/dv6gV0BiYLXrNy3FVqXBQ2O7KYy2ZbsovWCPG79s6oW4Y0KW1oD2LWvSKDWSPi2QzbVG
HVGl9+/XMKUiVgAv9xwbfDwvvXWNZACU2VE5LQOL3wn6qMJy6AiibQ1HnAxVBgsr/lGQ31vZQK11
AJYGck+A0JFdMYE6GsS1d4OByzRaYyUFM6W+ROw4d0TrfP++spAS+Y5DBZ8OJniZqA5jhCByHWZO
8N2yGKIzgc/oK+9vVpfdUW+fSTtmN1K3OLFaJQ0lorUiN2wLljPNE3vhIHic+Fgw8pJ4JzRlCsmQ
5IIa2wiNwYbjfUV96saung8BeBReWIZZ4Sr1mdUHWJT1kS6wc6lRUJWE/+Yfi9AbBTO4YxNGeurj
gkCFQ4thCakIjnnGGcf/6ede8xVGDKgSz2muli6rt2Dr+yOYITf27RujkYb5FoPx9HyD11YoNNmD
Ov3B/oGAPJAUzfl2u4LxG7eG77W36T7TdhMD+xuXP0Bx4xC+4Ov1XefvJtcJClORS6gJcf3Y8DGe
O+AyDAMtRyt9m/wdk7SneLt4NUPqaVymSwxSNXyu5hXO3X4CUZqCD2Yv5OOcND/nPvTP2cXVZ5r4
wejjxdcxTRpCedDmPbQc85aviGR6VruN80+IiwvHOks/LxqxlpE43Q0+7HlLhkmuWifn3bmbdNM6
gw0pQCksaTcbISwsV+fnbf2Tp60O/nZcf2np4xlZRHAmKIWHtmxZV3ojaFZWLf7lTR/gU/LfzdgO
3yqOSrJTk0PwQAov2zmkEzu2tDTP4efCii7f6ISZzBkvmZmioGDYnY6tNr8L1331oEF2UvDDWbPz
bp1D5V8hkSPUAdVwCmPLOqo/iTU6ir6GSaVz+HpBgbcUXFYrEh6MGMNQl3L0d0d2kJwIoUu1+8nk
f+0bPX38suGF6eSBxPLWWBAnVQimdts/986wUs+6pVmgXoNDz05ay6brsaILauM2GVRskvrKI5ez
q8XL0mgXHaQ+w+X6gkp9FY2qZNEBk6zlvkAYMrjcEvJjBdNdCMDszQ+cOf0bzC1PDtCyF0/iZXei
ObVX9TIKQDgo1KiT/hTUIlDZx+dY2B1nIyMhhFFK9E3HCZhkjQMGzdkqSNaI1cbp5jfh64XiHMa/
J7RgvpJtdZH5ecysrUu+josQyI31+8lZYhLJhLumJADxFj2eHfNzl/DJkHASbDmlJBm8MfxNFJmA
VUjoAutoZmkmimgVizwjEosK+rswQ6tDhEpwjlRgBG39G7wf+QYirEG0OK6QOjs+pqkXrthU3i42
xJd73wzcRTlFZjY9GmXKZd5j/ctDygzOEAyyB+3njmOQ4Ieer83nkzfvny+Owd5Be2o7V4vefaSi
fZ9Cfa5wTzdNduy8m+I4TDyA7cLiX4U+pvoMMTciG2qkf0dflGXRdfmeAwITHMSdkQBUUx8CaRiH
m5PMgcoxWXf/REmI5Uk6J/FrL+ID3BX1XiHBcIrxGoxquo0ZjTTJJKoOBCtAk/zN+b3EU4xLUmYm
E09MIGG2VyKOF68vHzIc14V+8V1LGOsprf93bcEqPzTmx2UihHhw6FXxHMOlW2iVrj3m0m3ee74j
oKH2EwzmtuYQ5VwJpz8hS3DYkt0NqqyyR8f5zaZoA3JxKFAebJioaqJKymomk5VTek1jCzk5WA1a
hTa/ONO2N69aaCeZOOdOnnpH4p3WVu4/sMEuCLxERcSg8CBkhqbFQdPFRRHb2PDIXFwKs52c+Pcg
oxM7JZhVYJl/4aVvmalxQ4Kq6k4ffvU6mmOAlk8gEKAsGEiiRAx1fWcfePEXLJjNQlWa+CxvEVVC
0hu4D/mH+C5cKMy0tUVdNH41hOwdI8vFjJ663bTDc/BVv7sbbNTkffkM+7zys+YFE4L8F4/G6aw2
4cJDYc/0RU6/yZlSdpoeOjUo2V9cHUdHtBCYto1JuRymsXiTHWb7AeyNoJShzxQB0ccGuikv77wr
nzvb7KKw2vIAoDZ8TqtVlHzD8KqtBeEGfn12tzX02AfXy/HWH2VU8s5p0IfugW1v3uQXyulo6t8Q
xpLBWWOpOGk9esFKWRPatYkJCa55Zq1mqnp4T3VF/uidg5xw2uc/PoZtlkYRgUmo4Rgr11JwN3Dq
KQuBKfF+UgtDZBGpwZEZvZmazmGnK4iO7tF4pLDKrlnMmJc9pGVJ4wL5mWro2AaJLIxa5nyUjv6J
3SUu0kmfHjUhCI/Ba053tAzLSz7SCGXPuOS8+GzBswXLPQTdGyqc0/AjnhsKIV/NYri0TGBMT0H9
DXSrgn93fK7C9P0Qou5ftW88O4XP45eeyleqsUcdMEjTYE4puKcZKcUsC6fJPDMDEkxOqVxKIDSR
y/I7yse+0qz/zzTetkc+aViqMuigZHTh6hO4DJlxVhvLKrZsCSXizFUr+LPfiNXUrmOJn8k5MsFw
svVCXDZFvn+RvDvRx8dacvWXpehxPnvzD/pu1IuMErSXWdwJqwnA0ySj0OnqWGZsJceegv39i22n
6ecnZDE89WNx1nmYfQXGsDgrSSEPpTvwYPpfcw6I2pA0DoWwdlvoSfzghOkF7xpzxWyRZ6BALiJw
uULT7RT6IUDAxdyJ4bZZAdEkf+/tEjfGFmtTH9xA8AzQTlwfqOiLEJePzIS4MSsg14Qc1TlULfog
WxKM7jg6LIdPDQFU+dF69f1qGR/rCqTRLqoAtmyVMVIRo4R+wbkRSBrQXfj3THqeDVoHnZkZRlbG
tEHaVSvN2Wpbhgzv27jXzkTO7LRUu2b8FlHgukgxe34L9zFMa+kB2AwH2VxTbb7XltD1bB+xgifk
eRXi+oEC+3nbmO6dozAKq+yxPtS1HYnKGvBdTpzSz8xOQQNcnT00YGRIOQCJrKb65UQKV5E59q7N
ZtjzAUEYzEhqKZRhCWzowvgkxsM1vtvtDCIB8urWCeRTAOvAhmWquqdI1DXIrRd5Q6K5Q/EdasqT
eJb9fEMTxmO84o7SH5fHU6rpTmj5qSPwkZQKNIUszIPMu+cnrvgmFPlNUfYkR35drZUOdy3H4UMx
dTRsWLSpGjpvkF9LUQM76RLa8PVkafbdy2gLG33jmd1rkHEHPYJO7txf/D0LKzS1k1/OXsp9RF+K
6hn9tehuFpBb1vjrFHGYLdkGruF0MSgGly7//lTk1WGg1ZIdc/b1+KWtRBVnGMd6FMyuyjECfbAv
GdD4aFfjZfekYZeKHE5jPx/DEmpwe75DFC+8C3vs85oXUE17qZERf2eobHyaIMjlwmahIoUCQQLO
jGfqignXxwv5jsVwlwdd63jq8CuAXjRVpFZAugOrH9A8Y46powkrtrTkstW+DbVQX33RqQvCSpcw
aA4GHpx5i7GnSBtpOp6umYWBVW6PYZfWd81GzVLpfj2qlRCiFKY5d9Kxn1mZ5Mv4KTZNtGgDXhFB
f5025dY59UtidxJ7pAUNb87ljorkyFbuW0TS65TBXuMyW0DAxrmsaf/u4Ge74hgdjnF3qfAHIeqz
jM+B8NqwM7UDjwQMmqNi6CIZqmQVv71uB65nBGjtTwe/9I8QVdDQ2q67waBSQP6tNS3jCbw07e+O
DyiflbSi2nLmAGw0KJdi+9tVoczVACZcujJO9IA5FbLJj23fHvAGqMsZwPM45oraoTmzOyAz5FQb
UfINzulRB4Y8qIEI33zleZmx4ofg2QKn7iQatHBjQjUhz7sGJAd40J3ScTFNJOpZlA9Mx8jxEgET
inQfqfsM8ltyyiLYTy7+74uBTKu7CK+9thjKqyyuvpA/AQhkIfcqfuj2EMf2Cf2Vtj0lawpnfrPy
qQvt+OVHlKhWepVo3FUexZ5yZZJW3bh1Jw4F8hNRbGd/Vd4OjAXQnKwQYAe7aFJjephPOOVvg9jt
yvnziuE60JhlstWiR/bG+B6TSDqh2A/h+MvsoxMtKyGrMWSIRVQRuzPXmPev2ywsZYzOI3Ua/ChL
5kWAljq7V1b2J6FWbV7A8JaMlGaMKbZBEeSfreYIfciEDf7Byb3Jtlqx7k01U6JjjST7lBsL37GG
ZQLaE8kJWN/FB424rlYqwRldctqKe7l7XfdVhmI3/WcI2veTN7wQGfwvFEi/NlwiNHSyELbSJang
oY45X+nibE6eiGL0K9WkqSK1+7SFwjVuYsV/nzJeksTvEvUmfqiEKn6DC+QNTON5nKeSlpFxGZiP
lv5ya/87MF2pIYVS/MENFvz2e400GIsP7tZ7yY4cpb4K/+PZDjE8VaNYMeL4TfJWt+o2eR8Idaqq
fp+0Lu/y9LfqooBc14r25KfOxMavrzKeTeEqAKTOx4PLjkueOEds9LsR4us7KdqKAvBycjG+dvQi
uQzQpJnD166up1ZYT+DdkNKPF+3FZmBg7IMyOUL1E9Q8ucjOePYTAaGW0qV8DwGYdjilp3wz3DMi
yKQAnyhEroink514UwubQocpj0elQDzWKUTSyQxhuey1b4kmBHRjDQDHUbhGH7ynyIbI20WxxUYu
3LXI/1VLt1sYKlKs7w13Yuue6co+OasUTKbikVHtSrw6QSJYEmaaVPINDLnYqI7fGBHG0REORC2d
HgVFX+1Qzmlm44yv1BQ9E7n/rCBlLOLGk8o84+BgoLDYTH2BM347Da5WSslNRNIw/b7T4lzbm/mc
KhEr6WpOxIqqEhnev51S4JhN+S46Pr/KnlyKU4vxTU+jP3XQMJmrJsHHFU01kDTY03TEjqKPSDm3
F+RNcKLxKCu8u6xMkcqD1gc6PpOoFTlgHlDQxaBRJkzt5gKU61LhzZrvFUlmBPo1zXiIJqBf0YOl
hsxmexKTxrEeTJnimrJJROn9Snuswf4Im0fB66sRTizGXZjFtruDBUiyQh/7IPDrna6qK2wgREOx
u6aBoYSmGhyHauxcCOFp5t707ViWI+MesliOxZWRQEU1jOXh4xVev7QXEcBPiGQrJpwMZUZ7yXr7
6KvJlMAfsfWEpEyQe8GPpAktl4kVVNKowkt9npTQRATmZ+Y6pXUFjl2lFSvnr8PBLSMqYRegs7zM
K3okJ/CHOzb9Vca66IppzpKskgdaJ70MnwUCfIeF14Bv8n7MT6iWwg6LAOpRyScntMURDkp7gb2C
xuozIXOkcUhC9EQxzVkGLFjhKiLwBwpeNqzT616B/fD7QewujeHs73uv74cUfpQETZw86NxPvbM1
smPjzQosYV7wyvL3VI0qzl+01wMt0YDiEIRe35XscaA927FDWbVzGOrF8jjKXvWEYGnGxCoz/e1K
GN9+Fd66r2BR+U2si+JcD+EPMsdhWqaDNS9L+fbfwK1HpXmkQF4FaMolpC40ksFwDJFydYvFD5wZ
DnzMQURD/kSr3jCDAHTwupy6l/+/Sacx6dWDyGC9vB9kRxRUi6Ildwl0NLBNMXFJ337XtBGs8GVx
HyyInYtjlLB8LWMaHt+IcfjMP++P12zs470X/OHgXlMyJ+1nt6DbxrIJTAksUjgcrDEHP94FTh8f
AM4mYGbhQeqZ+7HQEjwBhI1PBwbJ7OL9jIn/BxLfgkSxS+0IiVDI6zOElFywPdxffdSD336Fe2/X
KZ85o9ZHpk7UnbdlF0TeVksnG2EWYd2AVcjPoZyojeyywe4VU3zgYEqipYPUJSsNMyttSxyyZk6x
XHfZHs9izUS1sUwAEUuw/aK+pxYA1ForQcPtLTS7KLdPPen3bSGPEMBrnjEDl+mmNgevRALw5NHC
EfCHnMjCQdZT11Benejz2R3RYMr8DKwFMhSG3Rg6M/M0YxX4EPQinw3K2hP/f5DUMX8BNIyice7s
Tn1x/mvr53dwJvnewGBm6wNkzDpyrPdE6jRNEEAOGXHzko/laPkqo5DHadj92hOyJAwVHsjCL+Iw
iuYExvz2Fl8ygpBx00Gk2P9YuvtKXZxG0id93+Xl6pfPVwwZCHVCNgZ3kv3818C6jvLWBLz2DVXF
kx20QX0iBmtEFLnczM/JKIsYdZSevmf8Zv4d2OWWXjxmjWQ9mj+JRE6qqjkvWlBmyer28jEJ8ZEK
5eXQJch5cPUUYxbenlQKTylrohciumaz9mk6zEGKUPdcvuL40mAEjQoM23rsOkrWGjyPaTlk6m+x
6E2LUG6XqfDNuiM2CQHDtCFGHV0ckQxmKQjoaU8Z38miWpiUNwcX/JhTg6peYMCtXix/qWFmWy2F
2eFJgj9QzwL8V7cNSywc46s5sCq4mHjpRTwjIjpoL5EdkYBqK9pZkHmBCZGsrT2pHqmacionQCnV
Quv2+ug6ctGf6Ch+mFEpgFkD3wNTRLsyv+QO+hYndkpCSA/bueXvPPhSGxBGM2JY6/gKNyYB63Fj
VeBeYvbTu3zXi2zAgzL09jqvqyaF0YaOE40BnTab97BXaf8rLqkVS/uaOm7xp8GgLeR0o3VQsUDn
d5+yNtIVDE1b3U8fjOAtTAD3Zm/bb2Qi/7+ZwkA4krlXA66KLbPwbV6JizuQE/2GhepXYPiuz4nc
VcmXRYcm96mY0nvVMJc8gySXF/9QkMo4/VBmAgcRBxQhw/XBMgGx5l7XVQWHDajyynBXSX8Kosti
E8WAxVeyKWY1EWltcU/rQLMHh6E8JIHrOr5uv4ybCrNNgg2+oNpQ5oE/JdTQVoxDA6uZjAnPRLw5
ZQjLyMtrmM8i3CmhO+tpf6UdGyXYjJHEYLXAoJyE5CdPOnje6QbQHcwOfUBHajOGecahyys4KiEk
kMqiGv7hqYgWqJtd3qregZkoiPFtNrAlnQXU2tU8T9JX+6QeX6BDZVHNaZ4nnMtirwboIGpc0Xb2
X+c/qtnMsMpezSOUyp94xuuPkROH7jU+d5oO8LzEjv0hMwyxv4SiamjimzH29oywMwgg52nTwjhg
9wbG005Nr/7PG9yRhbr3cpuByk5wKH+NIh3ht8+DIAh2XpoTwIk5m/dXCsxombaWl4O69O5+ZcdY
gZR2MDQ2r+BPGXJQ0zf5f4h7xGqo/GgPeG1wKSO7tuNDtdBzFYFGgbVxic4sC+OgXQSXP4pE7fDX
aFQj4edht34yQmUie8mbzGSRz/guoczn/LmZ3hp2L00gi2fB4eFX11Eh9IphopSJaDxLMVJxVieI
/GlGjwvWTNWv9cb2ath5cUR8RtxOqseUZLujwo7oEYqHjPFa0+6kwYKXvat1TblhXNreMT/qIJYc
H01ZtjmYpVYERKEZnlCKShVoZcdMgX74ya5RwqWVaHlcQchGN9f0wSYemlYK+0QocfUWH0TKieXT
S0fj2Yjdk8b/5R8J6F2fgIEI1n7as6R5MP+mRymMoGBHo2Szv+B2AiP19ErikRPnihEMvqzJCAqX
n40YzonyWb8DFCjzjcZIIacKPevLh+adi5KHFiF1JRT/joCXI9Yf0AIGjTMYKkwrPSRM4yTCJB2P
WbQ4k5+cgZ6D4Z12Kcl6Vr4uFCqlSIeA+VkkRZK2cHvG3jXAgjjCped4ZCxePd/TPup+DImWDYlw
91+EqXzz40KYGhSeLqr8nwmX0DiCtJgQPgBBAtSIfcXrSsFccKgJryOW3JqqlirZRu3hgUjHASc7
DfVibgFVL/8tBmFYkhVP8Pw43UeZo6rE6t/P4hF+UZbukoPRxbeldlEZ0Bk9Z9m32/CLkYqUF51x
zITFZ4J9frUrUeM4s8spN6J1webnV4xmmrfswqxyWuDl2kh5VQR0+e4RqLnD+YD9Wy5PY/P6DZce
fWyOGmCz4AFFNKLYy1E50Y/3rX2EcPYdGcro7NDQ9Qm/xUIU1xk29EgkVeXzgzaM9HvM34uiZlNq
DtJVMPE9j8bQ7HC10GzNGvjuLrGDFrKUYzuvI7TTqkAGJV/UGKobDOxnq65/f9r/Dsf7Qk4/YHJX
OQWYKshWpiNAOXzAUn/A7YnUd1uJtVumCqVzqDVImCE2oWjaGGGF7ipq6ynRvpE6khzPc80+T0/B
IMpdNCXF7SQaC0/+VO+VFA2Q1lC+mWxZpei5XePnV1p+uHzDJiU1wLBE9HvEfkd1nNebVTliu34o
ynTL5paAEtgEof8wH+gZqufKWxaY/iLXO+VWDuioF0iyDi9URwKlOlMHKtuoPfEj5fJzR7SIkkhT
JXUNoOuuXCvB8IDZqf3ToK6cNxhG9RSwPsrmPuRhYFP780jkGJ6Q31HABC+lHkowhbjqvnC2AJDq
TqqY18eR8Wzzsk71DZnMcSkxWu3585xopatqWh7OWHeP2NsEBZnOTu3KgYBFjQW546dQWwx8BC9b
yFEkHafE+jlAiz8nvoOFso0PtNPrrlI6ky9HS6kt1JcP1S5WpTKbY0MI7s53kx1hkfEnqreQ/atB
1jBB0IyMIePLPNEs1axU6YpVYl4qT90bc9zYFQ/IwBZ90qT4nlkuM2B6/uyh2SWhaNG4pkCUd1vM
RB882hL+XjbsinXSF86JzONRfXt27ZNerELab5jE21/1dzapcStcmqJ4fn2NiOy2Y+bktrepZm4e
UeHubi9zgaScDUWIZ8TDT3ekH8AUpqf5tz6i8TLWZhlpWX8gnEmgx6czgduS1Dj/HopikLMHLhmg
CH69qBSN97wsdVX/nRri1xFWm+YDg1QnxLZbdud4aSJzkGaeLsAVNWLQY0b6MMHu62xSL6xMn5lE
KctnAVhR8UoxTA0lubHtGnFNaRWO/oQ5Wxyp9jhJOhZe5ouavPoIjJxlI98sW4eKnzFCEa44ZYgb
FTAxnhvjt8ag5m2WIJG3woAnZV14OBFaZGY6Nuc7uxzYvbqoeTSME2xNf6lgE32jQSP5vFnRmDzc
9Wx2vnxlRBp9LxvW7DV0SlwzxYpqrXT83mgYXJ0Jy1LmDMp0EY3gUxIfQ/f4+V0mygQkNRuz/NDZ
H32/G9priZYrI/whju+OqHFo3gxTTSoscxikicoaqC2kJtHKqgZOhZIP3m9mdda8qxHe9goroXOO
jOnIcgFpELffPBqShzKyFaEqRC6LylfsqCfD7Dno2cDIuAmGNkO8PdPtQvuY1cdMAp0XZbc8Peaa
kI7ZoEWsIV7tgHFgzNLq7NxzJf5BeNYGQ5pjdzT2uXK2T5Gn4yc+bgIAoTQqx8AJ/oKnO1Af4HcA
CAq2wY0CsAbwH7XvSrdMUCovnZQlpUfCPu0RNvt5Ob4yYEeSk8CwWwTHZ1HsbyeBIhZNQZ0P+GJG
HHCSg9CpB8D4vaMv4JwhXi5TOJNw+ZbPMvNcFrjZe2kw9SVQObJ/cXUOO77OYlmASAEv0ztfWnRp
LUwBuHaJyrwsil6eF0Gse9P4p1JZqFXbAnI5xQKPRbWFLMPp6TMABgBTd6WBX+OtCQVffPnsJv8E
5sZAvlxeF6jvQ48/8F+hGhL8kNxMrAH2ZoSW/Hw92qM/bYfPeEG3VDjBE9NK6090TBqeGjV+5NBI
0qSAcsnYExkNdP4Q4o+btvnYFkiNff/trtyqeGQ2zLPgBrSaJgupSly7ceJXpRF1zMct4x53IVT3
uMkG2QBs5/B3W2EsReXj3f4gG07w+XO078lEbiYGqc7eb6nwXi1zucDhCxBumjQFSbUGF2RYSchv
FD26IGyetI9Txxc+itwbFtvKiyHFoEPnPsmB7SSmkLHT5EBP5P1YhAKZ6EhisyFgqI5sXCR+XaMY
NinBOS5lRci1Fum5e5AgFhsgEvIIYlh4/E4tnOcAW5Hahdl8pj+5MFUhik/KGFIx0UO8iCMfwfhk
P0uScZCbQVtCBGvzQTxck/Ao3ZUUTmfveb0PjkhHmAboR3chc77EqzBl/L4dGWA/s7uoJHRJI/jf
x9Gq70DaLYbBANfRcN3PlwAQAbXFLXudahhgEJ1AQIyApi3wHZmP0FoeMoKoWX6WF//zC6QV78On
zHRN2YG+zvgtUVgAwGpDFbeFARCbglwodkq9Z3oez1ktbY6zHtqevVmYQ6qFgI0d3oEN54f0VQEI
Rr8LftjckWDOtXUlGmF87QKKj2E5Uld30EcyP1/mw6dT5xCRlaOmDlZkVjtH4v1kR2r3/X/cy7PJ
PtEVYAeTQtV01ro+xDNxEEGRCJunNNIExmytDRMYx2QHNxZhlftpgXrjH6Z2imDqY7Tip1IIWLp4
XQBIffI9EAfv7pWexRFU5HjtQHHukyA01ANMOObP90WrYNNH8RPRIrV6SrVjcuSGCg2csybzm1QK
9MKI4GADnuMnEDRzFBaBkjxf1b1BR98HjMZRdZH4Kc/wvanESnQ55BGPj1cAjG9B4c2vlW9q43op
vjIYzxx/bRaUxNizExq+y2aPH2grbl95kPfguIweD6BZeTRDO50jUd9Jew88xJDHsnVl5WR8qKw/
RNkBhDttF9wOc7c5u3ZM8YVMC0YQ0dO8Hnmrft3yY45FO1jCI/sCQRY6XBOr2iyHYaKfJcWXimD5
en9AIsLnv2E/lK5qH4A+dHZS8ifFZBJj/KfP2jnUEWfDU+5oFi09HhC7W0yaWeizjSGKWgLcyvUt
r0zaG10vZdHaSTBozcH3xrXmtdeOtjyNwRQVit8zmmNg+XWyb3acuIyyrYZAascOJsMeyNzGjkfD
pX0s4EcXJ0wTJPHTcpBKm4yqAUHn0nEjC2/qmaqEuzA8Z36TCtFgmOylnYSuHov8NScUAcVAmogs
qT8WXRrqASPHENEX3SxDVc06cnJF25rskE4YGDVXsfG/rYfofLTw27AmuGnKGh7QRU9t+hZ672d5
TtPsuIRmw9MgT20QGtT6v7bshNZhJfDyOT5gkVKsJOrtPA5BxHh9ufbt8v6C8fJiLxcf0uQovT/Z
4T9v9HsCJ51UL0T8NG1auroxWKrXPEotPUDPwJ/CDn5z4NDp3SbPbLcKXzrMuYPlj74wnF1BYLhQ
yAs+j09MEHSYHWTmLYla/PIH2Zg2rxMiCMq0fOapjTcf5UKSV+/m2Y0cLnN4wGH3RbhvPtmr7PGm
z8VWWaGaO4/NZkhMPCsENYBpBNBhukmFoQ9c0HHeSmtlrT/mIFcRYlTz1ETkaCiXFZ+n0uTilzGT
/P3QC8aw53RDMzOpiIdAuNdM3KjBWkOoar5RWl0j5V7fPzIO/5NmGyXea1REy7Kj/nOqO/i64hng
2JN0tPviZ+cKfcjrd9PdjFHkMQZ7mXeZ1rcoSJ2IE6bRp+CvI+NgfyPqLmhFL+FtS7uX7Xs0Ddy7
Sl7odgUa8W8a/4CbmGW+CzQ1og4bbGxKDVmBgnqst/vuOh8ZtZmeTcIZJkzrvaFFvZeIMBPVS5OC
HMFmbgQ8kq2bU4iBGC0gnAf9TYf46BkL5OY0/FKn86dJi6zRLeLGiM/QwY5VAGJdkM05cQ7oA6Tx
ox0zes2hs8Szyv5H/mazNYJwN2eBcvZUr2I6AyJjC9ESMyLUlWHWuLu2xzgC+UsLNw/X7KGTh6Zq
6sK/AzeDDDko5m+Y5kgv3FxRiRvsBxGapEn3YrHekvbNEP/sGGULPImLPsdpwvAX8xRhadBAv1dA
yBD0cAxeh3VLf7VPLmTMQHBQMQ3sIhNSgxrIqwWwLGVZnyaQp62a0Dm5xjTCApuey9Fd6zijJtlM
QDXNWnv8CWPH2QmLmmqL7/jgkmoEysV4GMMLBFKJodo4w7R6AHznbAarOZoMvYX+AA7jPQVHNwmB
5ukKqMTYFH0suvTqFe5km0OSVwiTR8v3CBb13VRbH/tTrmuKQhq7hqQVzaDQGopVKy2Ctl/GRVQJ
b/QnF3GSGEBZJk4837NM1PwG+bTi/7rxfaqRekMi5vOPogJOVcg1mM9LItozw1rBjLvjQNMlWw6c
rnL7/3L12HkcmIDxsmEM+wPEHT7w3P0wZJGK5xCDJhQ3teU9McRQ1BjPwdw2qk3AUqPS89kKqrom
JRrCX/eu2fxcaTXZB5quMjvUBEXqtNWAYBpejBwfrcVl9/MPVN/rhcuOk3YgGwFiYntsRP0YJhSH
ZCmpBTopJLcj1kBthT6hlUAX79Mn9MCEE+5almoVZ/zebV2KKErhgI76RXIQmG9qTS0HoW3SUDj6
k7VjaROo7NzSWLW4wJbL3POlGG9qVYqv/32XI+b+BAtvBEDro8sSSsxzV2wrFKNITNPROI0AYr/x
wseXDVs9TaLJddcK2KB36b3asl7v7bxeKiu1kLUbk9LC9w8uSoUkV6OGtvwqWDIoDBTrRZDr2bz5
weepgM/xgTDTsz+cri2dur1+Cj98WIF4LHPWhTMF9Stv8r7zxKyY2RVLsdZor5mOrLhquJd+rNc/
KHLhiblH1T0y/clOsyjneXcAj/1i7ANrtyBQlgoAS7b8zb94haAs4KRyVwSI1ik+nnavMJpv56kg
m+/2D9QP71VAzQjW7f/J5PbFYCBO0NxrTmHOLs7Kbqli9PgLilYc3I18NZclMOleITm66AU1ZT0d
Hefp6i4mta7Z59L+riiqdJqozah914p1n3fyRyf1WImg7dvcJe9lW84DJ0uisuRpUFRlyf/X8z21
vsS1QwkryYxjW2dbnD3RNT8TydXaxjFKpj3mxBla57JtBvHegoBXi0+wkM8dIyv/W5h9kwMMIU+u
rQRDspBBybED+ubHayB52BOR+wemY9+3g4KxsuL1OK6pSMuuvy37ZzcMX70oAjtmzXG0MauKa8zu
DlmPDsy7t7UbiL+J94bJYLZEvg/esWkrbilFZBphtC8UmgXuR0ueesdcMvN/c5s/fxdEwfEW33l7
BSqya2SX4pHkGC08Dafkk8pr9s+FwUIdVNFKfFBxNnJ0vIscwh1yanx7wu+ARjAmOX23vhLgzPZf
7icc6IrIi4NKsk4lho6N3momyDwNkCAUezCauRQK8crAmzau6oGap/6B8Qz9fdvOyosdNyaH8BdD
wD2zzsppvAjM6kIC8CjvAbWKZD3Gs5XuoOefVroG7wQcVLJS6qRgQjE2majftvmScyskuvdibSRD
65N+/E4pt11IjSlcFIWa3nXPZRQOal9ixkYsgqZcsGVXBRrgLQrhLvo7srKcNs1IwAEkzFldX+xV
cNKmY0yyF6Gmcvjaaitm6JF/sb/o5Ol3FrpxLl3mR4d++foEO/xwzXm9vP4qUGCDillI2L9SwOaW
kpfpU9V3qnhOQKIwndDLgtqDRrn2dDfXNoCjkOA8kfDvgb5OQvg6W3nigpu026mwM86mG7s0LQBf
koSQG2Zuq6NgLWJv8NgEX/sI06H8AGm8gbTHLmwbXtndkfAEoeQn5DVeuxkHpdePwM4yQJsdtK6+
P4kwxG8c0HrScow3vgW8zb207Rz7RLdxDVaCilSVaVn5KticlyIcjgSrPtwIp5brRS5lUmFeWWS9
TVCIetXZKBEd1aGUWnx7LlANWi1FtI9EThC8EwkdVau0UOrXVhATv5cnjuopS9nB1sGdch4PyD7X
wE6uegIaHneUYcw0uegi2hnAXM9Lov0Qykr6lokARTomhA4Ym9+1IUvvq0R1/ftPSciV4Rip6awL
o3PFSq+SyDCjnauNow4S1ymh3BzCdvYBP+3LHgh+rWqCeLrpWUykq68xNBlKm/qTWvoWDurnsHDY
S7Ir3PtGsgkue7ONaLEcOzgTKPgOtXg781IUt2PdqXMkRrPtWkxxMnd2mCwR3jnCnRb8v63pAzIi
xvfu52vNvTXbEtcuGCKAK5S1bEG7cwM4A/IzUUwOeO1+V6huit79VX1tmOKsNhee8XoxBsZbhO9k
reF82nIwmQIILhbsqSXTlnSAf2Jq2vPjWYK3k+lKHC9kYLzipMgdBhJxZtAuAqu+j6cQSeX9gs+f
v6+HQ9KMrnGYiY4IkUl38aTyavOwFKDBEtHaNivI3CDZdiC/pc1WREbPNnDFcr7HnXpczl7TeRAT
IYINxk73WgxjQLlhNHijYRIQ4+vfZg6vIbU6MTt1+7aqEPSqgfLWMeUHGNqkVUCSUwqXAUzMQvfQ
xq4S4yTiNkKcOF6Oa+XqjuYyKMf+NHI9blIsyqMwIj07CTe8d8Z+7jYAlsBI12HeWGYppxBtNtxI
Rkx8XCUp/COgEoKxnLTGpeiqCrhTBOeDieJIqPb6prYnjiv+aHVVoz3IiT4Ld1i9cMKZRZehwep8
eHLDp6qyg2yIjF4neaKijzojBjNu8rhBOlDrBQcTvBT7/89xGpUXsvNFuWppsHieSor8wRr64trb
0onNLlVZkRBniAx7SXfTT7rN4S1cIRYWs0ZCiFzxMYN/jLHrc1RQYelcFxN+nIRE3fwloRRupW8x
S3uWNdeyqwEdzt5r+VAeJgF8LNGwMtSE56tP23qKafoyuBeOWWA/ZWH0BDrK1efDRs8TAGQZq54o
gcwzL62JXziIdpUpYbqlLhTHl9kNwcnP2aokU8wOc2SSt+6Cdq19o6SoXlbJ+ZAX++zshSmw9zVm
mQwCeyLs2qvHi7WDltRGaM6gEkinvmFXrFW0RqIU0cHinQyOiEui+0o+fp0zi9aRYfjHTvBoz6I7
1OSH4Liq2eXz3LwAmEMHJXLrwjyinxW4jyzf2TH9rEUC7Q5igKTiAfzjdmsEIopNTi+UPiT55Bg/
ysxGsNZkLtjCBmFJkEO7LXJntwYxyku3nLwQXrrx0NRSd52SgqkqwFYEJy+xQJIHCjaQO5iLNLYd
NOmIIJtqU0TdYsgVWVDquSKG+7nsjiqD0DHjowiPOf+cJ6Y8Sb0iF8ZnFrecek7oPApTlp7d71iz
DJ+g8SA8ZulzLsXmzRWn/IbdNBJrE3JBghG14G5ep6pMAQydfwEialooOqc02wvjlh+PFu8ivLJJ
JvJQqnr4wJOk6hoAN+TiW1j6g9HQDGbO0aqZqpG+3tTaw7SY5O/r2QeHD8A8jXBaqMwzK640sLDC
DQ4jXhc02M1SlwK00af08ckKhZ6i6dhbohM7Lv2KaMW5EqS5M94aTJRbW6637VuKI45WLHwq9ixa
mZ2D1y1kYPnkyPzVJ3OY+I/kjzmxf8PC7LibF1riE0VBmQKLkvpsXoHXRQ2ZJrWJDuIC85iWU3ad
j0MSiCmagEbzxHZ/Nna8uMP3Nksj6wHu5Iyh93O8N7dJh/SNK8FOC0xOaazpSGoImJBH+JLwKYDm
40axNTNl5bnniJsBstvqC06nRdHX6RYp2x5tlmdzYGUDiffVZUDfU4eYYJr2qG2jiLE4VDidKRXU
U3bsu1HoRHo94kfowLM17WGnREkKh4DK/Q0lrjeEq9D26wvookG9+p186Qmm9RZ6WQJcipjN4vsk
zbxwupfa4m2XCuJkjC9l0BDkjN/2MJCotD2Cym/D50NPo3zcm9SVAz3kr5OkZYsbsyhY78Zu4CKc
AHrN63WwCUN5syVKZkDWWoRbNAcNaG4sr4/KxmuQ1fXS+IvOoEwhf/maRf3PsiQQwQiRNoHI5EL2
+B9kV9TjwM5MW2pA/CPiqX4GmiazBOgM0SqT0tiO0ulrOoNhhb5nzqY7hNMIO8DAKYFlBEEdYHtd
r76t3RnDvbZPclqr0zbdHpFxpmqEFPN3e0SIlFR/a4KsBVD4SE0NtmY/EmEUxCpppnqB2x+83Igi
DZQh07D+Ss74xRBqNEEj9KitfmDU1CAwCKJThC1iJO6eynfkaNYoQCNP1bzMmeofJ/zkmwolZbCw
1OVnrEF/BFsv+GKGRivu67ELtB5ksfeYq72QU8mDI2qZxJbhf/DSb+u2aJIbTC5UuG817PW3MsT9
f75K7eUxEFFFYWova5Y6euwaB2WuMY8SANHmuOhLPehBGtMB3dTWayT4O6qCj7V+/2d8AmNw9rii
/YbX1zlkQ7DD9pNURyrWS5UeCCG34C4c6LnEoJIJ8A9M+iqp9wc5F8BZ2fwwOPnfGgbPWhtxCXhs
B3pLvQ7ovR1iFjocdzFbbwCFm3WGSHpiOFh7H7IGlry9bEAq1NeKScJ3qM5YOeuu6Rw6isO1vJs9
c7DksxtkfVz7FmGYiRFln0Ah+iCJA9pzwQX8W01F1zdExXk8qNN50uYy17Ul8fpd5KKyTQke4YTo
IREtLM5DG30MDWlcbpPpvUsOxGrbRBCH6PvxXCbvC5du1OlWnciVOVew/zPkcxWYBquAzk0okjoX
qthXOcfcUn81gZOSa9vOgy8dqKxV0LVHLxCvkzfOfgNIMRYakSWEMJj4+ITcl3ob9sM14jB5PLmn
p0omi2vmo8U2V//75RwUAF9FD6rwEYbrvIttKxKff1+oALQKdWUOUDM0xIjHvf4v4/mlpiGX/YMr
JggcVwxdpPoU/F1t8B+w/kZdNVYRxWTsrJGyh1mCeAdPdV23P1dT0vN949cFILlaZpBEFp5EilYC
UQD0ZsPFfXHCigiUPfTbFVSs/8gmWNFXTUBcXRa0xCCSvkt0f2bHzJuubPV0MnJnRgDFAH9BuPy+
2VnAgcNpPcpaZGxcnVbBj4o/gWk/2AWm86Y4DBOSuZH6r88RehHJ33R3R4QxEcelaSytRAesWG5r
dpacHk/bJPLZRJSKNRqmlmayo13hZQ7SQDgsI+12lCDEL0PdEu0jjmQBPvLpP9Vnag9uZNsQfvPw
hzI4JvAN17OiVj7inybv9ZGknciEXgqxVRO6A/Lt06TITGTy6m9CsvUC2fhVUMj4AgNoqJnvUGX+
hOg2rqVRwhKFfwyCPtFaeKMxx5td7Squipj+Tk5zfXoyyM1aq+K0zjHlIQlBoArZerXiSwU/D8ik
iBWo1yfl0TPiR8/MzlwixLfSBS9k8LeRo9ODzsiRiyW4sB/lsQStl7vRs/dPrfgYPeAbN+cqCj9m
biICwXalfXuNEr1SYvp8A8fFpfvEXk6icZ3Po8ydIvUEPP0Wysnk6BLKzWy7xsII4ryTjOM4RBaU
/n5Eo9N1RFs9v9B0UTx0vl61/4gOpb9gFRLhooYkndxOMz2HvVace2sj1SRL/ssh+j9kGP8POeoM
5sflAUSf0+UzAIenJ7nQ9knDGaGAAkWCGlfX0FbJ4rAK6smLcymeq1/D6TKugCBTxCmlHXxJpgH0
iU3mxEhjNG4mylcKNYdOF2tMmNyz+xZXIYoWG5DqTxbYqEjxw5vYoSpeZvuU3Oq8TN46ROjIrczn
bNcKFoZaxek53h1MD29K5oIhg4d/pFeJ/lO6lBAfOeBsiYFVZqkJhTuguSTFlG+A5rizg0bqfVEx
WOyKIa19Jmk+a3T7iO+Hs2dOJbg9wPW525tAstJE5Ww36j1osvxX4q745rR+lcrQMGzv3XH7lAqP
HJ/rguULu9Vism+SQQgjkMoAOtoIXjg3okM4qN10vXiSovP/jFqIM/JHJCkKVMeWuXTWEzX2cf8r
odfVJvlnxKn3LMDJLNDccoZ1XRZJGlxLCNPN8KxMIBPsONQUQnWrKd2V8qOGc6vhdXQO93yDj03v
eUtV3PRpVc1rT0iJZHr1s1F3T3UsJJKe8iJTkTnJvFD355JXQw0zR046vE4VWJ4uEHdQgRQcXNn1
y7iJ7RsInL0WK0UwOP+Q9AUpZX3H7zOAM8N66c0t8lkY/pF9tUWLA/jGUf9Cd+vTRXeQzHxrWUhY
cbB7wnrh4KcvA3ZQHLk2UP8cUqtIDfRxnQ0yB+yFJEzfmWrg6ghPB4oDmC6fMDKBxcmOIxZHLPhC
zMjngjmdRkpyyyKEFvqFkQrcRmbbE1gOsztLDrcFmDHWiGhmXjmRcDAjgcu9PCBUwS8BHu+3S/fm
yac6SZIRan/TghindFolEXrWoz/fkoqne0VXT1C39moiz9YYNz6oIQB5NlOZdSJ7XJbVn0vJpmqE
kNQVPnAhKtIehC0/u+F8sTcvKGA2vX1yrSU+afcF/FDo4sXgtIMHjSG3I2n3TnDiFopBXI1IJnWv
cXoix09H8WT7xiSQO1DEJsX9cOUXTOt3zt1syyPM9S8ZG7z+XQUjsZdpnZQ0TqzXmXGBPfr/8zsJ
1hHi7l84AdluLCz01PmWQZIduFzhBz5/yuZ0370Er4jQyckhC5IkG85Zp7AhuI4lQAV5q6NKxKZx
Px9aS46Je4j8FgFLexHCKpT9niD7OAFrfJN6LxBwE/2QlvDCbrEOKIrNPR5WTOta+6rkxPII/Yqy
rpJWwv7/qADAa8da4LUsLQ3e/BHsk0stDawIbXBwknqhlP8okA7tqDRSK7mwtXSoyFfuij3z0y8b
nakbrNeBl91B2fzyK2zzRKontAL9PH+vCwIXKhQ+CbeLg8a22HNlHfzczEkUjs8FwalAM8L+d+49
9hSaNCm9f2h5YQgPZvF7EIiCmZUuWUyJPunulcw2zit1yuktBg5zYyMHD6bDZduEnKwAJb4defR4
1pZhRM/RfmcrNBbfYnFWtp97eRCYxjtMIBgepNAKMTnHtasvCQ1fNoR3rUbZcV04zXkVhbltq0cB
93ZuQHtHE/Ctos0JTCjw3+S4T+k/9QJSwDGOPQ9Jk6nUwc0jSmZ/jaUObRS1waE2oXpnhG6J0cZT
J0sLhjzIy4lxrMOElT6p32AXYZk30RLbCWCyYeuzevlLUpf0YyxoBdmagWZPT84afw9PipTgXdfe
eTLshpS3L3LL571lKV9QZKDbiCb7VDXgm/oB2YvavT81G8n4BWbAvzPxWkzFqaF+F/L8gjmW3tN4
6ixxAtk4S19ZjUUUahx7aSzMG2ygfcoojCGxJBsepWamRMVR12bheqwdrtcVPKoond0xm/9bI+PI
/mcWi0thrZIXR6WIRnVeEAb8JQK2BjyubY/nHszJI75UITx3hX40hjk6qc/zIvNPtEeivl22TyHu
BKNzUj9TIZSSH/Nt12wL9Af26cgNFF6DYMabvEC26SuCnOPsIDmdquGdKQRkRB0IlhhMorR0Ao9N
0hQ0rzjgoq+tZcUf4o+J2TneXMf/bDYDLait0PsSM0GR7N3bBZGrShlaXVcDXNEbryczqi1L1hT4
YXINcj86O+izluB5w+odI4UztoAMlYn+usg6wz6T07Pr5rdDqxSwYgbCYUhIhZS35Vjl0KckI2Ct
OIHp4TQdBwVIb6/vxbOAlQIReYbRcNzTrxa7HMQgdI5OUbfqY9Rs/tagb3CVJF2xaYPB8Eco8JtU
FmuGwV94BxanyeRKqOkaSxNaqOnoDXlkABqLpT/sw1aDIYdsMUof+8H9E6vX/RA8CGNF9AlW4Bwd
xwLiscB49xbO4kPXpgPBX2vm4vfqV0mPB1cj3mk/qt9WDitmnP562uaKkThF7zyBiwanyHO/L/lf
qwsV4C21rXl3A5AFbGiua630xbvlLnH5Dh8Sn6RE3shzaguzSxdy6Vcms0K7Opv3BiW/mFmd25qR
djOHeN4asenLULX1Zo7ABZ3o6JtA3u/EaqtTDGOblaKHsnzutb+y5lGeXr6/xxbrzUJ0WfRl1CDw
Lr3KUtNOSnLwC0DpGYRYSO5IshccYRfI7Oy53YJOQQk759cOO6O5hzBL8WPuLSogZIPJPUc03fb+
SYo08oV5352Tjnhyvj48tpmsIw7ZNJHtUVDlO+zZBHlnEb50gUEOg2YuHzDfBNxhvASyAhGWMAjL
tT5dX2pdcRUImmRjmqZ5Ymhr9drAi+aTqK/BaSv7nQbf/IKzQtI8WXbIsIwCCQGshamXbqTVdEyd
Gjt3k42BOGdRWDBwOVhPNgMBDeu9v30ZMFEQ4MCMrCA753cyFYFPVYBzhmvh5uEYT9UOlo8rsTeo
H07RJQKSfnTPeLusWJQ2L01CxeFxiOyQh2XhkPmEjO+fzRPXnC4mkvpVOXizA7Vrbb3OojYFu301
83Pbp8f/YsN+Ik3VgTiGHtGtAmkISq0hFX25Qp+0PtAy9jy/FprUJEp+KCU8nPu/Crxov4KqHsr3
TsDa0RF23x2eqLOzbJLo2QHeE6Z8yJyGNPsDbNAmwkkBvczEtEA0/G8ItEOdqzNsNdAM15bPtHpN
JTA82SNoZk8agPgDv++w6ULEYHvqiZSvCHd/Wh5Yf2m8iGLEg9PYZC667WwGXSZTNtdm3LK/dgqH
+Kgwv783LAprtOSke/7d1RBbWeY/eCM2pLswzNyg8Or8mXHJ7t3/OFo1lFgN7uEUHybhBQhshSfa
zisCy+7CpScXaUKfnjk9uWdod/+9Ere3N888SkqZFCp3yT0d4S6ChvjHksXrIF7zUD74Fo3Z9a01
aq1wAA0b3rkzYmRKALsIbG/0swhA9ShDA8ntHVmuQv0l8dWegxPJ7oAFT84uOIvgrR74aGOfkDeF
A0JyM8YnGirpYLRN7zfLKlV+HmYaHn67t7qLXR8sIPiaSECNICjJN7UAfceQH+j+O9OgTErOuIIw
6vE2710oAFqcdXXh/pH9u+o7edDI6mYE66gbgd1J5dz8dqcThPYjZ5VfI2FYzPwcLXW8TsnU9UVH
CqtnK03FqBUsQ/Y0keMB16ZAAApQ3RTpsjkqBn3gzL/D+7wBfOBcOR+lYWpJZtmqaAzJXYetEg5A
V4JdmCc5ssLLooFntqIUoYHivFeteJPKrf4Vr37bG3+pO7r0UDBKfx7THRvox7uB2iWjOxebbDIr
fO4DHOTNo15rwV2gI8jBUn5o/pgdnmahtym3+eB3V567tGKW6ZEQkguQX6qHrQsOhDsSvCGrnqxL
keTtkgvjn4tr8QvGD1Y4wjYeqcyTz4pSOsng0UfWu7/rcRJjEziKoraXnFbOdRASMYN05xAQj+c7
jjHGiZtHNp2+m2Vf91Xno5pyjGNbp+HxzZE4J9dcY65szWm3yFn6imLZ4MeaxYK9ERHXOE1dg9wh
+UITiJxnLK4kc4T00yZlsEFDO+M48+DxbKJuho63HjKFLv9ZwX1vs38C7Kj/kYhUKdRO3L3xTCmU
Ta3kfHjEe7Q5gzqqmmWKixd6RZvrnKZUATbjAvfy+Zpzg09pk4vtaeNA/whUpOVBtBguCzZLgtax
iuGgYSa/cOjjiAl+PSrpgMhuCGciy9RTbBVJlp78jYhQEJeFaV8gBuIRtI0OfRICJiWjpULgQkdK
zWQZQu4yNgJa7961O2m0OCSjQWUgZPhc7WBhnJAVpZsg9a6Ub72OEJ7EwcluhANpsNOLMwu3RvKX
/rRy1KqAem7qPZN25eC9Vj9zN7YfMDblm+j7gWZbck4WG5hcDLSIgVKhU5WnU949VWf/XnwcWSCY
Pw2CzY9hTngqvtv1okuYGB8nvU5kfbSl3WLh6WbHTY3Q2rXAKfk3nuxPVnxeqK5hgAIu/HjkiKzS
9N8SbxhLXHKgcUaXjArcNm4o+VP9YfGC8l8Ip5cy8KNJRKh9Zd09D5409Ovm1YQGWQN6rBK/9+xR
sEdD1i9EWrjTFo/IZZ8TIxAy52468c5QyTiRAXek40oH/9O6mP9Dyh7Ug4EpJ3LyDPZmAPJS8CDu
nyzLajThA2Xs30dQ4pc9KNlGeo78OTiOOa8eR+dNOOpzu8THdhDQbXj7EzNzPghm1k/nPyYj8Hgs
gUrN6vLTJmk4EOFl1JDMCGeAfS3WCfYRPCPcPuOOriduCNwwNaz//aopbSukykICwQIYRQN9dkat
gCLBxeAp7fbGGK8yDGM3GJoMBVhR4BR2PJZfPPw2vmjrLrWp12jzsZK0/fNvX8w6+z0fy8spOxjm
08SHHCqbKlCHoZrbw7TZJHp6M3lv7qvKaeDvrXN+8ouZaNpBaRf/sJFhDkBmQYOnjBsa1LFzePWq
NYM8cArBJF7HzeBexmHyAtSC8HPEIq5OGrJ3WHnrShNH76nQCHINmxPnbcz7RbXEODtwr9GRFuxK
M3xunPNh2U55kW7+AqrO3vxY0yW0o0miRTBIqQFO0JZzdVtEjc5EnEcZA9f8hOVV7UdA0G8vIijS
BcTeNHBURIyFZ4UCndBkh1x0OCT1KQ8i5d4qBTiPVMJE0Ccr323WPchlTFY8aEQywnYTQupwe4jR
VjeDORoCngKOqX83ORWUv8/5bbV9XiTgO0/C1pN8W/xQdLCBS0uKx5vi0NAdfdA4MdX4bt9tEwgE
hxkEkmdcVKQBFsoDW687+yvr9TXD7uoqQy+p2HRbqmqjnc9/fQ7c8mWNAY6Yk48WZ4fDIRTiddO+
zJ/iILBlSLmDmFPnVfRUVzs/sbktqcdBj+iS0ka5zsqbzGQQl0K/UMOdYFEQpZXykBodEX6rcHFc
N+IAUI+fb3vWEF9pgyrJFkGkUByWGtBe5xxSnO6j87GSkBqmGO+5NZo37sdppP+Yjm28KewB+w3C
pdRu2+oGpEpn7qYAkGN1KI4z40L1i4gt0hpnMIfWO/bK1Zon33iQtNdLYHD+H4Dx/3m9WouPbiMu
Y1R7YFfzqSMabv0NHKHVU/bvGc5CLYjO+Duq8vg4trhIXOa+Sr/7j8XRh6vDAFWARtU2YCTJrwDZ
smzs+qQTurmd2eW5giPF6ksGQQoKQMD7XEu8h5XB2ACMXD2un7mVf2Ji40kzt4raeVr3Pu/E7DYo
YJM3woDmcJmZS4eo83pZBHNzTAORmXFOHi68eXPa4S2UXJDD7sBkDBz02VrzGPabfvxA1gBfLp6m
j2OH9LTMHOQr/I1Rif+L6EB3mY5BjZUQtUbVJV2Qp6doyWb+I6Q0ezzmy5PXNeqWT3vMXtr8FV7N
5teUOute+OiCV2OviyDwvJSq8Mxg6IgHFtHBMdpHjaEUfCWVwezd+S3AxouVSlgLOP5bZxlIrI1u
7tHKnT4a3tCthjlLsfrPAecVzT9ScK2PvK0zgJq2CHGznzS4UN7NzqrmAi1vXfTxIddZqjLeIdKA
yApVZ8KwX6JuVN6XETqhP/rCUHtk0m6s8XAs1yiRVM3xnBFXhfw8rRkFD4SIpENz7R+9lkWtHMWp
m7bp/30zxjqifFO/NlJJm1WfffUkmLJgRHoIzOZsPx+uFk0c9DgBH5fmdf4yahtXvrYL0ecZujHO
JQ8xzHf/ueRob292DWmFqOsNPi+SvRnIRMn1HA5QiYurvUR2kFOy1cmpB1aCp/0pr0pR8i3NQ9fv
oxaxuoB38fdohf/NICbN8AG8eAIQD0RKOiDgdV4ZUT7A+jyTiyGyN3cMEGkvzmHIbJbYTJKhgsaf
ur/McHAmSG5ceBHNSDNPRJPD3IyMTl5n/zFoxLWbpNq03+cJt7zz5Gx2veAS9vkeGoYRNC3WOAtj
qgMkYqvyLS2+NstX4+COxakNyIli5SCRyCKW11taPrtp9SMKAwPGLTxwjfAggeo2nRwdOC5/cuAj
nikdOykPisUxdXmJmvo7PAXcuXNgBY6BqIwyzonFd1JcP6hgKeMymkXGmqGHmMqUdHXwZvfMHEOR
QjrCSvFLXnvKxXkpQYbSX3sRrvgExB0sIwKlOawxkLgJ6X10YzaEbK0vMuC6/TNd+Aq0cfPHUrtW
sxUoFj+bcBtIMf+It/tzHH/HG9SD6HJFcWFB8AMIs7wjtb5v3pYyjGuweuWvKjI7BWL3MxSvmeLj
7DUuX4mS/7vzqvp2O6vACAAxjE+JWMhntwcv1XL5lj525HGDuC+8geP2SJMoRAzAVIWeZijJKaTf
lXlyMIyFMfbiHOZIsV8RH/cqRjqe5FGWSKsxg+0/QL+LkmCF2OOI7cl7kl72PB1SvhbfKeeq4MdG
+fok8oQGssEthcK6T2ovbMf4UoAkGRQLPYFmv02AJ5J3smqAX5WHSQZzZwWKiHwAv6ydKRTVq7V7
y+JEypipt0fqfTr9+5nRM7mnH+FnlHnpLOgaF/y28xO9231GeT4JDeH7NQXHS7N44UukeO6OD+tK
QDzsFAdkzPgh07a6lqJV7mP6SIzkVWkk5reIvlFmVq7j1AJYpQ2MnrxX6D6rR0X+WF+T/8Aabr+B
BHyWEvujNNwiW9GMfcjZAhAHqgCYkprve1Mx8iaohh4WeEJcDGFrGXHP/nZT11/sl3kC3fR/Ebay
CSR7aNbJSXesalFVWVHbEEjrAW+c+0aH9HOKPbx4wxfVmMQJ1dImasJwGcDku0X0pwpnqAahf6Eg
EujhVS7rWNrJAb/XJljSfYytJDs1ohe9u0dxIr307WW75GGN2FxWTAJTeOGJjIyIHHOk7sl3KXGI
j0mCUR37Xg9WjFtnc7Rl6dgM8zqWNLu0IzkL1tktaEa7a0KJgVrxXSRFWoiLHkdNXnqXmBYC0INH
k0pWw9/MpTzS/f/V09QJQ4hTHqibctCVIaAFWGevI1bfSrSUZX2CyCa3o4ySgzbzMi1XrGKXkzVL
H1Knv78YthUqilP/NUa5HvXUJKa43yj96p2Jj8Pvp2HF3vk/ORwQ6XYbdPU0ZvY3LSALszuD3dxW
22F+iL3AF66clXsYGe5DMD7s2xq8jcw+whXfTZl5wG/Il9XSGL9cCf7EhuKBc2lWhjD66KC9pgVs
DeYwIcncaar1I7tRBp2siNB7RFLK+839fMBzAnQJxngIWY60KHCUV18cjHP1xJT/WGpBXkn5yZ88
KDOZmKyVQyhQUOFZDYTrFR9zfmDWlcffSSfsZIfY8vRao6gF2Xp2yvgF4qimkn1B3Avum6J9Czv+
QxgnTwDBEMu0lTzzA1ydNdUfHnlT7KjTSAtMQdEd+SFsCjbDmGFCClv6hlneF7qDIF3XFHjpGTGj
Iy0f6RHN8niZKSbX8nUPAm3NZj7nXjcyK+OC/ab87/ZBq6rc1fxF4VyNcpUuDoyl7l9Pp8Sv0klM
mylxmj2pzycVclT6Iqfs069k+HZ7/x3HNMTUHE+FyvDxaqaZgE5VS6HIf75iuR197qn/R360m7fg
VBM+AFERzHqLFjkiG5WngJiRg3XsnIdWwmsQHzmrmZisi9lI0XvIQ8DyD/DtuOeqDO8cv8GZUUTs
tV3NoQYPc5t9duZec1XzECSKf82o44t40Y4t4X6dzHVFOTTRk3zQwTitpGZrnA0zM+e00ZWZ0Atd
ryVnb0yxIbcUGs7ery0BjbmxabbHgSnW2uzIkJe5jdkhmv+j2jnONia61rrcvaTjSAWEgPRiDDlD
DiXjkiSH4Z7htB5x9QrsxKpciYNG2bBjobWQlVwjMc7HXzQFEow6JNc2jVhNzi/HEAtn8Dq5vedB
3JoxnkQZut6d0wpWQOIqdYsGaKMRj94GgOqVn/0rNfYLuzgt4wakF10fxMWXFtmfQuIX9vCf49HE
BcGxHUnm09FtYOwJs11LEzWoaXKG6O3k3x7K4DB52QEw5N5BSdRkBYdUqKtbGIqBT6lEwV/VPda1
6R3zNxt2nmtE+aNOnSpxkq65C7IWdXkGAb77BJwA9Ko50QOcFEs3pRHvCn90vMLg7KmSW4KtbUsq
Ip+ZDUPQxC0muZEvCgk9dS6V3ceUS7b6yM7OcwZIvRYUs1v3WADxOkwY6jxQYG3Rbyskgb7zxkni
hOtcnUlgnqy3TgDrWwgQa1WKjfwGUO4eoaiiiA8sTOWlcaZit0bH7iUEqq+Ee9IcwMKOk6VnoZf1
22/HHoWlsjfxNbWIj7TRmYmhlhkr2Tnrm27wR91adgqLYGZBHiLVtTSEQU2ujp+3i204rlj68pe9
3OClw1+ifD8CSy2G9hL4vj1n2VY46j6ryLLH9L1MEodHKR64BsD+TXkckYgF1t2+3B0hzf4IuzEL
KBovdjDSAl+hKVYuw7KTlK80k8kaleApxZiDPjnDiXjMnijG8sHxjMVhlRSRoHB+3l7VP8NQLYEp
HBTW7g3gJVZ6ZILh+TnNVYj1n3qaEp0repCPsBBVyG+VAgbAUp9vYB6x2VqLxV1MErHhTFtxCDNI
XzBOJTPEhLk3S3mFNYuP0aBETdypuIYELJTQspLpS9HGFcA+x+T+S0cNbAvifERF1zpaUuUOOKEf
j1ZF10jotIotV1XW5ivHEYBbBnL88nsob4EL9HWkp30cpmNiK/YSBmA9+/p6EXQ1arnUH698bxla
OHvSRdVPR1gAbOgb7jiXgd3GotQlwGhfGGoyn6QtkAWuTZAfz7IV/164shsn/PpU4bbrH4uubGeq
z5TE3OHhYUUFD3u1ve40UoMfQSMvM6O2bZwXg3JrGABEJHDvbBRf0A8xL4ps0pz+wW4ApkaGWzvO
7pGWzZKztFfVu7c80FGlCcG6U7kHQ20UDtCbVt7cO8w8pDt0b6xx/w8Jm8pe2n2TV5hki+njNuje
nh9BzSb5ncLbZu3WztypuOPzi5jOgGGctsGjDnCYEBiXbG+3UxAMS7zxq8cI2H7V0kVJ3kqpKKpW
QfyE7x8wsyv2RPVSmeq4q2v0e6k164vf35GRYd2yewRqd873yfl6ZVAhiL3oeJHdFgwa+FvgePB5
bhSfTZfILj/WYhp/BCP7DArsZMaYEx3b+dWnuH51bbAdZa9lMa7hEU78OPGcHIlFXkPovhWFYrMW
M2J2jU8/BmsF2C8vARGE1qJOxE5P4oNdw8uKxje7OAWtKglbdDVWAaZ3++o258zRu8KVXIrDZEV1
o+BZsLnL/BxJ5o7WIHtVIYnQ7ZyoA+VUwZxxFdULuz7l1PHNvIOHJ9Q4snDeQ/s5Yi1B2TE5yca5
1+KIa+eqxypOnTLK9hWID/w7N8kTInAEkdcQJ30dT2O9GVxazk9h/aWrsoyZEmOVlJri/imk0bO1
47Bw+msP5t05qvrpZb5HbKzEhrs7W5l2u0dr+wvG6lX/DwgpyWYm50yUW+tth4lu3kBwC+l5yt4h
D91KlF8LJrahnR5BzumTudNMxlqVM1uycfTKNrRXP2SU0sT0SL93JK4ZLlh5AnRahdl12tejbnHr
zVWwpDklqzgZszqFTC9nn0+quBdWgOv5HzUo1H4ZrjAXULBuoBimBCCLiMXfZrQxWFPz2sBeh8T0
0rPFV4LohlJEW1b3kQNcjQeqTIidWmQPKGZNfprHE+fSD8qOBDiw7Cv5+jWbXSM/DnUmZhpjG4U+
Vx/nI0jdwaN8teVcUW4SG1pKtAExpA9XQgOsjdGaVfGb2f4vzdCTNG4cUOWLKFZ/prQhJMPM69GP
SFs5KnkwxWTlVfdrNMbE6tU3CMNK5R0L95OzIEo8qAStDzb1ddEQiRJjXVGEih7lt/gQZagrzlYG
CZUNCKUaGdlXU2wpp6dTHvh0B02xJKh/a9NLqdKvDlwlk54tnY1UXp+nCKy3NDqkU41aKj942ZUV
8JKrnAIf2XWcWmi7xGoC9TmrVgax+rCjF2glQ1sSm1WWqv/MduUAu8u+maN6vN0KnEpjPpKg/MqH
9TY4jiGvJKgFXVhZDKqLLroq1zaKThUQHb9dQ4CTvmxAtWOTHs1+Mg3ZmParrKakea9MUSI2gEOI
4ZpfMGtTixjpL+0LUUwBPebyyuuRI/aH9/vvK8lkmCwgPCQLTWmqY02ESHE78CHxql13a7hrqT7/
RcAJ4HVUXIw/0S33fbeOcAV8pnDhiR/HwNGBZvXy2ttexFbB5I0FX5wu/AakzRurfps5VOau0BL6
c675izkBtHPyCvELtyeeB0HRKeGucIg2vsPWMgxx7pRKy7uI0XW1jRKH7F7bYfyUGLC9To2ha22+
5UQjBrzAll4qeo+b4B/NfuP/ynK4DfHMt6N9BTLqeHCsCNuQCrJ1LVSmqrpSjWVeAZIOSwgw+YAb
YiytCajxhuJpXXLB6oNB5s1OJs0795pnseNbw9ZBtq1noHC3/+X9gfWn1JNI7ai2Oxl+/pqg/zzg
7yI+M8LVmPLaO0WMj6MdcrrMR19/rzXlpKJt6bcvpP2q0TWb/PeQ37jPQbC/jouivXLwMXU4Ak8A
4lcDCmKPQFW8hTPQU3C0iPwhxWySJLkABBvoSJXliFL5HduDf0E8AihptekbOe5LOW8SOIlfOAF/
WYC0HUY34/5rGIdkT8i/ng2COS5x8UyBhebLZ7NyjrD9TU02dMRvkG9QlW4HbNbD5Lw93rpwNMg7
+11UC27SBIeBzoy8VV8OyF6bu9jJsjy3gR1rmLot6FIhr/U5HcFj2KBMql0R43hhI9wade9YrrP/
836KA5dj7heT0r46HaJdFnN6C6oo4x2DwULJoU5NFiea/AytttIlN1NhXjNBRSmGG5RVE45Loiyg
5e607jQIbisavAIZ4mP7Anl327B30XgjwoANgolw4/Lgy7fGJYnrobfr0jgyedewYCSAwMigSpRA
7ezzQaXASUJ/CjtJOe70+N8viV3LK1jxrne1ak9B9q49LUMQnqVZhTY6OwUS2vQNko7p+qDsFzkn
1eGPUPVJ4Gu41NMP5yzSCn35kcKkWP5+x5NJfOikbjNFEVRkU7Oe34MWCyh/kz4JUOX5PURftnKz
aM6ZC+Q7DgX1BWI6qYDkY5QczNYrdDbMOFsowwWmbmo/I9gERmtOB+Rm0//psh3BuCQLv3S63soV
ZDjmolXHAPZkswdnzG1S2KCzg5lhUmED5FqC8fIVMR46jl+oJVHiyFf6kKpHQH0/uw3tALnFVagJ
xtSyQXHCIlRQUWWq0162vZpe1s+ydlgihL+t23pdusKPsvzOrxPxbAnNV6ydB5O6IYnCJNLLAYZK
xDevpi4gUf7LVjBW0YfNsebl8xu4PWPPzp7BYRD4lHfszuC8eM3T9Zqynry52C7f+S4I7JTlRZXT
JUs1tTUrOYxwBwDEHz/WlSLYHRXeVMVBjSdZcmRP7XRaH8wysjCSxMq5GZW4cI05CHNtN8q+vmfS
3HyLqegzkZAR3qX7KkmqZJ9EHJYJidRiTlEnlFWBzwTsmqNma/nEqXe+ka0vvOdxC8Qz63f2QtFH
IS4bMPuQP63/95lCxzNMSRBL44P3WQ/QMac2MseSLy2rxzHJa/so8loSf6uWhJj1+21Fok9FOYVy
xbgBlx9QnQo/AnTFJ+kiYW18XudE6hHrnPVe6tJrLhQKpMfosAu3SV547hbTlnKoKf1VFIziBIB6
f7Jzx7JfWkRXVqvaw6BrNmWFCXMG4Pz1DfuFpkTP+v6R37Sp4t32wzr5gGfsf13VOo7gi2lJ1TX4
tTyV9/MPFvQT1Py1b8Jr7zUBbgtAG4FGKd066mFYpQgjvwsQHSovBoUqlz+un5dKuEfz95eEodtp
ARncYiSsaSkg51mDfPhhmERjYsH1JZPxjFJ975OayGEJSlJMgSv7eiS3wKNdAwX88x9ciFANz6zk
yZDI6CwEeuPSFdg9Vs6YBUpdzY0XIFwbTQD6yBMgvbWiigU5WwS+pmT4rIGWNAQ7dgOCM/9mUK1f
JZO1d1hd3xvZ2J6HZJfYdK2p3qfrXQquwgLys7ST4Hrno6kSxFE4KIecQl9ipr5BkSiAfNQZHxMn
D+gSQo10Nkt4HvAdVT+nfwntJL9bqRqG9rPSwXPYW70dHJct78rj94oJnf3qL801ETqFYMMSmUCW
ytNBqnmD28pKyE0PT3DBUENiWzQ1xeM6+gfd6d019MZf6AHXzjckjHA9dP+eChhb1m0VRh5NYavg
X4Bz4cCF7AOxTYc/bl1bv5ep78HC4LMmBivCoofvkgzbtmK50EhARq2YnpkffzzzE68166xd3wtb
HnLr3rNYvA0fn6utc8q+yKXKTnt53GICijWuPgrE6YOIAjrxU2r7LAyZcqNc2WKb2L/hYknmWkLm
ibNmKD1/tL0JJTd3IYMdU10L/K3ZNX7OgoTKfHep8nwfeVHLmi53N6eY4TYqC1l4fkILLjSGLuDM
5S0GpIOZTAjhhFR7v17nkYha6qjOk9TipbCqr/MJYm8Q6ZmzgOK1gRddf0IORico9uAo7GvSZwtn
STTmNJ0FkBjY9UdiDyXXt82LxH4RyI4Ut0yM28qafkWpw3vXKSjykqrEae2TQojvKnLJl+XsIGHB
nuuRvPxkdIju9m0WVqgDXUYrsBwf1MPj5AHt4l1u9SRludAvBzlwkkHDidlLFtj5joO5H1WfZ6XW
CAuuvbZAiMEYykUtU7vviDtw6YdkOpBJI1VFYhWkevnjckStyBl/zM12BnbkGEBl6sovqqtezCtW
8v19t44j+3f0/+7urcK38mzdi1IafEWZj5qLzBWIfn6RlXTX4b4gMJnTOZTwVEpoBOUCtfpOl9lM
vSPxF4TSgBD6Hgxs02JidXhVCjaruEuF8WJDgn/eWVMgMtmlKcC1mEKspUahewFLHy83ksuL07od
DeEztbTsMN2NN7xNSJ82q47LcDpY/IgSkXETxDNfiMTeo/7wA/x/VfKUEkIOaGVYuyZM9FbvzkE1
Y00gBWQqxpXZVdKNbVj67x37g+jI7Ob2omT9IE+LbOcydhHpUEVXQWOgAphepAlj/bIjThjLC0GY
lyE5jl4B8K/b3cK7a/zEPg7ToRT9je22XF4yB6O4oO65TYwHKt/q4hXZNW1BT+LEVwTEt+57B4S6
zUNZzY4mkoP3HrqOxJ4tqTDIESeyNI3kDcXZiVxSAhstsz1ShbdlOS2PYO/ujHQlr0y7WugcKlvG
dR9ymVzEMcxrdnNescrzychXx0jjMXA+aFWE2KNHugWwnXvvbfAQgeDhGPG/eBnT0NFuf9zdvAV5
PCpnLUQ3XeHnALFSnlC88yoO7BMNHtK7rEoptfFjEy5MfEz5CFiZpD8sWfQjcFV+DMKtMYA6K+ba
mMl6JWSk5snxt06cKbCrg932ZtboWRjvZjaz6Ei1zx+8/12Mi73UwCRTCezoMs49Z0A9IFHzh1IN
yK8uKgey+PVFKKUp218XbRAMONFkprYGNbYICT54sKOrAxrTp5F3lDUZDpNQ/HS2KFhqxYmBpWRK
3p9VTwjPo0ZsX4Q5Ear4Ph/eumrPjTfRFjFgwJLCNTZ9RISrcrzesu8FE8Ztb+vUzZzCKVFop+Q7
axJNLkvoCMYDfMhjUCLPKR0bFSkCtST5CLBbxuG+NN7QbdGsz28YHCDi8SA7j8aMmK+O5tIdheEc
MZnHIC/QXFMQebtTS4IyQpGb1ykPaaX8HKeo5wE/IWpAYEOlImuHutkAdiYMSReG1Q4mcnN4CtWc
0HsD3BuZgvwEziCbJFfVBGboirIo3mCKId5AMR76kAyuom/T93FA020m8cvRMn/VbtH4R5d4kNJm
P9lvbDtcbA6sm0XeU7FN85RUhtVubwGmyzpW0XEccdbO2azMl3OOOGVrNNxuHddPdAkuRItGKoYW
96xu88KbE2MeJdsB2OAx9r+uGTxWPE4JVTBk8dU54w5ime2kCtFxPrFgSPiuHoNVaLD6p9aKgl93
l3BecxvIookTOS4Dn7CyV7nO0ptMyN45FrvuTFnFqw6DDRCCOJswW+GXNJBq8SjFlIeUOXrL0Gra
KMZB3I8MfAhYeMG420ghtk9MgAjDyr1BO2Uu4wLK8cRD327aXGnsLchowdffe0wPNXQUIO1pedzO
xaKra2ivS1G1SBiUT8NN9xmk89Q4b3u14EnuxkfXjI07W037oUhSuJf6tXn26nLXSdQkpvr0iBaT
0D6P5pANwcNVdFtoKj0J3+06fnoiwU/shJHX1Badc9KejL9D6CdgbTk9iWLUXoM/1NwfSr7E5Pz/
VrAMeKZuBnZAZN3nOzA9MKmsTrswPUEXp8BmtUAxW4Ja8VwyKluJsA/JzO9AVrZvZR3/5ruoDjww
EkX1iYwIH6MniFQCPaeujXHFY7zi9VTWVRKdwTcDnhJAkTEtI/QaWVDn/C3LFP3N3oeWO6ujFKBQ
DzzeIcLFy3ztcFZS8t1I1sxMayGPJdQFcQ4PF3X9WPTyFoTtMDPB1onAsdsLn9CtWFB3sHewA9gk
PBdvI366fQvaYkSIoIxnb7g7b2ZaAhkAnEO9YOqTSDtFrkGGKRHOmrQu45bmb8gn441GNvEbFE6x
ITtDem97EWEOZhobJa/odRl3x2dkZ6fSWySScKAlE7EOPVchnrbtb4j0hYRrJHnTjoL2Wgo/3umq
F3dG23rGRo7wGnx3H3I2TbN0v1uzsMHFlAPh7Xb734+7t3gYAi5qlQDVGWprtWyY0Gs/TELCpOdz
/pA0Usv+Q0qqHH6sDRQUOAUzVSaGTO6I2Yq57/scTmjsM6pIn1lEeIpt/pV8IhGkE3K7NHTkLAso
s/JXnuIuwxokpeRHqzPpjNajutNHhitjurnd2wCUREJfAtAFTr6Yc/ExMNmyd2nA2U7UASZ1rh9m
tec/QAwRJ/495rjD5YbgypCzw5imwppBWWHSC6iG+ALcPesS0oU7uZYYBKk4xvwXeooNu57UTGlL
rwMFZm8G9xxh0C+lHhRW11Efh3wJF1KKEQiI3l1oBz+B5Jgu7PPyZu+quE4Nf+RytGs6O9nZrxPd
sosXsIwLtCCp2/xleaZbgE+vkyUSVfyAtcyEwbz2kFh29fUj6O0vldbFo2EufTzK1sDZjt07YH4V
s2bHVR2hPmcjlQBvgIA5OqbQk4HdbaohbIqPuw+QKi7IugAitOKv6OUMNhxD5SBpQ81SbXlptqqH
esXkZojf4/Bd88Wp1zmxu3La2uTePmhOHqSMliXEcijIujxxrC54vgM2WE5OjxzuFvUXV7188+rw
E2oahW4n4ECjJ5cem2Jm2JX5rw1lU9X1lM3Ghejgm600iJ4htwponbXNzlnctGkmjO+yFpLI5irH
p7Yq6QGgTHTJOx/czXxcRq83ZL76N0PniEisHwi8DBXXPFhXIrAdV3ThCA8qKgslB9PNvTw8N7Si
C6ZD3xMs4BnAqMSpjW0GxY8nT79iKf7RnXSLoUgZ+4qA1iWNxNstuMYCAWgyliYarQJuLxehE/B8
CQLMikP6kIHZFCDFGYymwIAeVxlay6JD94GXQjcRgLuCE2usMLoFSZypbtCJjFnLWSNQvgX6A6Ld
cPHJO374/MSAK+vxEJWrGNuwLt0yDFYN7SAO2KukXUozyhFTcsgwxaZ6DIu6DFJBKBmpiw9taeCT
/rPxiWbBkAidqditBBeO/UAVcVtn1vlPiRFCT95RK8aK3rFBU2ZOnJ0B/knij7kBAfV4th2TKDV9
aqX2Uo7m2HVsB1Badczk690IoCedIVkWqDwrXbcUp3m2/FzdOZR9NOk1GUVzIqPsPibZ/+h6uXUn
x1sA8tiV4KD94sXQg5n7fp419tDxDg3ZdSf3R/nS0z5gLYrOjjzhw59nz2RSIYfo5llIs0yui9ee
6QtagzUbkdJi7ooetI62nQ7LKzKm/0ry0P9rOppj+q9//ktcvFLXsoTzkUCZHuTbT8zQqsuu0KcJ
vryhYBL+9GHJ1GEWnyMitfOJ1ms0iynpcvUATBgNbJoxD94OSdgD/iWNYaTrTTqvoIlGm6dgXaHs
+N8Ado4JCUEexetTSIfEOpQzOhnXh0O28c8U/A+p4LhyrU6ClyjoXUYbVGijAH6caJWb6L5SuaS5
lntqUSqy8RzS+cjaco/yzJsVqDuynbzzQolTQOJjLmCBq0j49UVRThN3pgJg6e2FCdoomo1y1vGc
dhZ+NIN4uGOGfsUOJrjN5ZExbbeZ9hTnJ/zNYKMqSwZ9AxBOsIOZx9+oT+8dkI1SdpreA69lzk5e
DtT5DzZm3THOWr8Qi7oQe4350CIo1TEkYKb2Wc/bZ55lIhXDDj2HZYVlpLPl0hAk+wwMz2xY7cgn
OXOsCA82vis84XQlq2+pharf3rkB5BKp6h9cS2cS4wTzAwAfWwLvElhghwjdnMIxqZ5g2Hv/dYTX
rA6cr1QM48wH4pRGVCfKUmkEJh1Ro8UqZisF5ulueCQKViCkbBJkM8OaNI6wMl3+NL+ntH+eBvhk
pDsx3GqzASNtOll3w0XasewdtApMq2IZWQBX0ZUhGxJtM8XcTZPnvBs84CFXE/ME65hfL5URFELc
FkFz7IkgvLzU6o98M+EMKol43U/QO5rgkcWE4QON0biP+IlUyE0FsEvI7zh1ppuNNVDVJThnd1VG
YWbbeEbhi7wKa0dQj4Sv+28JrdmU6jCcU0tO268IgmtNgbz2GRlA5q7HOrOb3206tc3MRqtUXiFb
TErvu1f/myhariQOmuNEX3Cf8InigmTpOOM/JwkcLOp+rh3K0iRWkNq15a/4jO7GBIrQ8GEjfIkB
+8ScME9QWTEFs/BmEFe1Lq1imRC/vDEoQnpL4xOABoTio9/KZiT5G7IZpMPn8RO/BGSPtklvAzl3
0cxB0hVGvudpLoejLnIcgMm81dMBPRfuZeqsFywWKNnWf+B2AtDr8C8bmxo8mqxoVRwzhypvQbp4
BkwM4pHvkhZCJ3mOP9oqFu8GYH1dYcsrS+hW40ysyRX+OyWftyGTiVCiIajf1DW04oULii335Pc/
sPNkD0cTgp6Jaqa6qGMN/3OsdSiD3FCsoPVpJCP8zOtRy3b6nfoNoIa7nKVNMPphj/hpDD6DcLkt
OS1ThKHehCUxfjqUAsBmA33UAv/YVTfJWwD0Yqzr2evNrqB1HW2bSD3YoEauxPxJ55tQBXrFAvgN
Q4sivzprgtzD1d97VJTkkJC468ARMv1yt0uBgVjZgTGqPLYuQ6L7IPgP5yNImtWQnV/2K7Ctvcl1
FkhDRDJxPelbIwEnrnLc+Dk1dZbIycdWfEDm4e1FdFz25tKYb+0U70f9KlP0i83URbu9zpIczi4V
8QVsQFiporagPsYv7Tm7YarrhxdD5CxbQXVSmOQOxEseAk2nk78kRRgga8lvRRW6ZpJk4y1PGvsO
rOvuhB7clnWKQZT/4U/66vrllup/ni8LCDmizEIrTCqFgBSFQLHERCfr1d/GnYuVx5iJnEH5T4Gu
3IMCXUTqtfC33JgnkKgpe5J9tmDb4VS4B1eoImH+4c2SxleEVBSV2N25kWcLY0SYQeQ41mGUCq+C
iWpSwZ9Q7BsFwCLdaf0JFh8dmI/DB401m7LR7raa3Lr7qo6sUeVDPHwnyLOFbJP30pQxqUf8A0Wm
IMjUhsWK29GYIU9XrxOKrEpbHJC0eX22pLc3WmwyrsmCiy+oKbqefzDgrwplNrYYLBlqPBTVzIpE
lmsyuaQBeUuB58jkXZRp2d9J09ZpQgD57kKyZSPR1mGUVfRkq56Jbb3a+Vr1t9CP8yV6aZqVgAFM
/BWY8TdRmdnTYfZxAVx9/azrk1PWUj7G3PkPwv3mi8isE6X3WtgDaY/u6NC+SRoQxj4CGTtHJlcv
Uaq7Xa93LcH7xwf8OMSjNZR3p/U+pN5Q+TqkKU6ihFeyGlCDdxCZD94jhU+Xrjflo0aY3TIb9Siy
eVWl91+tA+JLqkTHJXEZHxWsiG8h5jyrqDW0X9yNeDpGB09R6XHr0JM54y/SLWbkV2DlcRidgej3
8E0095xj4fnJ6eq8g7RW5lQZK616cMR052UZW1rT9d9lBDL4LqFkAmrwKFDaWYftRwOBE0FVLkct
ZibI3TQwIoszIw232KrBYlM9dPFQOzXq6WcS4noq1OPF0chhEQDo/ckvQFCRdVxI6ZM9CgU6f6Ac
rJTvKqMLDRdxh779gxNMz8OTsYKfG5rmr4Zm7eMCOkmroIDl/9ZebKc/A2Oc3vicJ4HQ4eh7Vnyl
d0Fx4sCxUTB5dP4VmK3p+aKigxic3hhnr46XZAJknTFrarWShDq67CKp0ds0DC59HWEbMiCWParo
2kfWYYzed7LaXvQdQzpMI5PWU4BDpRzajyDzwbr5swocH7HxzFOvRKeK8JWuMstOkFdvtQcigUbJ
eeFSihJOyAyqWbFNEGi2kGHogX25MxAGfe/HKPIpJ2fWJQDqCsFTFjAF/c8y7YRydlThYmcEUVid
bZ0KlN+bWQqvIHwvAh2Gioiz9HBW6udLZSjGjdCtPclcSz15Zqu4Fa+wAPAi0bTJllP5o63V2Z0j
k7d9M53gjyMngiqJBOtLLrXtVEaU33u50jcOv0ALis/izDrwsKi2C9fcijE+gUJ8v59lp4cQ1RDs
468q8EVFmOkL2OC8K2WmEW4h8x0s377xnXGsSHc+Ebd8BklGvrnxiSeHjv9R7F0c61CPhaYF6b7K
/XAw7dpi0/yYD9oY/0bSOdMgIRQ3WIDCz5dxJ6q4Kg/fpBD8gBzLMaDuC0S+8Weotp0M6OdnvCxD
hIGWCTnBnWa0qy2cWKRUzs/Dn9QyhF+M3w6TnbppvCHb76BiObmsr04AjIQulTIQutGh+1Cw7C3v
ENaCnUVrExhWqaZKG+PM8k49Mkaa5Kz97Ao91QjC00ANozVVc73dmmVVIWm1s4+Xqe1p+qG6nE9R
z3bmRZUYTe62O8nuTUm2bNMSlFRhhC4qGhyyB7xMs8F0nhxO1/NFjbwV7aGhmJiWfHd2/QqcUJWS
J5NVpxXxUgFM3bIXNhSNMbgkdonQ6j6pOgJ0qL9aBdaus7HfK66iuWDJqArpJmBhnswkV2t2HPK/
h+RZdlf7WJ08kZrG3Yyp+x9b2okWIkgcupc9QO8sRkipiuAxj5cGWQSGtEoInnfk+1bUPYaFLQvM
ztESQWtY115ETIiketwk/nLlPgPzqKEceEVHaYAlJ3Le/MNSGquibMddwwZ7xP05WvcO/fHGw6o1
sswZSRQIq3Lj9y1pOkUVS/7tgv01kQ4MLFNgJeNhUrI7vzzfd2lr5NnHg7GherIaoXNJt75JazJH
IaXciu3siyzw+lgxnrz5JESxBwEWm+ursZ1koIu2/UV7JH7CH0yabew+7DMrtV/wbtVWjENG3pyF
mrg9z/ej3K4y1uldgj45BSIX6TTxRCKpeOTmAsLK9T4/rDoppn6QxLU7KNKP57LAGpptiG6Xn3d8
3MYFMhh42RSHQt4boeKwDzPRopliVLJfgweSgq6+8biRiaoATtViaex3cbQgF9eXSvNe9Il4wU3X
60KW4m1ySiZGOMhUajyvEn3N7nVd69NA7VStebD4F5uVNtjKvPJGW7xZf0OlSZ1ZNzhSJnA4LmHv
amdN3HLHKBqvlYkoCcYV3vcGL5NugfORZtGnm/et0Y9Ybn2JeEgz5BMf4FBmUOoxTgFbOiK0mfuE
WUi7AA4HnqGMvDfiy2t6gM09NBoJOuqhNkMNrv+0DcnuAgtMoI3Mtgcw5ndeOBivCH88nakTDPe8
MbQdA5uDAq8KkKOzvjPISz1nNsm2VA/UyiqE/C7H1O9h1GuRBkuThXkshGrWb4w/dQIRzjktvtm1
EOG7CG/sOid1KuXem7WVqg67xUwvUkptIYelXJpYW4FbvF7ZaXPMwKcYapEMUDrOhMQHe3BoucBo
vqffkEZDcKrnCjz0K5zwnRRbLSIXvTz7F7SD/zP8bu71tsW8n5Li2G37udlUGrj2OtC8rRmIG7ql
EB/WD2sRHe6ySV40RGv/8nAdxiefBRA+LNeWapC1T31oh69/yWTptcM0lnXNOQXdC5En3emmnHXu
jO+738PeB251//imxZQi/3Tkrkp/J+wfAdSCrbXS9BbAVFMZlYMa8YuNc+YtSZZHvT68TaDOCY3q
VhZQsnEBFpzwlpI0Vejkkq8v9XES2glDVWYR97yL+BtRLwjFCLdV2Ikdyx8OrLGZFG2c6NXcN3wC
4mWB+9IUdx4bttArzVoFqYSA+WEhvuz6S/9PbzgCspG8WzO6FNyazW3EQMsRwS7xNfG1ZOvR69+T
TEedpJv+toNRTh5C7VTweV19eXJ2UDgSsuhkcQKwFdW1V12D7UwHOSVa9M7ScFsiH64MHF52DMvt
Y4Qomf6MSI8B0XEGq6FM4z8pQd/eh7wzdjQAg0bmE6BZ4MaDJsWNiiCkivOPxNiuACRr3LHn6XyS
VeD5tjFKS5q/JfsHKxb2Z3nOknpyDTsYmCjArp88GO4VhZiOzR2I6lr7iDEf4DZdeHsvH4iZUIWZ
LJYlINcQT6hryIwykhSbAjpRsmvLm+7vG8e+fOPd1ivn4GcAzrBYItzvpR4a5aL1kaC0a7aO3Pf+
7mFmO/h74UswxULjXQTE8SmXs3kNDG5kRFNFRrAtd3D7opZx+mnqD09XOCT30hs8Vu8DScSU1q+0
tdk0OAj31xQOUzih8NRd8Cc0v/eaoU7VgOsLVn9C9GQYfNc/gsgdE2vEN5FpuzHvYCE3ggqZuvVG
8qIjDo/JjPJ5x9P/O5ujBWQGRZze4U7PLBEUN9IOx8r/RiCXEVmUyu/9YXFvdc1t2hrYTEcxNkYS
A5oVvc5VkIyy6ntbgSMb29ls0e7cdmaImdb8OtwxLTQlxaDQBwr3ZaYKXpoUc9BX2rJ24LYhlwgB
tqKZzUDABDxq9CFRz8KquOXPYs1GXw4ijBG9zS6GjjSNwxJwNAxBPKICNXTGGlfCP7goM8gKauNd
W7ic1ldd8f6p4XT7qTjhJrBTR81S4fchNLqsl27RI6dJ3gkyiA3RA/OzGk9fcLmiAsNEr9dwzc1Y
tkDYTTptNY2yjKIVsA+2MQlYw+clZhgJtXrWvl1oWRaVJKlKdepKkdDk6kBLzKaG+e91YJBpuPVK
lYAqAwh3F2sjbL/Zm6F+spcRwmFKlFT9QmQcvAQ7zm8UZEs+TlcETpHXS9cHIB1AliEgsnftJChe
Dh1bAyD+GmOlH0anW5T8I0NcBHhbf7HdFjZcad9M3+/SAEFNnNM46+3wBzC+e6slfiLfcalMPOLV
taSFI6ueF3vVPWcblXdBUtVUTl+kzJAM7NHy5cHx1Jl/3TGrpVXQOv9levFfxhdvD/Z8TmR4GuxA
fdRl6P8OESINRkkzfJDwT8b6zo1Ftt5DqiQTd+QcuahQAUQV3IyxMy9tKvUm7x4tx4PGKgdCb+PX
oqOPWb8jewzfcpi+lAYWA7F+9z8L/yprGfHTtPwqvPGv0WxLKAJrLlNYhk21OyV9kNDJwlIVAova
OY+NidUNWOya2rgc93SdMuJpePjwYHr2QPFWZDwuBE9WW/XWUeIZTQFpyp9nSGc/qiDA1+uz+f15
h0WL+jggt/BOt87oIYtMICEs/+NC7jWms/Qwf/cxoKiFYLPcny3dnhsulXFV6RpYP+hbT6Qx3Sfi
JMrDFkDtdMp5I3PTJmnUnhcjbWYv5aQeaDRC8ySeKedZGmxcTDVCZoQWFZjTImYVuZps2OZRXhSx
5q/wDWIMdvDusA6NdbRv49EopPB9Z/teFAQOB7TG1EvY6uPTumvrwuDoLowHiNzi6WW/x353MRx4
sxvmywPWZ7emrGr0U1qxRCZFN69dHZQDWvP1+akK/n8j/bVS/5jUQ7Ls5BMvHBx+b1ws842/89iD
wSAhsRlL+UoyYOyBqiFowVLZ5PEyyMe4u6EoBglrRfnrPdNi2Bm+Elviemf/ECzs4LJG13MCzeSq
zbAvdjLz/U66d49BQDCwHseWwHy3GBKNyrHK2AbslagHueAlfjbqnbfhgqgxNjrGyALAKMJsPpsc
8ioH3vZ8q+6yk+oJ2lAfP2bokr6S/W6m51HsCnvaRw2/mJlxNHyDxjVYDTT1nAww63STBkfdqqxc
AyknoninbmWU+dqWi4tdUqzcZPfrEwup754wqMOKgPatyK7Kg0dMNGHJP0zioFSUGRWC4gdfiskC
qrq1e0uf7q6CkvJD2hyjokvvWViq9GOMRnLwu6t6rm1l+j4MirX2GHgECXhRwT+1aKsNd2uVAMuq
Qs3QSbUPVoin9IZnVVVTFUSsfGMtSdDS+h399NbBNcUooTIaZRG9kkqJSOfYQIDDmJixpUX/Ak3s
uskIG9g0RM+IsTzJBemLZJgd7Y5WsB5lkVg3gQu7h6BXTaZGiN2FZhAviwfYZvNC4KSaa9Aq/WW3
7FDoK9sblrB2y+8rPR0wOdkCY9PZPV+Pd1ncfeR9jgxr1XhP288gjnNH3LLbHakQeF0lw+VUpqGa
6559Nup/SLJY40sq6qHhzlDkcXkdAkHMmHbYoWRWmbudS5gixi2LvO8WZjfDixA6pD9W2BvLofuj
cKl0oPkPfLimqKSp0utuNAz1Oyra6HHI1q9zCQoVGtGG2iMthW2m8DcGsm3h9KFm9Qq8vy0ayI3W
ptuaqoS6hM4EXY2mYP747Qu6VW00MwylB2QtZyth3Ka4XZkwONZnAGLGVim4mXRgApAqYjEg8str
BUqo9OX2YaL1IzDGAEsNNg36hXpYkQkWRDI/Le9zf2g6BFIe+ZZTdfcfeq0OA3JG2lm9beMZU9fd
FJc20rMN5foegbuzLnu9wKCXdM6dPhNb04UPCs3mZK0MIDB9PrdiBHxgkDb7aRJM57kzLpouDeYJ
hO4C/f25ZlgnayKcHa2cbuXNg7KOEKkSE8ZrwC1EYo9SzKYMc6IU4s7j4NX0mq0yYGosh+Agfyc7
oqXxjNuDF4k/OI9pSUloolHYrIGjR8cskpxxxnnqnJctEzE20kah3ngeyR44q/5hnZ5jjapuZZVX
AN9PKyPi4HgmgXttgV7AeIN73AnX9IxVs2R0640FRC/vW98Nx3boEIyU1DJNewE+bTuogPBIr3+A
iHlAFtFOmaH1LbLlNDv1u6z2dxvMCDprAzitlTlKzOUnxJMdHnblgDMmyV7yP7CnWoQT0YHtJZON
dP/eaPJFuZSYIRtx6TxZ8KkiCC4sjLe+LOXk02JCiM7wOeBRF7hD2ehpFhKEerx0FXapYCddpS7x
lSgTJAR6n3iXDNx9taVpgRwZzwKUc+T8kuzJfZ+OSWgk93HmZxxkr1xDKxDNWJNrtzZsYBSom81w
NwvLPL8IiakMiIiWzQE0RGnODB8J4Kaw1Dn/iAQHDMUZnFtSahA828YtBGPOybyYllXo2U6Rf+yN
79/+JcYXvr5d0hjZyffNuWmFIB88M5upoT8HC3azVrJQ+jPwdgZX/zzPHX3rZtm6umsVd6EmNMIO
Tn9CgX14R76OvPZ7haJEm5MXudFvefPD8pv2ZD9q79kp7yEoQYtKms+8ATf39I+Kfw4d+Hqfqcuq
ulnzeV7HdlWLQBpGDt/sTuUeNc1DTlT2gjdJM81w/GZb49oWdzL+pedO9lqatVSc+4Mbilgv/rzz
eUtWLXZ+Kek3VcmH8EDqoANlaxKWVWUGHost5HCHdSJJoZhi/zCg4Obo4La7hdJS82qraoesetsS
p/IkKxQZLGLU50qQOu2ddWlIA8fLo1zPDRNDDYY/4QU7H1iCbSIWxKQ7IYrC7Ku4mWuIPEvIQaD7
ZN6R0PuuST3sTOdg90Ma3mxrn1DPz3/XzoWUbJxMqu/YdalbE9LRofZk9sgKLpSdPsfpTL0BhQ6a
BZY5so6R2sIpS5QqmwCszodBoWT22BMxosK5mk8CYX8GeVb+ge1mpq2S4eHPFQU3+JjiRgQDyrJr
Xc0OMUr823TwqfPyr0nclCrk8lgpt5T+6BFfxp5MWUdz5VWUqgJ2KGq+8YirvQtrnTD1u4IE5Lgu
sMsflkdZ8mILqo11cvtWWohJTCGy+zpj1qoMXp+DGKAFUl5+X13Ma/E8STagire9Ayw8HadInUF0
Y2in9/ViV71fjgAHqKpT1HJ8fgp+6D/hmmPUec7ja+EIYoaMHYs0iXcjGMuYZvzUltJz4HbK61dG
iKmaPvqx8loA84nGzicxAuFSjtYDKfogb3dORkwC4l+nAqRnFP5zp70Z2ygdS+0YmXnbaDBy894J
2tBUOJRXpd0ZUiSjaoaAuKFFvvUUP+W4ZoRFi17mTStKXaAEpRBRNJLKwi4TlfTa6TtUzgS+Dw2K
gXjBQUgWRrnQpFOzzY19ElZMWhA7WQd937GV5yC4D+8FoFOsXkne6+4uUmlZn2Sm9I/Lk9Q1Rg0V
bvoZ1vh6eVoL7M6LvQKjvMz+krmOcgxPyTQXfS5StJe30EaRiV83flegt9NjvMSnUe9g5bJ85nPE
OFx3C2jfQJ0hKm4Y/tVcfnZ6U3SgZ5GEyw+bwHhGKbiSeTDQtDXxdsSvBjW0mgjq1Z9D9PYlbVtg
D18nRUULqx6uJWkNWmZi7ZxT9v2S5q9G57GtDzDHVeKryFJiEjUeZGW0i83vqktRAgP3cMOqwkNm
1ZqS4SX89tClZ3h09wxaBwpsGObkj/rRnm9XQO6yF97pHy8C9zlnuow1kW1tQXrPSF+zUY70Bznx
T6yyXCU7qkNDGpX3UazvKIWnmNYHxsb4d8LrGnhwzDNf6VeZzGUtGVLi3+amgbRthf5I1Ny/xGR1
9hhxzl0VbOkEPy8Gnr/v1ilgeopeCcKmnUpsPvYapdomrRfRnaAl4QlTTaPphj/4OzOj1RgwczYF
RE8PdlTbAp5/PjpWRM7C//h0PiM9JUpg7aSoxOxZq/StZxRRWCHe0kEnO/kdvpEnNW3PqYdtWYh4
ik+Fx3THlzOz0I5yYrVODCp6cXyUEat2KiHzeSQSkq/DC+b9Ws8Szfo+CAXZaQjQ7vmAkEscYRnK
6a6xqKF8wDq8TCvP1e1oeL77E9H93E3MI9rXd8p4LTkR7DhOLOTy0va0UWhpwHKwfB1fTORP/6jD
KyGOj52pOCtaxsEjAAUN1+wpGS0JszsWgppOaAFe4fOiaF6LThumw8fGLfHuS5SpZWvjoedk7SAD
hfwYt8plpcHQLQJUFsex6eAMULiQqPWPtrfhGEOfKI8qIeKk79i/qrEKU0ZuysI5EK+Ah3u1z+T7
7hAuVm4V4QZVaxKDYLN2Hh68tR6eoDx3qW5D8aeK792Q24FB/t8v0FXDH6pbgYDaRUzS1H0p+/Ql
Wz9frvKbOfyzACgWI4AWoq90ydGNlIHeLjmHluEHBE2vnBKS0KXs8xS0AJIrmlYvT66s19bGoAq3
0S1Ox7tQxpgP76g3V3HqSUuxiqJRO4DOMmWAPdSB0BKZDO+Hy5AvqqyX1AGdP879HfN+Mb9EHya6
hshhChhyOm84oYY7grRiAj/3At6BBcVcTChqTAtuzCT6953SM8KCt+4kq/trCbXc5xCRFrnJWzYA
o3/JdNEz7y4iU1ZreyU87Pp0+Cd4NYgTOc4pbm+iO438V0wi/Npev1j237rLF4RFuNpUo4jMmTjU
/Y1DxZ3AhK9KK1EVJrEbozZ6DVsr5WqBSgMQ7Ija8an/nig5OSFqm5sdj4hkq018gn+BOIfTUr86
9UpU+yUeQYBAXm+vm67tzP9QkhLrTPwRGb5Ypn2z9QK4e1h+rnT+SqapL6bN4d0i90Erjx/ke761
7a0VE/Jujph7nrFI/IXCccbHjMgHt4nolhI9u/5fyEHElnsq76PfOG6gQAkG+BGY3ZyA/FHBDGIC
/r/KqqUsr1nZ8JLLmrgWAQgMZ9GfcWM+ASJEwIrZexpOpQIlEPRehaHWISOEBPz1hppwx+jzd5+7
W7Th6ZWY1BdA2Hcz3duFZV+wEajAFpSbULfJv7rCLPTJ1Ts/o1tE6AxqHHWhK50MBFi0RgjUGFKO
bbuy69YfKEZXw+eUpHbKrwyaeWPrnnl8B8lCQvKXH2KQ5Sy048EgKl3Szer7ZdIEFM82MCFeK5Q/
ydQ+KlofuE18c4HWoHvaCzxir10kGTNUZrGvogVOzHPZrfAR26vvkmQEd8FHOOu6Mmiuvk6+WR5j
aVTQmU79ASIwpPkerVINDK8C+cR/kTirXHK11GCGPugwPKSFIaSAIttx0U9ui46FHh0DIcWbFJl3
Tpt11jeWDuweKLB90k+OS6GZjPknEJ5hGU8hVz0ixNiS36zfEt3pAEYmmzruYNnWA7L5hSefNUpY
axJMpGl/fR8Q/aJIGloI1gTE4NoL2ZGy0kdVMy8Sb3nWLq+ubpYl3MU0QK5EjuzVzNGGwCQ5lUQi
eP2tnokyDjDcfivKfzH76m38KiFdzTFZ0AekKNy2406KuHBx9ALzU2bBcRDNMHM49Iv6II6Ku1qc
RxnpWw/+xG4ZT8V1E2srbcATSKl8vTatZ7CenG4vFZ4HEpVEYRtWRJlsmWPF7IWa7D2ETZ2SngNJ
PvDwjpRRLOPwC8zlc1phVyK+GKYfvGVmTCNC/IbiNUm4vxbxK8oZX7OMi0VjbHHgYro5a3Ox0vpu
USNNE8BVJ8KcgINGiCr8TVyTe+Zf6PVHTafxwX2IXxCNsfYKia5mAvGADwKTAaJuIvc/JPK9sQKW
TWLK8RiMtQESzkUDsOD4YD0AV+xjpU0I1bl0x0yPBYwIeNtEfNC4eiz/rSbrNAwiLWx8f1hgs2uD
EFVWpvTcYCuTiKUHX8CxFcUszwwtO495iVzI3zHxYpFbUKZvr9DIUZvxt/3nvZQue3DrwnD3yyuO
QRqtpldkwjP9VqsaB38vFYKUrh4uSidli2Uz06wa4kXy96DLkJJBrWEmybr+TlgKj2Ypov1TnqWx
wGu7ml9pW6sdnhcYHvb7QsK90UnCFN2Rn5Q6FQbguI0r/MPieyxd2/HRjTQVF5J3qTyTRMFgCm7r
dqvc0LDiTxO2H+gEoF/EMv9tt7+tY4bVyePZJk3wFpZ/+vbHEY5LeFVXj5XYvwMNSY+8pA8aTwFl
sxqUNcMtDtxHmLnRUHozAcYryJa4iRMuL5RZ4VdYR6BzwHduuyfQd3s/DtIzO1mgbU5kMju/oqUG
+5HUubLV/NVxlbE2NJedYH+ka2Rw+DnuMRYXpG3Omf60Q649QxU1yUYmyXby9LZW53A7KILVoYtY
i9w8Sm8VIihErJAbech3KOJgOWEuDQ4KWQ//jQOV417Lw2bq0KqwqUHowd20naeRewHyCzvyoLNf
hczdTw/sBhH6exlqDsbXjZlsBucD5l0Eycnm0LcZYxfIe9nPGQw2UKxZNUJiJjRalrVB1S47CawR
kUaiiWTDxE0K4AXOg6QzXrahf7y1uero/5Sv4QyuqZSITE0IXgd3gE36MpmO+yHS0dl3JxPOYzv5
H2hwI+SiePB0ly266RLPvoj3xQwMlZp0HPLkqpXuZddf0Mp8a8zDwE9mrSoiJ/vTy2l1SSV0mNFx
Ew4yZmDxWEauzLaBKtmumSbR7go7wp0H5Gc9Mjmd01afE7frOIt1rxhn8ROf8mFfGU9Puz8W7SLw
IhscsE8v98gjni80F/u3hYH5rhOiDxLFxNuiFOLdA6AfvvOw0aKSRUryM68cvYHzuzSrgZMAXTN2
aEw15CekiRTX/PCuIw4OLMjdds9UgWiL35rRHoF5YDpCiyreApDuHCSjUWeorjX2vDTa+757AdCk
CmtkOjQOWTgAXkkynEzAIV/oKWiixyS28r8RaO/IZISM5bCCtMr9dpBoQ1zcR4rdlXhBn07Feo7z
M+s3P6ZjTAco6dFnrrfGu9twI2yp3iLsaQ3LGuyyj4PiAVIH2lR0ct7oYkbHFhAE47MmVnh14C47
I3RMYcYCeCIAAQwpAfgg9pvarAlYRHxv22Gs/Wt1b23+rB1CX6nqqPq4jVHqnMJI6FxHOW5BgINe
TgNTuq7OZP3Dyoov0ALRKyi1o5HjfLh/7bvi2RaFyl5tgETQ63wFkAVxv11NmCikhj4WyTG5VUMr
shDPorOefM2fAh4XOCKfmPiXr7LfIZOroJbC08htEDoe4N4tTfWjgN4/vLpbdiDcXNigbZd5J3WK
DcUK6EBFI/OMpguK9U5sJUBseRf76sD+ivh/LedsfbxnumH2z/1wGQSwpHecbhQY2nAoNwNEf5Oa
VyKt7g0LJnM3PCQm1gAqf0BuXal0ljn6mxpw+RG/fWno9cQ4PsqBiqv76nSEawC02dfwue0XHr0v
44uWnfiWStYC9pN4isY7MWlFnetmhtq+jghvXEKM+CYkVDE7PiagjqpcDfR7g/hdf/4NpvBRzSj0
Swbzd+eS0vcrhWlYUa2MhUHLkJxNdZO8xTGCe/of2zs+ieBiZgTaCWcGH9R6U8JJoNBlbfcw619V
fGqTKMZSjMHOVZm4fMtA7rrVwgA7X70LBly5yaajemWoTloGPeXB0gcuUtEE3uJdOvKhUWgawSNb
PHzMDmwkW/9mNrf4uXs0ZWlMkpEbDNa/mAobyY9ZNjtnI9bqhpl2FHLDrDrRRg5NtDr4MQPRh4KM
fQT3KMHi9ilKtyGkJJF1FxVAMz0/J2Wx5LbbDkTLYOyBchUU/4/jUt55vOmbQJppO+CxXU9s3LEp
Pwk8OLmrFJHsAJUKYKhxkg6KfQlNtaSAzQtk8xiTBCdgmQA/fFYujrMQA/f2t4tMKCfChV6av1r6
R5ZVRHscjx1RL/upfSg00eGrInavYikgOUvXPV/NG6/klVchDBTmwZWtn+Sl5E6etkrC0BuumOdS
ATxUDhf8sLTTrHbgMLHOO19phrUbJi3KPDWQYNbuv1BVl+7XtIRD43XEPwk1WpJNUZfZJXF8VXjp
2Jsh7joVkrR7Er/jMHyL6JzhSEtpBIReTVW833wzp3hpz+vJPm0KE/a4UljuCIESJBpjwVeNhMHQ
yKvcrqvMXxaGqrTmTF0OBaqSZrKeMEt6nz0Knrnf3j32T1C4pXt4rgRBPA4LFkWVwYRIqdPF05oL
utpc2HoO/WtglExi8LXxfDYqv8ct3/X0ib9gX+EzD305vAIG1yrFyHVhZhqzHtUe0LVGaJJXtlrM
69z2RkYQcz/9JQdLDgDVM3CwNIUD07uQfckdoKhdPmxTQaBzY3MSWqyHf6pZkg6wTNF0YcvQ4d3l
8/39drIM//ASc7uGqpfsaJ+wnrIen8kn6tixB3xKfazs9a12Vv+vVGWsDzkHziu6MrmVGyJqWjhj
oL13q7FTt+E+HPeYSvlm/POmRBeXB3vQ1iH8+qlEiut8Ppe8SSTxjqdtxNb4Ikb716GOsXkU5Ydt
U/fzAcjDTnD172BtWDRIws8MPJH0FkFbnsbY8utGpKT3mT50IXpXKo98mIKlMIiHB2F9eeEKzinr
zgsyohws+00JbVvXKC/LCjy+Hdps2G0eeuoaZmCXvXyUYrU1l/l7rudbrBfho74E2vVgVNJ9UDdq
qjLjZxpNNH+VtsJa1GCSrim4d9/1ZvxEb0wZBBRvrLaaN9Yrr5VEpv8gZD/UfLhXy3xSLrrufHW+
umbif8WrY+CPJckCtKOtty6/643SlpVOlu7WYnrdn0vxDV6HXODC7UAeA28Puz+l2XiEx62HwfQe
bIhI7SBlyXfjs2YW/bzw3qxWSvAJNYlWRqJx7csMY18oN8bQwvFc1uEIOWIqvXujy+HlAbSBCoiL
bQTX5q1+aJGSrFEBGLZxWmhlFEvvO1ec4NBNEUhrm/ionl/39b994hirCC3EGlR5ymLtVrbBMdYL
nqI2oEZGu8fDHbX1sJ0KwwVtVokTs2nSApwVNzjFsa0/lCFj+qTxqL5itCSrhifYI+ft+pFHCekC
W7p5ooH7ZZnnoXTa27iud7vTn8i9oohNleHy9M6HLjetiW+b5ZKYmQ6L/v3L8Gjl21r+K/SjU7ry
/ziGfPei78GmqfkBJEJtRGP5KEmsPfv3JtAaU8sIiJRnC+VBr+6GrwyoaCwSa04Ev6tvDPF42tRR
eeUpJav8rrzclFvBvxwMqj3C+es32ZQDXWJnz4nB7yT2o8kExvBF0k74MveUO8WnLtH71cC1Xy5r
WkLcFHPRNb6JKwGQFlC7D3BT6h2DdJ1O5bGl6GspGZE0o0mcHbiI3lf5pdM50bOYdaGfCHi6e/gN
0pYxl9eXxK3R7PjOhSr0uZnGNyWboAgJgteu/PtGdaAYuAqAUK6TyYzZ21mv0+bGYSDm+HI3i7Zs
/Qui5ZCh7h7/MmwqDOxasuKVNm+cze8yqGVBhUIL4ZuvJqWRtdPQ4LSSxEIMc2P55PMVblTkfVKz
J4pBSXZ8DC4tSjHEWbzDVVMN0ql2e//FbEoKS8lHAWe6o7R/ON6HK8ewjCTFnG4C7rJMFn06ZI3V
yjil7XBm/gLDF/UhpDA2ICh/30zk0/iuY8hhOpv/xYC0tCnqFVRD6BIDCAmBQ89+nnJWZCO6pAXF
gRzr9gdvBEAWT2GZbouYMJ8Q2pVe24dr7Qx/zvTPDR0LrhpBl9cvTrV87EgXHIk2B2SbQ8y31sBC
ADcpP+wA8mUoc50tS1Lf5wC+p2u8fvL8+cYHmD0M1UBI0JnorojMNxOkQvAZXzlJS5K9rdMW3aMp
7E8LHOvwzzMu93fVD8J0pyONjoSR1LYOnwOzYiMgW3LHJ77MgWPVTlISAjc/MmzYpEc4R0yJ10TF
Cwz1S1cdT3QvD1RbloaXWdaYcFVu75orlAF2cwyzVnmQqk6jry0WYnHz6zyP0XsAmxiJ2H/vKn2c
CtLZINU2SVeRtwytAtvGrTS4Mwr5xsJH9iSelReEJOLQe5VjRJOZeSPDs6w/udpgzx855788Rell
JdZZXLnPwF87Dp7CtdS3WXe3EWrSF9ENZQ+iJubCPGz0sRba7EtF0/vQBbbHkj00cs3IV2zSqj4e
FciVYLiqYaBKtQ2d4Yqb5mGISsHPwQDwjpR8JBnVdApyTlyaSU8VCsGpBQ/hY71ymSW9AgbtcF6v
nAT/XLgHS0kL8pZ6s2u1zYvOve0pIUJuQYilr65WVr4qIic6a+V0XJA1WtUNWpErZuOVy7NdUfe1
V5rDBEQzovpOgUDDBb86XJWIqRnaqwqRWvMnVzwhGYTxc+ayaWMUbG68VpfElc7YDQdpMII4iZnT
CbpYltZI4eLyl9I+YA3DPoFZ3KL3j2cUaJd5gkiEWzF5ea7eLfv2mYeNvEbXNei2re9DSAGGIdqD
aGvlxUXvOsoZ1RJFGKGzwLjZif5hphjPVwIXcFAztbWDbO24Q/kWef7+Lsu59z5CGF43qXH4MwRT
rfR6MrHUlL/gW2txSrHQnPzxiFilFPSRn25z1pAvpCfgrlOe0DRG02Ibod5OJ0iwMD1h61IZ6pwC
rz2jR2Pu93TVRNN71byYbBDagPdJI5CcK6PKxlwMrWdcMme4sSHCxgkRW2kPAXfiTON2cGcfBTDP
53JSSNXhlohy1Mj5DPW6vPgfy+/Fu87Bwj5yRiUKzZE1+4NTyaXh9pqxnO0zpVS6meZOLRxTL0Rn
zmtBFW91w8LZ5H3FGo8WgaOGueB4rO07GNTlowRGgEZPsTzKfMc69MYFCMSjjTLFiPwQXn3k2en5
HkJgSxY/TmuLcdKkNqORWkvXekQ9hNqGZni50O+yM8xJHHxFK06vIrxMTRWHWZSiBynd0EpYm10S
GTEvOvj8wtFTAQFNhwxVPP72vML02nn/nY6e0zx1lEt2tw0S7FLB9kqpCGBJFmxYkBokk9qajY3q
0Ov+TPV0cp8UWxe307MrKvKfg4yuvPIhFuon25QH1aIfe2HPMKjCgyfuNYj8uOMg9AvhFGRoDsSX
peFZfRxWFOgwLTP8IdpLS43qPt1L6HkY5t/5v/dsku4bWqSQfFJRRmvDRZW8r4SKCNKoNVMvimIi
TxuNhDJbNv6LL65NzjsKEscyItly/ef9c/f7H0DAechMvSoAsZmPRFndSy2BUMwcC7mMbIPDwRro
xS85ITYCr68EnoKNupT7iPva+kXeHl/smjbjS4EQhQInAo1XaC09G11gRf3DxyS4elywzg+mGJXh
k2UFitSy5uOhrfY22Hf5VFyVIDCLts+qS7CPyxiI9+devK8x43qU6k7lPdytm4N0eYZeArk7CJRH
n42jgAuPP6TIslP40NWYbZcDwMozfvNQkyd+2sLK7wd05z8a4v/iqKlwwMtK5e8HwK8rXZz9y9N0
MIzbrc1C2pJUmEG/eMieKoO4h0ForT4iXJ1E69jv86rjNUqjas/5VfRcmbV4kSEPyRpfIeZXQN0Z
qn3S+v2hMTP5Ps0qimHfvEchchu42OLJgz6pMyYmEdoOeeJ7CkvwOT5+miWmC7Z36V17twrt+Ner
rJjgZRJnej3WVdzEwYTRNqM2ShX85+Rn1V4jxTT5g6cModB1PTzjZwjxtTVJjuzhRrtTQCuPz+RW
I0kA//8yEhB2wOE/pk6F8wuUyou9OBngILizCdGcXpmIp67x18BTPrgAfleohU89FkunXk5Rb6gD
+Am4gDWULbIMnQJNOV16BLB7O+/qFu+0zC12eoMDVlR5Avffd6EKSmtHBDhbEk6bk2cmhDSMvdDX
EH0OfBSd1NbHPbvpfCgaKVbVknefFlwQcV1xBnNpCO9FzeHUkiuLo5+NWzLEayfLPo+6qemgGpBF
8rG3jeNB6WFTB/doQANDAVEa07mQUcBllT2xQ+XhAbVPM3WVBvWpNB6ueQQ/tt1/QmyTZIWJpD2i
XE9D6UFcsCJDuMdQ+H8A8E+CxRnKep9mzz3ZRC860ESovzxGy36kf/ar5Y9Q5VVvE2KX3RLPa7OD
iahXskqdCpO+Xvpa2KFA6y6rbeFsG9XbxLbwWYeeHADR61KO+z7kHIXdC/7WMPUhjfEtsg8DjWie
cs7UwVtu1h11cbxoyULz+izOWGZlvUP/FvCjL3Z6MNl5BZOtOJYF3MwywEj+eKZMuHs5t1dYWboA
sQMj9Gw0jdyrNgrOI0s8rj9Iy87NlNc+XyYoBFuUYQyVtIj1gyfKyVf707HWxPCCQqMK6wOIjelD
WC5eDulCnSdZTNDW6t4XrzyXHeSgXaZkpR2asga3ucT1xkjd+jm187BUN2itnVaXYwr2393kjdcM
ZM/U36g4MVS4+e2UTX8hDV9tzGcQKDK7v8irijPDQSbezgO0A+7lje2+Hj+t0JJhlbx9+y6ED3qx
FL3tqHiLoaa3D3bxzn/voVe6sbbkolGFo8Crtkg5AJHdAH2DOstXbdBC3fquMd8TMLzRUvlxLOk6
ZDgF40N5myKhYK984DLYouVymeF0ql5ggnVCgAelTGbPOm+qumQOmfPXNSuai6U1I+XV7GecN//H
WCG0nzDtCQUIu/ezeaM8pmYmmRgPTo5ziOSfVm2PAvoKb8bRgotfScQz8nS4YRet4m4FTVstoxp6
KYXLuXHMhmaU6DSz2LXmtejoE2Q+fKG+eX5reW5gzqeCqIy6ZK30qa38J2JoqFsQ8dIe92yzbXrv
I3gx7wvVpKCnwFIvDY/WmqNtkqU9bRiUBUGdxwjCMHTYUgESE5+LwBBeRHnsm61800MgVtAmAVBi
vX8089DkXLeQHNKKEZxMP6lOCPrlLV3XdLaxlbhks0qqQuKzkwTegldhoiwHDoOwUXcVWgATIioq
24GglEctPprXU7nUUDvNh3j67CvweZcxnRLBM1VSgA+5Z+ASM3k9KcnleMpK5XKoUMYVqs4XQmoe
S5F9Qx9y5vja118BUzu4VXMK7tLecYFCZqEVTVXHZ33HgqW9CKNRn/rDOmTuvA7b6+lQZiJ8eQSF
6WsVn7Kh/z+2K5R1rfe5iBaw2HgqIyvuqXKl6LVcqr6w7IzyvKbJAZNSqOFIDNDYKICGowasZClO
jihVS8XHQR7Qaa+yB9Zcr8FGEqiakV0JZmTy/8Y3ir04fGiHGRKSQBA56SWlnIAiE+gPa/A9n2ag
iTQLys0jeao4MGJX5PA5KNfebKeZ3LP6LOHj2pe/GxMgKOYE/KVrFAOjKdEg26VPaYUi1TGs5M3K
wvqeAcakEuBA6Ydf6Avq/oxmongzMzr24RDnIeDMUCOPct100fAxRf4HS/rYqm0WvFJXk6pLBahR
Ma/oBCMd9Fl36UJsb3izAySfECKQnGAiIbFdoR2M6OELIh9Vj5+uoqgT5b7FwX0Sb9WEJ/4iHCXB
a80RUkouDtO+/EPtoF3aYCGJHomZ2nKprw7y4/6UNbAzyJ5BFNlFEMQPbuYu/j90X4i6fp0r0a1N
iqEjl8JNEcI2JDFhaP6jZk+rFQ9cNruVsw/VJrysZgrmsmbsARAc3YZMBhrPLo6tZsRTpcSevQ83
A+Lrx8fGufTqXuMJ/xn33Eo89NK2pJvgviwGm+Cy5fTF/2tJlxTrBz0UKxTD752RrA/Fj2hfNRqN
DiXxvqyugRmjttDYW/ijMgih+kka1kvj3pS6bzm+QtZ3mk4FBQ8e+i2QachDCiUF3/JI/K3FZmWw
+JyGH+XD04gjzftSDzP2anZ4KS0r4AV3EeiNm1OMjvVoogszi1kMBHBGMBTRGSnMpYByu4dNwaV9
rzjlKd5l561l+nNp+yj28xIvFAxBLIZ3Ju6UU2jVulWc58sUgjDjoJPD7TLUGzHnaa1MZM1et2sa
S0LL0XOQGNiwm/kW6lSLZUSBa2vI2RccJOx3lapLwZZ94N4RwVCGcyaFWf5C9Tu1gHNOlXjQhAhW
DTrklEGuQaijf8yu9WUY9QtJubTWJDUqMFURdXKwI6zIhNw3ibQypCXA+Bq9XxiLc0qIQuzKRVR/
C4kB8G9lSmG1CG9kGHc0+jkNcATECIIoMNWXy7Y/j2J/FoGtT2kMVPXrgKajgcH5hIg7gKVYC0dD
2zDrNnkJLEntKhLZVklTtQJQ3JNEhylYq3P1K9Hvlr4D/8UfF+qJ5TpEEkfhjpGu9R5J3IZNuGEm
G0Yo+m7pEkh/KmrgNAX+c3sm0YgYqau3AhMMHQgQ6QIVSa6KU5kUfNS5rPCBvUZ5H3j5UaFXS+j8
tDL4u4IE53jdZ/Dv230ZE5X2rAr4hUl8QTbPWxbAqiJI4UB7TNFZCJnTzxy/8vb6A/3bDYQWrWpm
I8aDF6efvOw/uLLfuYXzmZlYZD9RBRLjV+hABf3oC83Cf/wYPmj81AZCnc4P7KPt51EN9TmwLc3T
kPebzRFz8fosnn7PBEMBY9nu0biS3AWh3CJaW7qmFpTnz5oB6DR4Fp02tNa4W0X5E/YyK941ycyr
AaSwwhx85XRg85+hFSDxkH/V+ZJMbe14smR0Pk+EC2LbyjCjM7EhyL5ADt/4f5FZUQ4Q78jnIZ7b
xY98W1yxUlqLFlBAx1zQAdVA5YFRRTd6aKDp1WKva3hL0N3fKfnWsccGqA4ktSz+Y6W9H8Jsr1aw
lVD4zBYKJQpsMD0Y9sYT+qwMtluxVAXnW+WH53QgHtbU1k39W1K5QS6w6W4s4m8xdBc8VD7szmEI
hrFPKbO43no2CUqUfm9bgYm6dwqXZSyXRWWlInZPLOo2oS0F/VqBL1PzPuYyw0FMq4naN0OJHgOC
9YxEFb42+Hhew4aOGizk3Sp6I8motjanrm2QYd/d3frM65p0pkSvycAEqe4QxjhIcbbu/Lqru0pK
dWjxs/BZtJwT4KCjP1J/y2KHCw705QpZ62GKUECbKyERNO/cxrm/xvfGpSff2NIGvbkyws/RgDic
mwdIYIt41hcinKLZYC0YI3vwF/GK3DGZDTZlVNKX1BNNMGLcnzvdR1Vctmlr6wsAswx4DkkyFzmZ
Po91jA2bSSew3aPUmQ65FFzBXL32O8lh/e9lF4ztVLkApl/+7q6s7UPbTVHkUjCvQsshzv9Wn15i
6fVHZIBPkrONwNksXT+ltZcgTdZd5fRteEpb/RVOUDNal9pyGJonJJ+/8yGbcLrWD9Fz1uEn1gGh
aTTV8x41e1hINU/20LLD9afmMIMnEwXa7Ugf9c9KYwTVk47NFbVjrS8k3GliNkax822JqAWnWhk4
r3AmDCvj1eo5WVFfFRu4ZiVVw8e2aVO6gt/JU32BD0WMsowlYgq04l00QtVw7hZtvjhAqo5IQTQY
Pywe4TF1F3XA9Fzo8G96Dx7QHSTEPHrL/TRarpQt8SfYf9v7CIx1MqDouYIOos7Yhv1Ou3qh8eTU
7P5lCcfCdAI+Arw2YXFYrGSkZfRFtee1pnPTjM62ykHprJClXdvEElY21Ua4E+e/temzYTimeboh
vz2D1ZwSr3BSVZsXWFEKARbHjG9PSXn94HTzkcV55XXJcXw6jHKeMZLDErXUYb/iYplv/nmIGOx8
Z7ddqR7nFbls+0vxmvGjoBN/hgGhGKAxetvUABy/+660LSe1XwDo9NCVodaIOKHLBQY4YD13lKOm
Yf65ZtCtBSImX8vSJ7YQUaMQCGJte1/J8UuUSvTpFeoVd0aznh8+TZCqvGfvWW0Rr5kJTJwB36wv
Z03AzygM6FrkB1ugAirxQguqWw14tGzecqofsZJUR0yHKtk+inbm9ZcIMOUuwJ0UcDz8YFNG3Q64
H8M4Fc8BoiWul97193Z3QC3IVZw8rMrZ6FjKLimrkqvJ2+rf/xNkA+w7rg1kvMQGBlQwLW8yRcFf
B8NGLyRGxT+T18OmumnndmpgzynUxlcPbCmdvqH9aJveGyUkcioS+3qW+zVETeKq4Rkkm0jHfC0J
LCKY2gdoXtPBSDMb2ZHYlhuQEr5brWbfXU7EdnCXel0pWgpg89qeIf+vGkQN3rNoRyMAiFwLpnaC
L5k3r371mwfpvqCAPCFkZig2ebowp2hDsEoPx0L3xel8CgGpauh9RCo3lS9eugIlgaLHlSKW86xF
fIVQ/kkrINRd5zmwrLrXBrKmXqollv1i4BYktp7kFWoELRUmDjIIcoQkyQQsoAPdDLHpAKJedSQQ
lgYnHGh1MEl+/PFGfYUttvhbxR1BfnNvRDwGO+fRL/yaejoGMVLbc2ZkYRpYbxe0Mv8yqQfM6UcJ
4/OH0+RyMmymHo2aENKc90mLm3DhbCdNwwz5RqVRiWjUTJHshZox9S6PEXVxxjWfT+ZQoLn9BqTu
2VCsrYwx9p6eMttDG/n5E7hML/T2azOx3BNWbWXj4mHJNbjqpFtEz3Zaq+O20OLLEApOwtw5nOYB
benyzlKTGeQHcPY6btXOS78tUwa691u3o9DAH8/oVuQXUDodgwy1CoHIPmn+B3Kq5rhWm4AYGBmB
7AZlcQXYAKUzYbPX5oqAfA0LKo/nUpi5/weol9BQ4UQqpIPYnkU/QjtHlniz+yvjiNKm644422N5
x4UmTnd9QJ/gvkSCKGEPMfSzhbpaiXjXyA/ZMjovfk7XMpmP4eis0iK5l8OVO2lHbjzD6AuX57PA
UXFsYc5y3JBMRAS2xX3VAo8XhUWTKnQJOipINpY0R2b2qc8zpgLFH2Y/L7FE74/80+9DIWbqc79J
Kb5P8HfjES1LFEgExRTcgNLYA5338Ffh9j2GeWQBZxkgmvOcFPV0wGFyITwssvKfYNcaSOPCUS+r
Y6XPssHqA8BgsBYYAAzjjwaL+Tm9OBh4x2VANhhZHacPW/1h1AVfniK2vVetUzSxzwmnud1fwmlf
+hIUa0JLN3KJfhFjtGrneSBXosjz+Pzc/7e6GTCNJ/emEFL1yhk7gfGYA/W8YvTTx6u8fedjN3ke
HBpI55IVqDhMbjquWjIB/Gp7F1CBmx4vwWNqOSii+f8Zcd9CovuOzvmJcOX0RIoytmgQ3lS8RnHM
kd8e5W9ZeUxQ/8sw8IFRtHSCOCiCHvtV7kZAPh/CC2p13DfBSHO7OpRQAr1LS+fEY5cuovkHQxXc
XJfxPW5reRFRi8mwHdTbHcCEe75Z9Nq3TEnbihXtAqMtjTNpZjOmaB4ly7PJPUqYF7vZTmyKxopO
LzJjIKT08CJ2MsUbIsqJ5PkbBdkYeU1IFJHTtnUdV5tHQAVc+zEYXmIFSI+FrhQA9EhZY/q2XIBA
Kvqa6DM4omMi/S+AJqgvgafnwIiRj+M7GLYPLSQo81MyHxww3/oWHbe/uiOH6vY6Xa6gNsmGKHR1
BpcG+3ail4MagJotedxsE1tEvwLFbRkA4/HW5szA50RlbZ9lQi66VZe7gA0aiZxNQQ9fbLLuxioI
RvAbG2i/T7ELqcbLqbW6X+g0yzop+utBUYtA0sP44JOaMTierJm5y5wqK5g0GQpxTrSy9UWhZ2Ud
xk8X0ZJdqXuzV6QfRf4tWg+oOhvGnf0uWERDWVvv5xuWBCikf8iEo2tMPirTWlzc6DJPvFyW9MB8
AGcUFmMaEjMW8CHpfN8RNzDwScVCIknX4uBKwCQrJLGe9DqWsaNuYiQBWjEzt3VnUyZNKJPj8Vld
ypD4j1swd+RDVxY9Oqy6j3RwGzLgYBQXVskfZpdai+2kfGkZrOWoH/TuSSSpXF9UIUCHl+2iKn5S
uuDSyiE95hJnBT7AZEzRMNF4aOC0fRcJhYo/eYi2Bz8PuKvx9/FnzxQPL98y9i/hhyPCM9nUW0YB
oSZVzFimWyxRyCJQDb7vuTPrpL173XaKCFdZ+yfpLm3GmFH35N0wwrsrbH6v8q9g+glDihUPci31
yMqlYE4MCDUOCPgPsIrU4dP4JLN7iEMvd0oWWyHHiuVa3GA0Hpq6fKMJmLymTSxW4HbIw+8Gg1qw
MWNu69eXYk1G/+QcEpAWAx2i2qbeQWUSbrpZGoXdYhVz86xPYHsCwjPeTiDfNAf2h/283i6wypzf
NdQz5AE677B/58J6oZ9g0YMkLV9FJ2gGzv/IVYOzua7MLk/GdkdGaCXWm4bdKrdu4YrAiVxBY/lA
3OSJu2/tQve6zWGfsiL3Y82QIQIcQvseD32H2pedkxMmRkm8TNo+eP4iXsTFuThnZK3c5OUIAXgj
fjBvY07VHm0gEwwuymOg+WXW0lLA4EbKEfh/OMcYmRnuDQJ3fXjBQli4E4Iway7rzJrF0CymEvv8
ug6aXQnNF7ezZsoisdH45RelmaG17uA2dlW/3RV7NeTwyTCEXdMMLXKNa4E20sdqYyw9hp5+2FSX
rjBDw8eK/H7w7n8naY8cyg91AhHoGqXpcpsUwA2Lfycm8CTEGmTI4GJ0pzoVMCkT+552vjT6r7jM
eycVYFdrSb7qTdaC6c8CgBj6kdS03x7h6nbNZfuB8flc8sGRA4h3Pz99kaKd1+4grbGqK0zigLhY
SbZq8SW71GjI+hXfHi/yC05ro0QsUr10vZxU1MRQAKb73+ePumxOido2F+K7DgHPUM4XwDsYmOez
agcnSf8neoiByQ5Eu8m7bAzOwWXKjrPhxYZo5eDZvC7Jtd2BDAEE3P7/YLPdaJ/5bsw3E9TPmFo+
oJK2/dpaun4Ab/RCvYGJbnIwxLLkOTlTxCk8G0+4eCfnjOawjd+sRVhFZHwdRjvPzDsNa3iaj93A
1vB+owzm64AxAQstbdVFR5PHLUVeKNjQ9BkNqoypUXuHBxAOJsCmEQRBRM4EYos55GMPDyw0qwvz
bbAnUGR2w8+glT7jmjR1V+mwQl0tklSROzrGGvWvmVsikZ9HylJ/6nApEkDD58fqiwZJL0hTmT17
nosWuqhIBCOGIh2m95GZmNhnJeMPb7F8KiroeK4VMg/K3deTJgmW0hIK+jDs8UzYuTQP6U4aN9h+
dZTTgRdgDExKeuN7JlZDkHRaCXsVqnehJUnG+q5iBB02hbCtiqhEUrfnBEz4pPmk7p9Dc89XRzMW
Dm0lNn9mM1mpsRoZ6eWyFL5HzDf+b/VKwUbMqdkl7Jgmek0HF8MAEV75UC3kYSO+F5M4A1HrxGAw
Frfa8rMolHxeuiA6frk8RJnzk4k7wuTERlSJJM3cTbHFDFxqH7dtW04Y5bJOn1dIz2v8LqHdxRU4
vzIExvE4I+46iTH9FcEAdEI8zbLQovxJ1eJ8QyYy/5jPjr63RSTGPJPii/qsvhoZV6AaNEF/gWuI
mGUVPWsp6h65SuNLFdcXeOhkdeS88ZQ1kmthXMmXNyqLEhLfVgs1n9eSEb5L7i6L8DV6KrIFmisB
ReJdydtHkeqxLIQkjA/zLrGH9duKgMB7OMtEnXLe7eOsP3VEkEV6wC5IrJEV9ayUoQ+P3TqFmx1H
B3gVB3aVr409fP6mArdGTnSEuxKUgwpUDZZ3FST+RkDbWcbN+O404Is5fNd+sdgo9GUIIveDzliU
fAigXO+lOYYcm7XI9G2ZzNJsR9KrRPhhXvG+wYf2XK6vdkzG7oP1DxwAXbUx8unYV2Mjjw9Cl+zt
x44GW1JS35YtdxI420E6RJF1zlb8tJDvR9Zp+135wNCd3pWXGppEDqEc/8mYoOIvyEa34+tLbO81
I0Fx7iQVXSKsxkskThwbzJ1eE51rz5dlYsxgfBVnT3Xhhu5R4XBvKBrK0CU738Pxiu1IaPhzLknX
MrU76JFB1NnQx28v8Wiqnzhz3mUClPACs26G26Ydg9QPBGQYq6yfdpwMwUhl+Vk6JEHLOKoXCere
x/3/0GUsOG/Jbc3mdDuQ00xYoKnQiHXSsDlTT/AB9ljluVwUfxQvPXmxa90Iygdu7ghxtqnnlYzC
V026m0WAefsCywyZQChnP2CaQkJMAsho1ct1qkSPmR6hzZ2YlyGJkVfK334P2uCaAjTUffkxf5QC
M3EpoN//Tj/g4UVzevMozgUt/HHKjaEmfBsRoSHNcDxA9gzoBOM2M2Wd7bvJD9Km+i7MfoSPY+mg
/9ooEJIc0fdylYKEkK2ZLYmnvDP+M4kTGIwLlGct3NcoGl1If4eRewvcylQPzRTJYrqxGIbjBkZA
bPtIHw5fAe6f+CWusMbqlEH1VFfyZ0FQ70A2CIUJKTvXKhn+bY7rorL1ghNhEBux6XL6uRgLoaJa
mcpx0aZdW6z+ByfeeDUG2+iPp//pjDhSOslC2dyoJMC2BPrjFwQwg48bU/xzNW5REAqmYFYdv4e2
7hwYxxQJKZeIcF3/P+p/m+qW2tUvQohD2X8aDQTDTX2TPCOblCZgUsfg3fK7FPGiFWiZUy5sxgFj
rtT2vbVmLlrBEvVJqRcHZD1cErWR/AFZaUR2ecTqXoChzNH8XldbpKQYbBjJB78LFddTKxS/875Z
aqjgyvs+0LBjn+KwrOpw78OxCuA1VS1N/sloN2C8OUKECXGj8CsX+LawqrtKqrq5g7OOEU8PZJld
KmD2M1NoNhWXDCS+QXwWUZ/JQ2SCfj43rDuQQmjQWV45TPjYcCV0XCjciI4gXLq0WHsym8z2IaXL
jABuivLHwwQFvkfK9gUTALTTcXj4QpDyrRF0ZnQcEqrhwfrqwyVLyoWfVNdA6hEyoWCPbYhRfGK/
9m3sBO19DYs0ge4hqtfinL4odY7ZUK/zrkSJhq6v59u7Xu9yuFBPmCWegny91XE/+eg0viOda9my
zNaiNzOOJ1SHGnOVjSzEiamEPldj+s73LIrH2TI2H9DeHmGRs/Qd+a8X3bnc8nLoWJZ+vlj5qWC1
+zT7VLJoAOOxT6AX1+EefCkgEM4xJfgDDt/MebcqoOrVQL8BfhcUnZJxGxdSXz+QP40sVN3/kyrf
SiMqtyBXwaMF2Av4DurkbP44SAfDtbuF8acjW9fG2j5MHkSH0/fBXGBWjMJBfqnnXtAD+CTaJhe6
SYNRPE0V3BAnCu6mF7qEnu1sQvl/493UarmBD8+iQtR+KmEQb1BfeMSMTHPJwR63eZWkMuMpr1vd
j3TNstvm+fqMZi0IVii3sEVQq8rrgQonnNE+U2eHho5Vno/mq5mycMXOTAMmLiSzU9xdU+ARW7Ac
CBjZKiDjbQaxqqsoxCkrI3/HA55PYAzLkMJQOjlzdWwm2wpZEli10e3W3vqLovxFai4GsEMxktY/
4NGm6RD1MWVzuUJUD+5DEhhnHM1slTspYo0Pd4QTe/9OXLk/iyAe18L59h2AiEO+aB5LYSvy8c/H
8XPbVKoXzFHvDTFp6InddAmt246bNd2LWlfK3XBlfpovkJw2KwVDGCPKSGiNxMYCwpAC6/q7ncp7
jLct+BtOFx7cRmZ3e6u2zt5w5ZaNCUAHEahO6NUdagweCnb65X59cYBglUv49Bd2+RTNTuKQKNIt
dSlXOVewuqy58d/ww3FFNuMi+/RkhEINO183Xa3oQCX4Ci3I/z5DV8ZyTchR09yL/9zO1V54rQ8i
1hCaHnTj8LYcDHRubo69RyfB1MzWxYGFvILG+09PvgDK5AN9mo97Ky6PV3ZlF83WWz2KAFk0FkvY
HKBU+PlDH29ZcjcRdL+GUp015RwysVpU8nx5VJTky7pW9JOnPEQrK5wtT0Q7W+yoLr4Dq3rcX5h+
5w+DCdnKLIsu2AA+T0yz7Vv+z5zetaEVlTRu7x03QGb3oEDbj4ChfRf/+Ycc7vkG5tZBYhRLqkAg
6Y41vWb6EME3Rh/CEu96UVomvyldgJweExGytWBD1JSpbUIp8DfNIunrrcrdvxZu90o3+8bMSiHl
nfDzAi64BvWVyx3QAWJkFaaLzw+HDt8EVDhoFb++rjQJ5yEudHClykJL/EyY3ocSjHw7Lds0eIkt
G0FlOmVPIqx/qPne/3Kf34f46asSBJT7c5CKldsHTQOWKYytwBjnR5GF0PpxNjFHW5lKhn81QLLz
fEWZ4b2H92fn+VdsA0UAGvuaJlPVfI74ePbArO9EIuvGAKD0184zhyzm5jKEuPHQpu8Q+8TpsyKi
kG3buPv/OrtSSrNE4wTuisJXJkAh3+aFKUnFQBu7RAgZtov1wmnvcIcBg7HKB9AurPf65oMhUgGz
8VppQdpV/QLq0x+TgCRNQh0nlvjMq/DbuBo3dsdlH/E1CF3aD4oJLE9v1BN1u0DkoN+3DbNIxTgV
q4AumE1smLQZ+SPBSYP4hsD0vKF7+1AJbgG1b+ZPCH9Y0ccrtV7sMJ7uENjg2iqSzpCZd5P5E20n
tewPREmSTCD6Mldz25Z3bzjYMaLZpXAVm94x6Z3x/hs+6Xn+WYfzkFRbVgBfgfZorGmRHnrYWyGZ
kPdNiL7IGsHD4E+iTrCH2hdvSd9Rh79eiu98ftBqnVNjOnBAaO/NeR95iQQiV8HsJ0vp8FAhZMK5
/pmvdn28lSCMELnWIQ09Ctlu1cEei9BHs2qGp6hD3H5dOgC3XHilMboGCYDheAQ2vKMcoS1siTSG
DAW1a9rqdAEb4AN9ZoVFkrOYrE2Rfb3IEb/JRaM7kBk3bfuL6KxxkX44ucqzuG0XMYUI0STuEo+D
aQH0RGPBJeWE9UY5siRBlsIZv+wbMx7XNV7ioG+T6zrrhCZOez8P+Im4EI78iedm39mifcgnZl/R
kFFdibyyHTbrvjappkmYx4jiaQ/NfKh2QEaCsSY/g4mPoe5SchE2IMDjTFVbjX7b+31yaYdiymeR
zBJSebMJ+YyOANgjrmKVyTA1wSmJSqNh2zfZopmZlW53ScHzXRsQ2bIk3vV/MpUnCkuE4/mMDD56
cNNroX7dRKQogJeZOQUxPUFg8RUSqdAMG29Ps6ZFAFLQ/lepxC1iCwwLO/v/ZYOu98Fh4McdYvb+
zmMrvcKAufdxlNCkbl1Acd+woOesWYukaiRtikCJI+BtrgegnEHm0SrUY8YUejGBnl6vjRGoJrlN
KnTW1EF0ZQQMsCfIvxta9IPvlHjkFw38zTuOkd3Yh+KyfCYWOLktQyj+1Q80nUUYXch6R775CY+H
/jJmU94grM0uP2g+stS1ekBFQU7wDqqWyU4TAyTWLW+gyO3K+YuMfEL9YCAyVETHDvxn7Yrx3QVi
N/v6CAbX8MPSm7GRLA7NGD8yprUq+6za5v0qqz00H06FmFQdLCdr3z3tAGSvAbiHI+gjzruu4KWD
O27XTJI/BcvFfUzT97xZ78Uog8VL7THA3Er123+9169GqXdAxA9E1d/+y/GSSDnWBpsJ1PJR6dTc
pvtx60WYtMXI4hG1D2jOVD5kngaKCGIUsV+ajG/EUQXUHc6z2uNSqRzCJ3JszcEbrruwsxYHeOjA
yPYH2WQYZktCLPi3JPYBKquw4QLaTN0yzEiRAoXFJPrN4BulBwSZAw4tNLNfAdOMTA1iSgF9Ln8n
Qpu70dyvD5ROjGlpDOFyrQ5mXPFBSYD1HzQJQUU6bXrnRlG5g1xkC9GcRrFlMpJpg6cKlifkhdnZ
Fy6eLw2HEw2sOCKuY8neYJ2bhyL3uiR80BDSany2kqiqb6Mvr56vwiZ14PmvSvm2zVP2oGhvBMQH
nEzkeQ2/iUZjahBi8V620T+FK/qd+B5IXVqiaWSAdhISsZimt2xwWGtNezsFrQMwdGH2MtZVuT4T
KrxI23QNvZkHS3c+1HjpkB3Vm0k0V2x1LJSD+E+givbXL0lQ95Bk0HlU0AzGABKrVJFISUwok1+Q
+Q3x9l/BQ7YZ6avsRo/CiDkDS2E54DHHl8uFzEIg+x3vAqriPEP3eB0icB+I+cwWQPcyj3mr8Phj
xAs2yP7VYniM+5VUC02Rdk9LAVfjxlWrAwaynda2anppiorSMQ9YhaWXBvFWfDX2ardCqJlc/lK9
i+xeN0Tyf7xmggDpXCS1EvRYgIKPLpaRfY4staxI8yKf7VL1KZR4MU1pZRW7VI/d+vuDe4oc5HNo
3dNHmsantzs6ERzrMUKqX0ym9dc7dAEsmbxBJ4nGhY46S8xPTl5xUUZfpjTqLKwfMpSFbmzZ4lT+
3DfzDzO9MCfAzjtIQg63VDzz+k/ihLx1wCKHetrG3YZG+bVa4YHJlmIrDSYWMqWglmzEDZXgAyWT
k2dbvuXse0i14SIYWKd4TR9kWIOZniWgKvUrIt2XPUiCVWW9s3IFHgydPX3ZtvmhZBv3yASi8M7M
F2ulTmLs0VjjT1qUroGompeBLHLzwICoTByKbdGhhwmb0y/bErSUkkame6pwUwQZLoEj0d1Okinc
/L52ovY9clI9NrFY6e4vSBNAALVUW16BYX3uo/pWJ3fGGnenf6ZOa6RxYZrXt6t/J1Pxkl+KRgsv
z5kKl7ucN/YIz5Bdo4sst3JF/m3/5pEZH41nTTW1jru4ORVSdfEA06asWEYn0gZ67eH3/6lVnU52
9Jj25BeryK6pKxNvbyciRQXJLcb9Sj9fL9xKtLKggkJTdlDeVw9zswBaWnJd0SoKIb1DQbrjPwYc
uKeu5YMpQw6vn9ikPFvPdAMTQ0H9K+aBDhXYxIqQmwNYdZo739qFzqzXb15ioIyYrbovYRCg0wEe
jEJWa/NqGAMXkyK59N6h8HF1H7KlDzvd6wjvWRddOdkbgMMAIsTGz7XpdnEVPSYL1cMrly9bAGuG
j8XHp13yCAZnq8up0SZTSn+03kiH/wrhXc7mFQG9xnKzME88yb5eDbxYw5pa6FSmMtaHMEGJ8Akb
8GrXRD7rzjRDgyvDdn1mUsT45WWfGUM5nrJEr/mmwrxDDlRqaFiSK3wtefr/K8Z6cjLiohD5ytk+
Et1IRa0vGtBlFg8Kem20AU46EzG1xJC/eAb1YvuxAy/mN+RoHxWeer0/pHoEQKOf5w2n5nnMkmsR
3F7dyWibD3/WyzLRzD88ZgKFBXg1oE/2O2hjPKNcf0/Qov5pKOE/tDvNdjuhgYqW/DwIqtfcdN/O
wiVgZ/TWnukpdcsfwWK8ahyvQxlSrQrH0rHMCP2lsf498r1iD+V81Hupcss2Do+8jTMWWwtftiYe
6drJV+mPrTjopJxtaJ7sV+xdIOqC6JIKD5vtAfffwAUim1z9yeVBCK5hG9LN55wYIdvEoQSmTe6y
XL1gTcsKE1Wtt8T3lfwlXksKmdowSWHQoOimjNqvpZphqtensgZvFe8DbuwKBEGMkvffiUr6shzM
APo3nlNe+QXu8FjNupyq7/4kJJ2KdPhYrKhkOTaQfIMCNHf/bTpcGRsxkKc7tlG/tF8J/gRARObG
nK2tlauoccqrzGNmebiaBvUEC7AnY70SyekQT6j7Q3IWoI9++anV01i5tnYRqAhgk1KFialZG3TE
1cl5lObbB5R2TizIpWeqv9GDtzJusbNnNBW2zIIqAq/b16Qe58gLZ1OgUuakHRRm+khjIujRJywM
P4XlTGpA2IoB6M5nH30fBOD8EauSUK99OQ0nJSa6PQBkkPUwhgu3NHLTANBxlq3ArQrwwaERISce
9NZ/bXiUVOzVEfljlv6MDuY/V/8liJ0F1zpEamHy3d4YsLVuJO7P2flWCrljnj+ix29T0u+5gTP6
kiUMIBH83L0CRJ23AzckBAbOE48vrytFJpHZHHbz0Xjau/caeZbnNfbXEOazxLu+E+WV4OUzglfJ
/HPJSfqTyOk5HwtmUhnu8s8jrwgNaoxJdr0U7DaCrzEUhtQ2ru+d99iPX+qt6VrkgQkSwubq2+u5
K0rquADvu+dqGp+AjsMpflb0Kkiszta2PiPSzf0UmLV8uwGC8Ua0y0pWNMI3W3lo4t12grIl1yhk
leJpbUq+Wt1Pcvir6MwC86Ll/27IUl6IJ7Llde6ff10bAwTsMYCY7w1xpzKZxNcbiF4aCHmqwJm6
jvI7FQbxaqMZaRVEPxgTijWzAiu+74Dv1zYpa2kp9opeUfnaKG0Ay/pjSXSNzJ+VL9McUYPLRSZF
qCxtqVlE0e8NW2N+ma1DG4jfDpmLbNWbQCloZYB4euaD2t/54wHvuC4qHTrIBK9Faeo4QUKrzB5G
efdQdD9eWbZbLRup5teBpsJC7H9YOn411qcp8Nd8FEfS6YsQ2cGmIn+4cR2WEsmdnfvsD9c7eABk
4HFXMrU4WAfFWbthhMA4qTHBOx259WotOIqNPg0w0S307REILEMKyaoHQ6QnAhd6RsVR+Ip96fD8
9C2vTekZuuZmY74OxaWJ69kdGqlKikH3LGNxTn+JQcFHLdfwJXHU2tKV+x4hPAmDI4mlgTYhFaxm
Px7acIpTqNopY1kzRJCdpHSGL6e05r/kxw8y61XM5EBYWiCPoSWjA9tUbtDp2Z2OTQVbMOsvjz4W
BLO+Fs1q43m6HthMw5fGrgilGa1KiQWvju69i8TTb0DOd7+VP3qeEfckHzaK9OPfP2qwydKx7PMB
C+t6xd6S1cHEa8+TpkXyGjZPdFhM7Qxd2nwWe/pisvMRAaNA8CPQhX33HAqiGdlIfLGYsg5USV89
yxrqrwHgpAAzXqCqa4uuwVaMFbviuqIRoS92NNuxSimMq+vJHYqC8b3H7CgV6igPvFKb3n9h52Bv
+g49xzr2traf7jrlnSmthfJLdk8wgiQarPqS2+kdbgb4LQGzvMgiWbOYB0PA99YLF+lYs6f645Re
pIAb2C2OvidD79QmvM2eMHHgYXkvRdv7eOh5EQtwM9N/S7J6Z6kCjQkA7fRO7ZaxlG8vJ4LvKtgq
vm6gUYGGTVhhdJ8BPtDyVTrfHthpaSP/qAEtfTlzGUARuzqsZ6IIAy1wvpusz41F78FP7njas9ZB
xgEdpzyxYyLrZkVQyDvezEYawILvQ6ge1bkAetegtGV5xEY+2iP3nugIaCSQ0SOnKSfYleXj+twq
jR34eMC9D9qXg2rzsPYpZmtgUMZfgPQcnJDGNpTsyGRtlBXWStL3Y++JZYesdB7HswSkMbEfEGE4
lba7MfJ9gsypP8aJz4lr3s+mqt+H86AFc2+37E50Y1nB9f1oVbqX+pCplfMU+hvcYK/Y1rgfFIHr
psfsF0wwbSrQs1mbJAZIHBKbVjq85T3yOaK8r4K8/QP/keebziFZsSWvaGPcqFYLOYF8KxgJ2N8g
mz3A2GMod9RRS5NrBH+wYWnbFXmPWkLxCrU/5iRu2zp/4ehE6Vbg3KQ25VyIHQebwk0Y0s5EnNbS
57x30ztOb7YWorfrUwWAs9EpIimNkeS50jyifiFgW8679mjrob3Lebbmw64kvvCYSX/A+kqzBXIE
YaXFYJcapcNqlF64T5umL3GZqpqvpcI44aYzQWhFCYAGgjGjfQtW0uj+qZrgdAafkUlkQxE8zCzj
LCIMcUJv1vXp5xrzNsK8Ta2ySczMZU55yTWQrGamZDGKVeMxUt/BkAVfuweHG+9Jg51Bh5lUG/xU
cULbLxWep9/iwI1NgVMzJb7g+n9cdts/KqeRvAN9la7pPTZ0IlYeG5ll6jhmN0kPIjxglPIjtmnr
yjejng852xzfsz8Y40Lp3nD2AdE4OIp0F4CrDJ2TeWBZiSx3qX/8Ueo4um4lTM/cCMKhzRL049kV
YKhkdiMLAqQ/y8I5ItISYgpl7pWGIuqfUc1uZypCJPF8cOBJLzku+2/1vKCDKL9k3tWc/EeRVXBz
Bm/0xoalAxWqqNjS1fAFiYDE1ucWvY07ptNCyP9Zz8wAozmH2A2lzpPw+WjdXMabiMnUBCR1rllR
1uGyq1NdeqZMY0kLSmdPuZbBjfgGSMAh5G7Ofyfw/qhXtgPsmaK7c/TOxzJbHAqlIfhf9l83mU4U
I200XrvgKG0pcP3B3FXZd884prMK/Z7hUyvxKU4mAGxKjBN4LkFrfXvPmRmS0cBIWCzTeffZWFvC
YAyuOYpu7DHGi0nqqFe5SAQLxV8dnH5Y9lKx5M5/mqzBbLVxCyNzbP8CNIxd4xyMsXSxZOC/cp1b
yx42vVPRwLeJBW4lsi0wvxhFjJ9UdmVzafipJebnqqOzuMLPRAVvDGr7ikGbIICDIrQhr7YVoM3p
FYWlI9xWDTuk5/0kYfadfs+bLcon/s9EJ+LwQYcI6zgP+NDB096u3ONoTw/axhIgYDYIXg1Er0Vz
obu8v9A8hcMZx2W/JHl7dmN2pVcR2JkTkOgkTvOfEg8XBC5VQiUwC/S86uuUH/CeZICHo5NZY6zt
/BQWcfVLvE1irEWcwk4jJi24zKdlgQ8Sa6P53GHzP+o+8SzVG2o4vAMw2MC9GETQgw1jd0fZArVY
Q8/A5AJtWEx+igYqJK9qCiwyg4ioDbUN8rmkwGSzrwneMWXzG+jCKkwRj8zoIgwCyAdz/MGiQE1q
CklaMlBy0GsY5qWfPaMiZYs11TW5uJufuCRJwiP3sA/NOKTpcW3UI3RwKe1Y+pYp/9ILkoQkNSrS
/O6yTOOOAp8fLSVPbM4AmT+NzJ9Ip8Q63DxAnAAkQhX5uPIBAXkDazbbk5plfP+1E1uTgwadrq9C
cDoKr9jT2sU08Pe1olmJtX9wemDqkxcVCAPIfKzCOTF2L37lDRMQzcnYKVHwUYjR9w0epUGMl5sS
IVjVEMKOPoEfTCydBOmpSOqGabnycRB3/H2itrtXYq4kbjbp+hh/9y+/6eN0UUWi0DBH2Uo1r6ip
5R1IHETquttB8rRfo9Lje1bqaYWYRKy+YGhf12ItqC+dJTVjIatK28LAkic5T3EI3JAn5k2awcja
szOH95AqNUeK1OI0dr/XWxlk47a6jeERBC4fYg5zJQ/OohFvgkgfwzxdDltSe3lMJc/P8NWERE7z
Gm+m1AVA+1yD599ZsUt0SGyEV/U8f+Z7KUAKsthREp/NZOd8oywZL3wik2ZWiFiBX2Wy5xflED34
5HbFfxwdybMCVBe2prze7vqXLDKv1rFRm6ikW0Q7eU3UgLaRUp1a1V13EclRL3rGIBJEMpJjzX4e
aVtIAtsCHOcz4yc0hwJ96EYZ7yOEDy4Ga4GYYuQFxfz/BpSnZt6AOGyzCupvssripqS5sm9v7qHN
WvNZkYj0zxEDptQFIVEkhP/G98R8Q5u8RRhjJoHVgKkoGnykQ8e/iqA5O8lo/PE/G+m/UoIpixbX
kEGOT3DS+Wm73746BQBUEzkD/wr1GlXN2SZmZaSttJ4HvKBJ5FfZVrmeRzBOtU2j49NHFM8uGykt
nDu8SzDVT1xDx7KxKfSG7ubUjNjMsFqBnp/GmPc8jyF3t6vLPw3ucJVBp+hxC6CAq+lmvVtaHEhi
yBjeIYOG4x/h2pQdr1NBcgqS5JUuYzYblv3rOJRjlSixx19zv6A1sy7MoJwry9tRe4RSxjxDD35M
6v+3Qwxxm8DYCsiGuG9/Em0OGBeifZJyP4KTZGrzGRX6QiNHe8vrdCeeNZBNVwJgj4UFSckBN8nQ
9ZeSYs/1jHJg9aOF6jTAxjBu7VFpKlUZYp5hYgMv38771FjZH4G/CWIhTJIHrzPoTCf21ooBw/7X
WJBZloqvXu+aPFHgUs4jwmcg65CP47qOJlrGKG50x1JUSmmqmwK/3w3DyaKcxA2Z+Dd0gyv7YGWv
+l2QFMwu3QOA5SRw5hE0myq+MUSgG79zAUTwAAbQM1ghkAIDDS2lz5Lu5Zwbvnsqrjh4jih4Sg1q
3ceZKg0YRas24UEKD9q2KXE86I4QihsQiiXw2sSrzRvB4R5sHo+wZzwKbt+aGO9caC20G9DZ+uCu
bQGvDBnrxIlHamhMKF7IZgmDZ8fYIbp93UemChgVip3TIw3/uRvm4aTea+LQhkRrc5l2GpoBMTcR
jbQitILVQXK2rks83yPgebBqFciooxiBLrKG+ggpYU4hw7+zVkPBvinMQlsL/MoWHLFsp8Au4p2S
YcmN43A8m/5be1is7Ybs04uQ6KVX1kzCEkVqmlUmV+aVp3mzbG7P8eTL96QOhnNIpYPSUKn18FPK
jwO3WjLPsfvcWCm3mmZCJzY/qKHj4CLzYmKZbhWy8OoqkPGB25xI3nAwTh7q/nNpADzCazsLXTie
bGCQnuNLYcGtQk5QyhqEvTk3vB4YTUD4uLYw+Lo432tFypq7oYu/8cTFRrJ30zwN2M0yvv2QD6TN
Dr9SlYC7FuXysiJPyRmI7zZvCb0phbwFb0WeMUiJTfGMCwe1oxbXjndZrylFygfEqxT3GctBR7f/
TLbK9vDbpcXr24UrntNREQPGgYoENI4Xk/ldRnoTz5HmRbu7b/a50IBLABEMQtFEwyoUjI47dIhS
2OvOT2JD4PB83+4a6cef1wfDBx1dKuRPFXLq2Br6JE81LTRla52rG/WiRSC7hGSv+TS9E9o6raPB
CVGvLv3SpV9PX44255Rrl29q9Y9eoWjAGn7fuBxiqJ6T7vCQF82Qn78lQsUGuXwTwtiHY/XJSMlD
RcKz0I5ZnmSJJFu/8swiRCpuEcCZMPS/LCDxRtNOeMtz0+dVTIFfH/3d7evZ+mhFoLQETNQQMFDu
tmx3iBXU6Jd6XQiZ8C4tY+rJHhtr878urhtt91s3yA6j5y9P//kfSM+TcBbcqO00W8IK5iiuiegS
ly+V1ueM1fBhm1BweOvsjtZOyHI1b/fDVCD6B/oWr/lRQ0IYOQ6EXqj9D6hXXMAsU5dafUrI1RuZ
nR6GvzQIoK8zzBL2mrIU0Whbd0vJgEtQgf51LxbuejdbTV/bH6EEy5F/yOJvxW3ihthhHL9MlEyc
Soc3OnIIyQX01w+nTxEvhNI9RsQywBTG7eOIkGlLep0mkc7oDHWfoz9WkJkTnreChWKC17V9KXEp
jwJ8pCogTWG9QLke6hAmKf4lENqVc6iVzEBnCmveyNdb3yZCE3D7si9fuOtv9S/iFpAbN99Nem8Q
jUUQA1aI9knJweSTqPZiST4nzHNFUITl8DhVbi8YSn8swwvmSil6tEJT5uCGhrQgiOSSein/TAEd
Dmu67WXMrgL5bqH/MEqiVy2ij5Uo96io6nc8xL4Z2kaBcV1P4kvw6It8EwOh5pYSBTpyxGiWxqn7
N3HDmWSZ11wNt9lN+ItKHgcmBA9PItd3tsnGKzrklYkrGQK73qMbUiWNstxVfq1CQDPgf1fFL5j1
TOtAXnk7phATEVdxYu4uB9yecFSB6OI1bFPJNsNLCeZcmaseheuT4SMK3mxHGYSI/+zVTUtk0ycg
68uV8WqM9R/Kb1MNTizjttWnxgogaBoWKfSyzosqh6qjGDVn+bl2CJrhpo8uupHdOd6c3GReY5rQ
VN0M8A7N4T7Y5H5LuCNb+8WNaif/rpvDxoWU2AonplDrVeSc6NVJBlnKyRnyf52Q7/1yfCsAIb7s
NQw2vBCTetkx2tQtq4aCmLSeaN5N0s9/ez+GnZoGGVDCnE378Q4kWCRx2HcZLUi44DMxXsocKpaa
XxdcW113pFGYU3ptG4iow8ABh11wAKRdAYUJEdNNlTwyA6JX3NjpM0IiNAVUJqmhjf/RO9XCJ0nv
yAXx7v7BDT9owGbYHcSU59FFPuPBmfe6tMoC0RU2R7tSiG8Q8TtOhs9O9iYUd4YgYXXhElr+ge5D
mOsDp0Kr9CeXSsqEKIj8iGYP2OvjV4UdeuwvdkxFIYdeqUzm0/fX71IKwjfdP4hVpSfI3ovdDGiW
KhYG5FEoDcfJdQjQY4e1xxCMpRfmwpVq6qUy2DijOfpmNhoProexadlCvCxknU7TjvZVKWcuakzE
hwe9cDIFCi+4fhH+kUHcMn4dlfVFpEdt3LtUpw9IVBHnFIVoHj8IOZ9MLRReE4YXTrNSKcpJPeK/
KLd5CY3IsBNmGgwz/wgaXlRRq519ekJXTTbemU5d6GkMhCtcr5EG5+acZ23QDYiOeFcl8ntzFSvc
Tymv9lWaiihNLCw5b81RpulRMQzrLICDhZhHTDou2EmSMnsliI64wRLm2JQgTix+5mDzw//Fqc81
ErKd/bVj7W/xvU5gf3j0C8NC9kjZqijlV70KxDRHd8f8Pcvip1/Mwi32KTUaoIRk2XG3zEzcoAi1
PqpvjnPh+KCtsP3xhzQ99TA2Mu6qpFgHu2vx8afI+o0gQCcrTs9rgmaTaht5TcbaPFIB8E/JxGBS
z0aQePJNz5+S+h+T8M04N3b5FDEmcYoscCHQI+hNPWLLP1qVlZpzhJB34cf2gjGPSjys6WcpKO9F
e3prQyidr/J8ewrlh+ZswiXkucv0cY9NzHDVqdiKCmAPXplo1O8Pz4ztFxz2WCn/dWjkG7waMdbt
9rNL3M6niexUttAN3zaB4G3bzhT/JbHSS6Hhn8SJ3EEfGxenr3Wgr2VtFK/iATFpZnv0ZjkpaLpR
CxMnspg4p5fUbUwotbfwiS096KHhqwCjbf8DoY03a1xh+YZcFRuzkZ1nBuXORHJc3WtvobpgIgGY
BdbRHAg/T+KvO26AOz66nZum0ioB5AdEg+ROCA7S4dIwGixVyo9eCGrBXJgTrD8UipSixgTFYFOp
jWSAvYIogcTczizBNRhcJeCMZgCdXvE3QnJl81vgYyIb/jjp6cuLBWhy3WwyPRKkyrzBJbDcFbyX
d0BuBIMahp0qmT8goJxymNsD4DYmaVHaqRntjS4tmOve6U4x69UxpGaws2ffUinnEFPpZG0Eu5hz
4Z7SsGJ9H1UFHl8pSFOJIYGa5nIE4y0D1lhk1Vz9F4caNFU3dXLGBoqT93iaP3ywi8lA2fjQRqgh
yBvvx0moONylm/UOqRaQ9QRmkE1VS2sHBROO6by/spSDt3+6kk6rjPI03vFoIFb97ij0gYfBRVsU
Li8Wbkeq2V6zmr3ym/pGGgKn6kHUwlYXgTteK2JMPXvvkPR8H+YIcuTlMw0IKfLR0kO1Zrebq5j3
bYnFUL2OxBxjqfxvaqJ4BFKb+iBKPQ+c36MPylv5+i7xPbM3mLgozURr4y9f9rzp1iJxi5E10cqM
F3v6sXmdsfGy4ZNmgCYXV+c9dGknZDaiSMpiF/aPsqDs2GwXT5LknL8nw6+E+sLiK1jla0IZVp4p
WyFGUAGQA5HKPIWy9H9tY6ZuCkVbDP9bOXGrix3+ZrGda+MJUxQmt73+N2t8P/WgUNE3Eqb6mNk/
LXxrMUjwzRg4T6lRcJ+lcW2qLptuInLGafieVFSa4Qt0Ypr7VoS9hqtzqNKbRVJn8z4L5hNm8ccg
s/TVCv04VqyK02XKDeYVQDzskmemB+vPs8dp7rlzZPlER00m7/qZwIZHvlBAIRwd+lrXwZ46Gq+W
Hli7gQ6IizzJIGebT/ulL7M43i/tBBrfuQd687Lh14ZIfYf2rETJ1Y7kVyYcMZyk34P2xufZDg/H
sEo7Ck1zogW9ttDvuHpYFwtxqlLO9TCZsvAlepfaXZEjudHueiZxkFeQYcy1o+d4OyLsLBDLL/1H
5NjjDzXWgxNzcKXxZU/n+J6f5A6KWJu1NANJ3oe0Ai9jA7Wi+vqXhzh560FJhnwAbRSkL/uRePqN
9RH67NRlqthSY2GPweRY+wduvb9xAd/XDkf2o9RsSNIRKlTTUjv9cjsejvd1te5yLzbBkmPPuvr+
hE6tMbUkAF5VkBf0I/5BUrlpN4JQL+J94ycvjCyEc3hqReehBq4lVZ3V0fUTyD2/hWvKmx5eN552
p9Wq/4L30m6Lmrr/t8zyaAoTuUcASiQlvXRZQfoLzG4ncLOIhjQnrhqgZ+FWm6KMVB3jM5cCMGDz
A8jdyXkLwGNeM4iZlFMyybd90Ib2nrL3ILnYRhRJ4t+KxezjWmdBjt8DM0MWy/TcktDl9efvtOFb
kaRzkDBQiBYPVWKec4YAjPzSV2+C2frJD/PhO4OshDzDx02EzXTX41EFz33Y7bPY6hjTdBgPaIOW
d5hwkgD1LZP/sCl4f5rRWnexUyeFl6nux0uX1pwx/L60vWDBKODsRpZIkSHW4SbEYJpCGlzF4lg7
bcIH5nuWpwm5L0Ul8a+H5z6dSJWotwdNfCzOopZ4fRWgb4RbcJWfWdiPhXa2OWjdnVR20ap2B3zu
2RqLXpxJ31YnpBFt4meKPVp5zy3OpjHPvuY8VySu/e6dcwdZZTP13jsUnVLVeSPJExwe0lmAI7Wl
BFBgzjeWgNT1DhT1lph9Cr9+8a63HGCXd48bLdPcEtbtMuLrLCUmqN3sp312YHzaZNNS6xFJpuha
w+6Tsa22q8nEepYHf61GmRP517uCpgBFnoKzSROhLQ/2DHskCyMs0qDoztIHV5W9aJukysBpQa7q
O8sQ2KuMlJZtgLVGYI9cWKZoox/jWiAU0ViRkLh2ev0y30wv9u1RtclS1VB9JlFgX6JMnNg//JX2
wN04/EKHpBlAjskW06RDarBspYx8D8hmY2t7oLqwdwxmYcoMnE0QvOczkhmSZvRd2wnNaD3mAhKy
kKHxHLn2K/bx1R6bXVVCY2nZyx5g1Hvu0waSdU9AQMgqNv0/sF/nkCAOG1mmfHG9EB35SL9PLUE1
TIk0IljFB/PzSyBR+MSY9ZXWKv5IwPChAafhk+I51KdOMtgpngIWB+uRIP3Y5M6UDSR37mvNuDV5
MVC8cr2IK79ls9+/9U/W+MjDqB3R4eLi23rt3yShpeV078Nf+6jMndME74CSyCkpfJOIwiL3HLVv
9WAwRG5vP1E556pufjWCQSTmjeWfd4GUlrYDj7J+jHJDyABsKT9ASUFr+o0HKEnPEAe5q68XO9u/
eNpd7LAb0aqKJTIMKhf6T0kyTlATrZ0KGI3gVfpREdX0gNlNztiYioe3aOTIbDf/WVKaUx7zWAi7
0X/uy2LGi52X+rsJ9wIBYIQSwA4Ut52lEpfDobvi/In4FGXKw7Dmya8g2GDhGd0LvSn1dVRoNk2g
38bZHiMiM9/ORlDkK0kfUH3aaRFddEAR8Kk5SQKz+TXOZC3VTiizQkOm3by+eBw4o7cx7yuadmtg
MwMnXvyg1gzDIdteLM6Pr/uxMsmK5kxNstxQbic9JooNPeCDuJxwtmzPugb/DrZSQq4uqIyR38fx
Kn7JtRH3BlYiKVidnmnp6+/4cWLSKTBdQc7vJhBuT6zV7KYJ806lQDoqUTZ2MDWMjmjNaFzm808Q
8nD+l4hcOOe6q3vBveDGDzo8F4AHSLL+VFlCaI9Mf+eiAQyAg3d0fus7NkMg2c5hmPI+kv12VIEA
AQRqBabEpmywpR1BXXfjEG7GUBhjgeJrpqCdTtUNOZpqZAX9SpR+hbb8p8oMeoQfEuhY4IlGoOtE
BzAn7OVv5uHYP89QrBc0oji3p8XgcOpYg/JWShHXZSjNZ5p2eMY8EbgKKWxq1pdr+bMJPI8BU7ff
iLFZiyexrulHORASomuQvlZsqXEgIFPmVa4zu9mn6il+ki4t1P6PgcKg0/kXEFfBed2DPUuVBGqe
dMeKKYbpqNLt0EthNUDBFueVXSXA4hri+OKdhqKAwmfGS+qLYm72g2F+8pqBkj3CWXpMO4TiTQzA
jrkFDqHZiKWHoyEvz0tkMW0ZpNf8vvcyIUcayvH933oOAQkz3Mf5RTwmXVnuaa8uK4mOYTSko4CS
2BnPq58C1Zu4CEgmGvLtzqIVI9Ik2w73qglNorOnIKORuBlxu/ENYxkCthXHMB2KaetkgAThLZ68
8susvdir0yHLXAUE/qQKoSs0X90YzW0o09FMXZvb/GrSPpNdzLqhBITP0iPjpmz0i3RSUfYhGKoD
WzD0aCZnODSN5FhNl9FP0vdWQW8r8QXgRzSlmJMPWkYk+jB2cwC3a/bHdvDcW8ETXmbJouoCfmm7
4UZUyNxpaJxNTL8m3aw2T3y3bLeq/kUTd/1y3WN9XPAiJMHXoYqtB9AlcO5Gr4eePCs9eaPDNGHS
MFDTUFGPiufuc7eAWzZGvKq/rUZPfSQL16sItAwSkwlhdIJcieUO86pR/S2HQWbuR1R68Vxld0Uc
cy4dQRj/UKWrlLyqMUp89fXmE6O0uWg/GOidkNFcnaheka3Jpv8E9YeMxzDb6NCHmdOB0IeAOmDw
Da89lHYrmwR6B9gCENmBs8ovO76SxVjXPXtbzsXTP5utcl6NlsG9k130ZvLyIhidmASr61gopeHC
gbwGlV2pKO4gDTKTQhH8N8NrTHJdJNr1fSXvFqqwJdd1XaxiqBzvrh76N363s1b0Cb2XR3Tsx4Q5
Dz303dIrCZ4rG1lHT56bx56dU+cYmrKhYmsRlLkeTNtc2HltOxqHFBx9rFVRZrtzg1dwGk3J4tyh
Q0Bxg1a1s00t9LEg5ruwbYWFTxI5WKbkQq8Dj3byLc26JFL344St9n8BCRrNnAohSBfDRjKrLCub
q1trkVT2zBlPq1P26loSmM0xl5TSaG7wSh3TuDQpBLajV5bvXUFohtwkkedbJgDxlOJlrO9d3qnT
cq1hvfqyTZmxoCmJgWQnjhhHM01FlmpA+/EqIB9YGJcYR0QtYtiI5EBwGMUgpf2fdO5x/gVUxSnl
kNjCRlF6bJPC7/5PWyQQz50Itf5iJRIx56cf5ECPdO0pGvNCLC3GcXR6Pfa3Y1N+UMa1mrH4ltzS
5LLpfeTqrm2LJr+/BuTOpiboMF8GhtUcyEiMx5puMRIXbQeAVoPG/2CQL1Nq+T20BwR3Va1YbpHs
gVORLPbBLeZINybcpvkwBy25MxkOSy/nFuJ5zDeSqWTGuEt7eK0X9ypEbDuwCFJGby53ruxpvAFL
9eynaLkw5rPjgB+xn/yGkCBKOFD2SlpvutVVknfC9qrqQLKBwrPglB4C3gUe4cQtjCaUMVTlBhOt
V0aa8nYfQbDpReRVQ/Q+BNoPNMYQPfZFmhsKZaqdKN3YQBRGWBOIpWp55ErGnyzcEyz/HHLUuKDC
JlwBJBdQS3K8TXtrze0Yfya6iHNm8vCQPhmNbei0QLt5NeDSEkthmYHLa5bJMTGiOFC7qwIQKISy
UURVDF6waFKazXZam0buO5miu9FyhJI3cNqzL7QQZEFMzwJuaQHcoZn8Bn4g8GsmW/6LqfE3tpPM
ASxQ1Y5b5qPPneAgDZgPpO7j7a+pHRvUfAEGaqCWSexYeaMmS1RxXe+ubq9b7qWicgPyLvW4HkyG
eonbMNdbaSTh9aNYttl7szvobbz1sP95MOVTu80Hw+weHUWsSnBJYq7YGKGFknOX/eloaPhtVO2G
x8h/SFJXOTLpb3go7a+T5p6efSCGTg03UltCCWRVf9ZoqzbXuJNFx1XckSC680/nE6AaRp2lF3zT
ZVUad/37+gZQ9iUJdb/34ZSi3UWb+HS1T11AoDshBQTk+L+jYdX1V4Qhl1qyczYb6rhb5qF6S+UG
QVIVOT4un4uH2X7cNGX1ArDRfSoSNhLSJgitZ72Bz8OKd9txsWPS/QgMap4aSMBo2DBWSZ94C5TG
0djDXyP2x0CfcqoJ1T4ztQUkCUGHqqlzbJn2clPJKR6n7XlZG1qzZtRpSAKuJAZB/KfRUPKPcPUL
fk2RZ+5qHXY1/k07/56T1njhfL3vEv9NeEG9PaOpD7pE+/yN6Jd6vs7fSRTu9KhOYpcKxN42Ucri
Jb34rp2QGP1QDjzdUFA0Glf3Mx8zsfz15EI+V4w2S2lzIsvnIqyMp6vKGtNgOKbFxuUhgMSAM65B
eQgggbLBggLJ+40J+5Gggp+jNAqAxhL5CcBKYUt6rehq2kq7i2k6Jb7zbtliesxo594WlFiIaRnq
Ab/Ci8jW8lyDfEysThCvgZO616nxrgg=
`protect end_protected

