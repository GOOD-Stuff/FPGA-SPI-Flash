

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
NtyLCYL5/3rfRWX3XIUWoCyJypNOH9cIu+d+Hqwx6gD9tTUVuLJoOBkvN/BbGHIv+gHzbebnGJ07
gT9c2od1Nw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
gOvt00Uo43u2bKjWtQoTcla6e9cy8DigekFHOAFvmHLARM0er2069D0sJrV+Re+Z0pNJyi6G8RrG
7xF3eUwAm2HM7vum+Ypx+PLpFTVtAE3qcos/KdoFVruQ+2KR4xm6ct5GHE7I4I7kHpb47V1n3A7m
KsVZ9Q4Gj78XZiTnAcI=


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ezxkbRJZF8baEvYrEgt01fk39VlF4Vy9oPkF/Tcr/ZSXWZrN3Ny/64ZRk5rdp3/Rw4mQWdsVpddN
NR61Y/lHKqyzIFy5av4Fc1hvtJ5QrGu7jT0itvr42t0ZsKBOir24UhbMtyEqR3CR5fLeSQGsmFTF
dv3KWzF70ty9bmZVSQA=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
qGx0a/xTrbWGkdXtnErSWmLH57NqWqgsuujHfQ7lkXQ/8JEV7zaMMf6MlTKUSECLGX+Hvc0If1o2
8pSBoaczpNUPnVU68eGXWinC4mD31mx47odaV1wlH8fsVQbGMdBKqBWy9TuX5hg0WgT32g0BqluF
Ofaj+TwzvjOXbyxmTJFJC6smWfhzgJpDMFRCbwUgDfK0WLgNt0hs7vmOlNiRXaaxSMTGYh92RFiS
NxDABUW6vw4h+bGTVG3JhrkJ5qwKlmYlO4SD/jiqQmKrtaue8mcj0lTSTYM6SCCabd0uW94N/8tu
lzw529SU01QAq4RGqkkbg/FyEhRVNeYtMYy67g==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
g0cGT4TvnX48hcFZPn8fyr0BfDW/3mBT+7tkdfyWZShlmQV898cMKehzh5fGzmgpbgvX00nKxBTj
WeqyMahjKMWih08yRdHR3vNUJnu+cL6RFX9ce+T45X4jsmlXx/3XSRkdmnxonh8czuQZQRxMS6Qf
ofXembsqKBHB1Mfw0IzbD7aczjkxwFftGUuZ5OCU3B2FYe98Uxzn8zJLzvzLLD6qQ2ZHMoZA/Twb
InQ/RCbLhXp3ETIjJwF0wkbmIOXTthHHlTDEzXaE4esRBAX05vSi+2cCAm8ofWSaUHrEc0c87M3K
dgyF62TnK+GOK+n/yPM+tHzqnQJ/S1y5eCwMhg==


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
XJM5nAzNvkSjBrtMy6mR1RzFhNDHeLRKo6RsiRuAYypLrtq9GNYqKE+wyYP+Vo7xVBHdMLdP/8W+
MnvqKQLx4Vam4wQ7/3p6kO6JOKSLHgO7ujNfnfqKtGP5+wiWMQ3ayWgmNFExkMDOh15tsG7/M+BC
kP250ud6s5Rg3PFm7qO0LeVdlNevnOWFcNZmchQ4swQ72GBoyxzYh71u7WHuvzvMmFL6nu5Ag6sT
g2+Tuyl0MjRDJ2cHrBEG9/s/oPnSR3A8+jIaMFQDUdNMGg/gKLbDe0nvtFEwcxj3UItyerS1gTi1
knhxeuAu+zuveWwBMOLo3qGmEy9ucUl/jCOSWQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 214512)
`protect data_block
4QbAj4C899pCydbwSo3MApfZlt+OVDAX5womdmM5R9edtN8JrW6aHg6hviO7xS22cRUPnfYeeLxf
ymD3Usr6TCsYtRw//dvnxfYHnC8QjVGcmtBlDUD/B9sSMIIRc/o9xPOA4xgeW21riptMefWAEDcK
jtWq2QRzsHXSi7n85m+Fc+qNC/D8NY3X56HzHFYzUiVHpYAfwfNb6oZBi2GL7J7yhcs4pQ5i7YZH
PQ1I2Yz2x5XlEvsivfpD7jiSBF6CJl0rkhbpcc8PnGMshq1nFU3oKvFgmnknjoRBll5UsTv7VljK
7sCEzhTUYDkAiXSWFapX/VZUzGSQDaBluApKBmSrlILQ1SzgNJK82Syi9Uq9/s9efRSxBA4lwE7l
Ig0YSOtcNTwJvbpWXyCcO4pxzEdwSCHoODnPcVmyh/e9Emn385VmZjMmaaKlHJL6JCL/9wclnZZm
7kgGTOW08s5h/uXobZgplwJ8VN6U+OdS5sk+/+YXZQ87W5xufaFrlkZqawqArI7BDVf/mw2cvLmX
kUdKPih7X5/y5G+a/ka8gSl4ctUxeMZyM/DCXzestufh3zjQlkXIOSdlkGayv1Q15Q6VKrlQ3GsO
k41ivNtUeeqmSS40Y31m4mVBKJ9fUyIx0GvaYQgvX9+BsJv0uxh8sQf+7irIp6lmJAIkotFj3UQl
JLrFZ4Ciwv4u7E8P6vhlrAQD7jSadT4GiDBWDWdqsKmRQX7tndk8cJGU8txjPZoPNDcEWNBEhzNl
w9ewLLRUVWOvyziN51KQ08TIviVOsp/DWQAVgrK/qbb7hgsgxgCShej84zszGaDPf8598L+F0AFB
PukPCREMpuVcprD1Ez2JisanWPbV7X2VbOkJXNSdyXEiEp8jSDm0AdXgk94YfGFge8m2PDR2irNl
/dvfJSDQ1YFdEApnDdnZPlg5mpyEQZsTpzT4AEKsUJzgaBTCtAubRdirWzrgtG4jsNxG5NJEFnJE
OSyEzimTp8Oyjp7dAxN+pln6+Oww9Q4+1lQ8lugKvp31vxzIxPP1b5hSSgBdMREDEmbW9QeyW7za
gVI8S3jNsAJDvyNMXuBT3oNGWMUHTywi9brHxMAhV1Bq6XSA5Qe/ADzD352NQqnAVENt5noppzgM
NYqiD1o5W3GrZ99EXoNO7idq0uzdyDDgJx7XpSV9gVKRxmP999Znhslu+wb+ebu343V0s5R6sV8g
hoF7GTqx8LbNAOyumo/yZyTxy4z377V1clkFzLExQP3aakbmWYhDDltVXQ0aV1N90fqopyaStOSx
JKvoVFvAXu8bZ8meZozUoX9TLuAe6+shxeOCRpqo3cLVWasgtCc4/EK48wlRbqzNrvtudG9DwU0M
JZEzfNe1Aj+qw6zDrt0Qqq3+D6aTut2gVyHDsA38wa8naANrX61KUOTDX3vcv8sXrhKsC7Slhjn5
nMsuZpXwDmR5OT0/E8zC67TqlPeAljQArPET2ML+pjbc0ECkzSdB+utFsjIvkVu3RJTfnk5a4YV9
IJEV8d/4zpn/sMvS2Jvuojt10j15LWGOnNLJF+bSMUV6EAmL8DoZmMDVi+baP0rL8jDD4+k35jQZ
ks150zBcrO59ClgdekpGOYAJQ6ue8Db5KyCZ1FxUWIxc/fC7HSHb7Sfw3Yl3YbIDZIh5FRCpn3si
z+Qf4yTTbRKDTcxxYFfcpw9pEmcueKqruZFz889/9D4S+KpkzDuug9SshB6yr5GPG6nXDMP5ffiQ
LB2Zxgx/uK5hvcFVi5p4LTxJwOFgr+wA8Zo0nj7XWLFTpQ/DjVf6YUcGceXZF3VMfIYZkrKlHl04
7O2Le2cCon7MzFaywiYovL75Aip4XP8LnXOqqNBEn2WiQpFjWZh8uwhoOWSW0FZTdrkcDln8IpUs
B1svJm8n5OmMR3K1vdYhUZk+nJulWa63sJua/+lFPbAGiqmzS5lEe0/Hfy+ADp31rMFlr2pgW3Wa
AxmPBgSAUxKSzhmBqU0oK1TrS4unOMlPiH9ZOjDT1YEaUl7l0eDgnbgwaQFQ9X/xKqv7rGBB/NMW
VBRvyWIAchmOXd5+6YhzI7cAnq4Rxa4Tq7SCW2thw6Z/+AKvAQ4yqtz9qub+2KKIYVMjpee85nZJ
V4YYFCz5/oRIeQdXPXKw05LhCzabyBVxOG/BdUoRDD5X6efGE/H/TycDQ+T4BGJO0DxHwi+Kx2/q
9oeZqXlRnYY9r3QMxr0JchwYGNP37pb6MlIt9VE73IoMaiffXhAcLqhjS4S18pLb2WVRFMWmh/DR
28rxUeiJgjOko1W/4kGnCpp6Hl9SVT2UTMWdYUm7fgy+SqV+VbF57dxqvyWADXjs2/ngi3C8R2a4
dS3XsVQKGiaqD1odvZ2MlHbpwP4SQM+vEdVH+HRFcjc1sGXkMc+BnqxltxBHTSe9Os4HKfAYBP7W
X0ngjP5r167XCajFKfcW07p+bydKCaomjr6VDmn45LsgIPdOAqRMoOGrbiljHpKzdyJku8cS8fD9
EH2Um666LOJ16REd1ag4hAHUXh8sohYGClCy8WhQ8/rBTSwV7vvieZjuT39YaSnh0MOZbiXkijPy
1FbH95TmsuMqZ6kGXmjBZ2E3Yo7uLrisQiIRUXj3XI6EL7+zaT3vhpML85bLJbGcBeuJVfZdN+SG
yx961gOVrzuQkJg69TWf6Amgy/ALH0h6K4l6qOneXq449Au8CporjBhjvZ320aQhfdge96jN8jo7
J/dcwUUiQfsFe4kkpbxjpcCqrcEOjwGp8ivLgliURDLYs/E8unqidzS//A+valYy5yklm1r7OsQo
SbthRSYSVNRktQs118Cv/E5r89aR0wS1VN+QJBKWOAW6KNKoo18iClYQ4XGbLYSX/AxR9HWUNI7s
1SpTlfxX/doO0yWkCT339pqiLt0TfukUiRG0ogaTrVz9PTZghnueT03mH2zOHa82E22/5nTcvvBn
ng23WVhYFmpt4KdZBAoyEv5rU/OMdSzKcP280v/mOEtbA0FitXQUCIWpJsdRz32ieoFNlYauQawl
myQRC3Ii2c++H9u+Dv4CbhT6EhijSMtY4Ez9qIQwXDc4Ky3SpUmTzDju5db+iPPFaJuPZ14JUWu8
aTeNOCa642FETd+OU3eQHpzRqoZ9Aqlqwe4FPx0ss4hmR1sIih4kzomILpQ506t4ffuDXyezgpnE
czH/cX4FVtpmNTUNlc3Kcniq2aspRCASHi3oCPeN+zkxS445kSyoci7jXwP1N5h5bTRFgpLSeLFw
rX32YPYKquuh5/Y6THBEJrJl07ILOHfmTQbiMGIYs8CTq8zR9Jkvxd/z8Lzu1B1/OVsQ1kJN1DqZ
do3Acab+nVG620PXCaCrfdHxE7AIHdakx/IKkHWHBTUmwFhNgfuSH2EDk7O93DjFRq9fWw/02XAU
tpAQSVv7BA3ZwuA8AVrB0ystkggQNsk9sCHcxV0uC76LIMwF2bsJPOCHcU6CjWbASz37g3xjNR0z
eOgcj++RZBxrwxzrj7rJELuug4dQ5MpNjN47AHB7KXisWq8YSFiKHy6/Ep4/kuNwO6BJhlTkWCZl
y3PC3bftd0mIlE38EinYk9HiZT8krsBRYTd2qk82kjrA4DKV/1KRhRGU5iT2fAQ2gtUKqnh7tLFR
WinAvveK5zstAekBqo3J1mLLTVpmfYBbc5002pAxC8zT2YTzyVN3t0Np/bNb7cANLDq4fdKsScOJ
GnWv+JaA5+HMuxqEVzEjiicKtitdDe4LxZUSCWTSeRnzb/Vyyjy1bDzl0g/qhG4i/si/kETpsg2l
9zGVG62nc0GVHQmEVD7FCxSKnpfbtHg+4IhY5tGqqGIPAzYMKfgYu3HSk5TFANeENb72ArdnZZRo
F9u16frugntj6L8gfu+rbMIju6FGiDqOwY9oZkW0+DjGobuDNcuHjctm8Ht0QaMOJw9NFMyMMUQi
H0IHtsWVy9DwpB227tceEe/RLnlWaS4F4KZ4eUE9WWpUwXlI3xM7KR1Eat0Yjm3j7LC6g+BadGGx
jCtfhudKpya3tD4W2oxO4LAgony02HS1ibbm959pStWqhvhpAQExkEhN9dHcSrL9GhQ1CkKtTnyv
OB0kPKFtlDZ/+4qGlxb+j3yGoRaqKej+Iw6+SRcVWZCPmNtm8O+qx9VIR92/WdZKCDB5lgZ89mFl
pAl0AsZ+G4/BvXqTNhB3x67e4xio8utTzkwjrX0zn9P05imB1VL0Zu5lWTqCFeIqRH5/6jmCuLbh
gA799XQ0Z4kXRVVhLTF0FD2qJbDLTzGvL0p2K8ObMhKRkbS60DFLjTmTnK00BE/R4Z7xr43b6frs
OOMi7niaDBU7dNLrNuOq7Vptm9wWk1k9Sm6r5glnzfGNvkIF9GOFqYQgOCphqVJACUkJvusKDGxy
S1VVAZAVRVtH76ZyBEtkifTCQsUismJ47xCrRVHoY0xECqS/sHo83JO5XcqqORtYGUqiq48LAexa
JVhWKnGmqCPNDzTFxHpzeWP6WNLYKbD3T2G06k//8+yd8T0d/PFdH+7Xxflukj6aiiYEklXqqBYF
c/DBeFWvZcz98CvvkV4SuaCwBhRq5LdlZEmbGbG0KnHoJrE+mwWsYUals17Didkvr+fDbKX0ps+T
3IdzvH3BG7O2ex4MVYWXHUaI193euBFSwmLbze0tCKR7MZw9oM0FWMZS65djuqozPRIXSi1dRh/k
EbPpUy8lQVtP0RRFv1Wke137M0ODHKzfmjNcMV76Dqi4vmaKlnku4C4/FVHm73zGrICryGkmOV0Z
PVFF17317oFJZuyQ5B2h2zO9DbKsVZg6a01VQaYdZO46kMytS40ibo+qq/PauDB9WA3iS472ZtJ/
45bWchQJEuNpbR/p/mN61lMGWtftd3398Hp0tJzndggaWuixRMyqy57/9/1HdOl3SkCu6LgLJ5DH
gtnk0D7Xt6DlctjvdGH5jB6smHOWxK/AE/92Sak7dkoPCj+uBsKycpy4U6y5EnWpB3uJ2p4KzQSF
yiN/gcXol6tLr1R/QMX/hsSnA/VxeI6dKpsgUeCK3fujbjpcQCkzsJEC3VAsu2BVRRoIIZYIocl3
VaR/wJTNp4YbI04H0ZKKYYhdp9rZbJ9EfJ+JX21wZmaO6mW4LCTDzQv6ZItNjpIZBqKDBcyCKO4O
tW7lj1SbEdkQ3AqHNEZWc6Bo+Z2Qrm+B1O4n90mFGLHbPtf1CiNBxcYt8ZLiePgEjI1b/xFo5xsq
2pRRSZqW7gk3B4Qr5eQBdoPDerINUPfb/VfA42EDLf1G+Rq66zElejoVLRVLK67PEGvGdS5ngHP/
MMi1FSkpkLuz5qkf8Wf9vjYUOTqz4JnX44L89ryCLePn0zDmKlMgvIP00e0fo7g3cBuT/qsHnWNe
dBsXS4/t9FWQRY5AQw7/QxB2MSIXA/QR7J8GfG/nNCSEcsVQdEZjQ5Wj2FimjSoKio5QBQ8Fl6K0
WvvO/63DcdVLaOeUW8VwssI6sdLvr/Xku409FNaXe3Oe0KYBwcsjuTgAx5fZEkpWQNFr8iywOnXY
gUO0IJD6l4ADgGAp4N+eBecBL2R7xIIDzKM/pjcow1KWCN0MUe4oe4hPACDoMUT0RWtoSC+cMICi
RDtdJqeudbtrhXlo3RFRPMr8dedie2SgHdjN7qA3fzgHT500N1+FPYHeYOaHEBFG085r8zBdWs0P
9Aqm16deE1936jtwsS+ymSGHBtJ+IHqnzdjJtrGUZ35A7Cu3e9gbXw8QPBZGZaD9HWnfEEIuGzhT
xkkzaVwxwwBEWPUygOeBHCTmrCaJ1C0jIb3IJ1tBvdT8Khc+iQhVSUM7p41zjQcckA57AgZt2FBw
e6x2+qWm+bz4nbJmC3JnO6vfTxfks7bPaGdma29VDtBfdu9857SVvrlSonmhgihy1E3F3RktD9a4
cLnrpXanSnfvZIozQCkK2hTmfaBp0nMJHurZbgQOgAJkduL76SpfbVs28OnxZL54o+VVtXWE2GGX
tD4pnbQVg/GY530qUh+RsA4UGMVeiBK8AOfmedYZfn2VUYQYS7avik5ErbP4ka3kjPzoSu8xwbcT
5G65hBqNH2Tc9tuA/Z8pCKD4TBrITdcGgPSkdBXFHxurwM4djQwvzl6iPYWCjVv7R2JW4K2D1Njt
W2Hr4XHoz7cIlB9+8N5cKOR6WMS/bu+ewj1P6hKvIB7KoTUmJmvp1Npgvb6DbvJj+PU5OIvSHbz0
ZCqDd1sgQhuBDwLThDvuWPM5EoG4PTyPiJhBbQ35xRcP12zQPEs+FozyM1nlegIzEmze/5AhWHjQ
qPw2ZffhwRdw4A6vQaquzAvLOWpfwv1wfLn1RjVi3Mp53tzWy1jVYos+aiR1U5JeYtJf660JY9al
lItPqrEt0Zt7Dh0Y1xzpYfAJgJ8zgsIBdYJz81AKMlHObXaKqgf7mvJuo67vDIKglRc7a1C6s9/K
hJ2L5oJ/Q2RW87cqYo9pE6Fwz31TKira4D/MB8wNa0pKUqe1na6d3AdQxuFMuqNfROPNCgTJgZVp
1eXtVLHGw7U0c1ao5pvI1zRj5/JFiY0Hj5HzB0S84km4/4+Q3jGr2ffvsvmUarxBHV+tXmC1ssjT
nbj4cD3odrL5bQDYbKXd+Q0QAM9HLiR6ZrxH/w/yaLx8EGNrlUp7VgKFFwR0JMxi2ivTaKMr+k4E
GAAxfRDljyGlMg5K7iKyYeRZ9emwPUh5CJCI4xw2aLDy2pyyZjzxz5cmGjd5xHpfHhLeNNMmUn2F
WzD45sPLqRF/jZymMcSWabFAZBMCg6BEJ1HpisJMMWAqojOsHrHeRVEFJ1WJIHB8X2B38DNjmPFR
SOWNUDNtTXnMXF9FZtAFBBQcRRxzADiJgttwP6haMhjgkYR6Xgo34ozSmhgUnpGmmAmpoA6PbXu6
YI3EkvCOz6ZvnBznX9l6uLjP6AzMinVlZgq5PZCGnl/CaD/kfbl61sKTSKyYvl7x3fvAtld8br5R
5W5sKdEP+kC/6ODof/jZ25M6MDq/fxF8wwB9TCi9tOPiZI94c9uYg15Lx1i1q+BtCi1wbUKvhqNS
bo/TAvVGF5dIAYIUdgIopQlhb7RACHX34hlNGlzsxZrt4StgXajRoP9kg5F4nR8kosIp30w1LZTe
bxgxhRV+MJx5hGvjx/nhzN3nQe5rmEpaNGzXJeinh3G9wcMSi0Ybsd4ywRW7/yZgtCBW17x9LU36
H4PvirIyrW00R1l72lnLRX2xX7STbMCuvVHI+EFEsbJenYapcYrW0wC18FkiVHfSkobpn3ZHPMqp
PTIQUeEs+j9D14+HYWkCjxQjJyfQ8RO3mcqRguf1byOxIm8mLSNykmQhD8LwsYWkYUSBfinMs3Ze
NfpTN6U4WEkV4R2bv9E8caTVBbtK2EPxEJEOqA06U73Jf6kvoedLLSDkZgZaMWoNJjmjguJGNCvv
1gMz198S+Ppa+jaxbECWOuelgDv7IwN+cpzWyiMe8ZPdxsj23VPuCN2nPhe+a8/FMbkF0Uxqbzap
mhyC7CSQXO7tzwQm9ygEulMiSjS9qlouiw0HHUiV3T1qGCb+h3g9+3vFpV3q99pssSUVJNMRCDm4
EQGrlpCTXC9g4NUHyxxhlLp+Ud/kt3hQlVFA8fiOUTcn4FOLAe8kVM6T4tc7R3ea8NcqMX7+mhhq
QdlOO2yC7Tr7aVUE+1qnc4THouVGMxH3Wq1N3hcwNUAhqZS76/0UHzOkNg893jLLAU3YP6UtgioG
gNvctQA/Hh4sxgk/Mj95FHzrI1y9dpVSMi76v8mfNYz7h891sYsWd8NrcXumtzCDjQm1JAsB2j1q
hwaAVqFLy0fDdHvIKio1oVX6HG7dygo8t3CbjroF+/+mPD7u2DuWNH8dCtAKO6RDHsTqXdY44g/d
/Pmgaxt8fLMQlCviNtQItgy2AlqOJnRa8PyVjNb9S7ukCIPF8qm0CHk3TpDkiv57L0jh5xjGg+pI
B385xS1D0NFCy0LcA8VM3bBZrZovfhh0Pc8KbR5IWUC8lMGHgl4frE6NTaujaqedx569yGbGNuDP
7ILVFud7546vaYtjiFqupUkBZlwtgrD+8RN84Hb602nI4a0RtDDfp2GDL9nd8Iuxb5llGhx/Ep8S
cZxEAg8reFvD4DAVGLalnKAYWgcc2Mx9rHloz9MTURHmIwIXwJDdCTRqzQW7uea3JqF1vTpQXkR3
ZUvLubrYEgRqByiDQuzFukWaBj2xCgd996P6a5k95cYdtf3MZ4pwUuTAC0P9bT62ffhsTWH5xiue
OoanYyNXzpDXBxWS4MBLkQw8cX5dnBKrmG5jCJVIY/Dhq5ok9zDcE6RKSo+aVtadahpA3g7leXlZ
6LU7qPFbk3ZnLgn9zaZcff2uw1ROMdrtGyZL7JIy1pGOU4UB7KVr7teM4tBG/zhDBPhmqUDehl7x
Xe0Erc9HUMrM+jl5P8Q1jnGLp0MLkTfOpupR/HP/uBdFkiKm2N7d3gwNv1lynKc1AtoFfb4aQUN7
J8/k4VeZK3hG48TpfWM/chmfoWgPWy6/oJkbouS0exOa+efceVdrxh4VOGr9Cva50wEiO7qu6WEt
6eQp7PoGbV9lALc+u8qd6CFjBb1LjvqOfzr3QU3NuzRUIfrDh2MKs9kZaDYpSvj2qDiOvdvxaRG4
vdKTXXKOEs3R6uBySN/uwRzSgQRovKxILDXkoqwmo065X9kT/6OX6F5PVzX8uXD6v53rDh5svZbO
qeMqIwBjqIwDtWzX2pceVvCYr2HJ4yfQDSaDL48gF2m0x1/ZK8nP/sGvL//q/eVDyOLO30e40tFV
WixgLejAa108EkwoJ5L321gmNcJS96cZC/oppoBVTTEIskoNw0qUItV9EG4TSgr4jAwNHX+N+3mP
AgLVmR3J7jK+FNqDe05I6cYmwLX8IJ4mRV3c10y2mx3o3MGdb9vnKWzMtiiLlHxszpjvXLRxIcGh
rCcBis0d3Rc6297Gh76WkxhT2OPpKBn9eOCVXmFuCMcFxTsYKs+SJka3i0rswkHj7JW41z52tJqh
xo4YBvCRMA2PgAaBmqZTzmgUqgx2JCwmTqOmGFyuKhffkNpr10mU5Fb918DAfAjkLEX8NHmch94F
0rz/Ce6cWT27cKMOXRZYeupLjGF0F0KhAhUUWdiumANdsTjwZmH1iWI5TUpdM7ZD2n0DbNTTpsUW
bkPLxuvjkcrm7AbhmG8CxS4GMheeJd5nvwjKMIRWuy/NYUi7jnEW+9rVXLTOyK9Ef5saYvzWbXgk
otjJpPsCi7B+EPLfoH0g2hgK4JgF92FPhsJ1iOpjAhJjiJJw1MCj9H6t527oyn+SYIOlyMz89fhz
Qmgqtkr5fNO7TKZLxWhkSxrgZA18VUDAbsLXTg13+bTR4gRPhHMLp8xT3EcLeQlVrGB9UMZTTwhe
uEVxBLDvXk6P5MFWadnRIWlGO8yYh8Xl7FXlhE1qlNGSYBvtHHnfVm1rMSDClLU1BNNfBLz/3zKA
lDhQNz53Gw0YrxwI43fxvXSDgMfN3cAg9JMkWyNPN1TBzUvRVPauObbXh2ikbXjq2slOka/IfYdT
gK+cl7+cjY5F6Hsk1Mb6gcIkKH09Ji8qXcMuxL2gV+LQ/FR0rU+WGPjaLDhzNp0nhBDqVDLjTcEM
geByZzWi9b7+2W2HaYTiRV1kBlUEHbhxJ2SgKvu4nPg+snZVK8qIvv5uKzmw6awTizPB+nKHmKsv
q5tEGba2Qd5diaQlsDi8Ccrv1IPjvhEb7cRyaVSPSl2QyQJhwINDRh6W06QKjhMP00F9I3hUJqJ0
zsbHpS3p+dP7r9n+olb8nLyZsxgzZXfnAPsBP+hTyOLa+sfNn/5arYAsBROSg64/6+rsX3J4tKpw
Mg8RsTqpiGnLPPwNRLITrmzwQ9NQAh7vnavilOB5yFVHlbm8qwZIo7J7Nkcp7iEyYMSCd26jKUou
JgOdHIwYP75sIqfqvuwg8YqZ9yucpSBNXBmQ8g3Ahfy5suw7og+FPKBZy3rAmZVY/Ak+ZBQKsdoN
JYpl0yB8vnA+A8zrCfslCYMgHsQmdJVKYKzNyeeLFf4fCdFlwQXtwPDN/Arm67lxF/hM10Fxr7MY
6x6uEaJTIXrOSfNyinuQTtSp1uzROg6wPi+QtR0srDDrsbGETB0I43V7CIs2k/ae7G+l9oMhEZLq
c5vSwsLpkx5jc1McTTlLxhgttrRZ6t79+CizWN2piKuw2/Qo8I1GPy7LcheBngSxdypR3tCUWRLs
+MisiR+TRY9Q/8HhyczI6nMKgRaG1kWsWdP2KIfO+WYDVw/yM85uY1LApf//wXvGgMwGUpd9qFdS
l5bQacYwUcuEfraozGNp5aWzUhQ1Hh57NkCnWztSskTUv3z86JWrc1Y051/GuFanJkFQ6GH2qmOh
NvWIy5sk0QsGzNCLOVqX4IRQD4zxYqWA8NFLcaKqfqmWIPv5julcUTQBG8l9EnImHCB4Its9n/eO
9EJk3rEvL6w73lmoMhXiluMg0AFt4G7G4/1ISnx+bVYgcIlERX7CocUe47dJDStXeKWnZnuwnmwG
Ro+1i2bZREebdUSvY7iTGN27qGF4qEQICGQZEaDPZolzPrCkjAtwBxwvpJMIc3qvs2LplyHV5uA9
OuggCzqmFISn4kmC1JViYqHUtJgPsfnWEsD404Z5N/gVDT/vJdCLJOOOhPgTptEJrdtQhOnmnqDW
3R05ZwfQiesK1+0XGVwHkZVMOfvm+baKfvmqriNQPnQTgU9HSsHOyuqhfhnePl742zDB6atoHLm+
5+QPOIBssTHLq2Lo6IERRRPIN6xAglvtcfZnespSJyIs9HvtUMuBm9M2PQpXOQYi0Ky1S5H1wzPL
O+pn9gjmP4hrvaKrEu12ACCsL5csuOIeNLoZm5M7U6bO5mNZgvBXf39qx3IIQJHiqUITOnutKvQk
A90zfQqboLaZ46c5mvh4xUC2tHvGOFfWm6UtKV14ADGKKNd/xGZ8gamO7t15ASNN+cC9xtWoZY2P
98zHzg9l/ELwFWL26kBDHytrFDghrWOorWqgJ+hBtUleKuTu4fR3iFYKoA1jnSYORCUmHmLaVaBq
7lsuvmKfrodtcGV7Kdo6n1peiPhk0mTTlVTOY+kUFehkEnkYzhpJQUp4vfvibPFpiEs2OpSC7UeV
Ozot/7V11C+iSGeASqo4c8SBRB211l4LRd+P28NCHR220ZcKsGAMGMGAhewP7JknjmsX7y5/RUkJ
7Obto+ezbllRXmoShZNNpAXb6Zovh03a8uFaus+qSfrAPNp7hlc3u+zwgjQwSlUttFtJirhcQIuO
dSBni9CX3JVD8+RI1y81V480UfG2NfQ3ZO04fGi6byospP6TmlDnDYMlst7sWflxOV6cOSVB8yKd
cVt8LWbYpkTBfzSPgBek6GNhQy8orUj3FZuXMII10letTl3bTVI7YXNxfUCy0CQirzx583r8CA7+
BlL5ZYywFTKHEm1ady1AEh9tbwUraFU6Ix9FVMMWKhVMNdDxCBnt+MXVhfENDjhWJfPLoOm5OCTK
sbelsKJpaqhBiFRFSEuBmhTItk3iFMBmvM2ayskKsa6n86KQacN3/Ulqbg11vsifa1iH1xx4gARE
u+cf32uP30RAYW3n5G3K9W0pgF9LvSxMcYrrQQpQLTEFWjQxPJ6UFIA0VNtLHUH4a3X7bPv4I5HA
x1Bd5XyUZfhEtZGIH4THkqorW4seLsxQfDq08QrU0Dp7T7jSUcbdfQmQcOuLXUt9AER9LRRal+ww
rX7OhcDzINtSglVBWGfd0NXrE9NfciYtG9AncTN1Zum1pjmZxyQyFlFP60ih1WcBvj1QfzcAu05d
gxg+FtMrA6jInVFk/a+NlI2Prg8iBUP3D5KqNmXIbbnhjcB2X0vMO6ltToab+NpNMscUBr6CezUB
zCKK0oOAgFwOAK9zQKSRay+n74eBuo/g0GWylH7UNpMyTDRyDiSlWiO82gT7QaIiXv3LwK/+FLWd
PBNVSOKf5Kq0aJ0ioLR5FhjpuxZNKmoenjSW7luzqFls+y7DbFQ7ul7+OL4IBIcG5bxNDGwhJH2L
lpDR/QLqTC3B+OtB3850JBbeYTmHlU5rS+4R19kYHHbHUzWiLdsdMQzfHwXlBsVr86cxUB5TyKPI
P+0S9h1q2xZp4QrsQ7oqFD5YIM5la+iVSbgz33lCqt8oZZQCDTT7JuCNCNeqE+HNtjgs5IhqsO/q
I4aafARQhdYNbm2dOKqJ1Chg5tpwQInUkLBkwD+U5qnHXozPjeAnlOsJVxhhc5K6nNfD/xaK5BAu
dTkSiOgF/U2uDDyDKrVS5W8cwy4xhT8H1W5/CL95V28XCId+3XzYhDUfU7sHCuCW80mRofV1cdno
JC8fP9A04gA1pZxoYKkIxYh3XTgxc6r5rVmGD/0eH02cFtcGxBTaORpDvZmnTMy7znCBfd5FhlTo
x5gyj1ORxOQ1E8BXLCYu3SwO2RyN2eSQMZha9gKrThDzdj67RMpu3OQ4kfQprr2GS88Yj50NY8Dy
vjhvqtbrBe1ZFpN70rTIx9yaJy6PzM540YjX46bDdb1Bj6c9Kf2il6mRbhDl46sOHA7LOUNEYM4E
2TgfHFcXyu+h/vdL6/iTRP7GLRnmkniPu3PMI3IYr9sWsy6tqDJfIRsT57B7wHkaMjGvUdhuKQ5p
wSOriS2yxxRrxVbRTnB1wE1UFO1GcWdverMEIRGbv7L9Ch00VZS2l8wgooutIEVX8nsO1hq0xklK
b2hIv8lAKwaSvAk+32VQMNykNt4z6O63hlh2Rf4HA+uLpINf66zO144G4zssX0JVfIDWxtGgluQa
nUB/6AQvdqPMsR66s2mcpfGwG6hGHJ7Us+cdh/u6LxaNol3/gD7/KBsX1CIsDOFxN0KfAxSG0kWk
55TCYSJtDZhKhf6OzZXj+OhJcpHwVIxmgqHEzLeMoX8Rd2Tlw55s+jWEmNf7DjB7hxFCcP3dDbOQ
ufFcXMrKzVapO0HZ2Njd7v5biOfq5kdgaDgyHE7V1yAi88mQUKZX+jGF9whMmINM1xAbLxM7QIsx
ET14SHxKeLy82kZoySOhY42CwbmXpUjMYryUWViwfvWE6LTTzuWJ+6MIX6vjz349KN+F043gqTKs
pVIn6c4c0et95OFg417e5goQVzjh+11C6bNa177543QhYsWT4g3nAa+/qREQLVDZpDuoSqVKO6El
5HavKf9wzXvS2UsrkJIUZlFBa5Wy/9C3wHIry/uDnnKZ1xggm+rIW7mgdimZhKb+6I0u/WAj6fe7
4m/k0KTHCsT4W/iWrbe60dGB70B1xBEMQh45zhfSsGVS2nGR7HEzmYEnkY0XsSo6HPrR80QCPwCl
d8Lw6qyCWFFzqt9sJPZQD3HDP8twQITVY0G8On/OhOIy45WhLfwBtw9Fh44b3vJP1dzRGjFWgiBM
KxePh3hx5BA/Rl/p5llBKXhrFyL+06zn6bUYoDuvvvi9Rv/c6g+NqB08Abzq6wZEPZRnSh8sLzYw
sCnbE3gduPjYR3WHzPhsZ3VJZqM1Z5B3J1xycK0aStRW/3Al8FvHxvu93zj/ew/WqJm8PN4y1M5G
XzH/UIvRMWFjsiiHedqrBRiS8XeM8/bLNCIYXHqFAVbZj89dkS9i2MhFo6Hjsh7HAAasV9HiSLIP
JU5qsoWg/VpeS3N/c31YjS8WFJMrWIKeyXrKCHGmsRU909zad6QroGMH9Xamj81lvsR9unbZ6NEy
nWINWl8zp2HnJGite9rOYv35XThtFVTzdpoFZXuImddWy9pKo9060c7G6obJOTi1iYdIn79MtWMB
foN7kRI+PhH3NH8E8xA/2eeh3oA/CzERhhDAQSKRJdP7Neot6+fKdcQYV0FG+8QQh019ROsRYwgR
XQt5nnNhetKxqhH6R0U+0BJLwMdbLU1WlgUeP6J5XNU8odhOw66ztuo5wkSuL0B5qMcAzNdkRB/1
kB6cDuwMAp5cIZYePxp4Fq2YU7YYTjlwGrh+z5bsccPyIYa0ULFsDDw7le3x61Ljpf88MFHEOPBo
PVA04ypttwK7lohyNfV7dApjMuYxVzkugA/LOKgPnUEyIPkZqWzmLjyVF7CoZ06IJsn0jhTK9UxM
JbNWxGvcB7tjFPdDNfLcIMLDUd0EX3hJ7792VhSSS+I2jCkGwixknP9U97bTvM5f+3dKfL8FgSh8
mjAcBw3SbGEvuP41TSR9uaLVNccISk+qpWP6Y/AesWWQs3BQ73gwh0DoZ0OSF5eymWNWFl3PWF34
ndRJGtVMzrLWsa3/qfy7Gajw5hZUTcKDMARs31Rky2ZiE/Qpi56c/AG7PLBpSF20zZL/YvVFk7wK
HQ/NUKdKcOyC7Sk0il6vUvbdV2wr0nFASXMtl080jD5nhgBWRW4nHm0JDOAzWbqsFvII5/tdBmx7
0vaAQqxgr1JzS86njr7HOyVEjcJ0Yfxi4FEmfGZ22MTl8PcgFOgCDtzE7pUk5WW1+BnPae9WN69G
CX7F7T+yQdl79/V8xv949QJ8gcm+NbzKoBFsfs8hwMcMebJ8RlTmKbQne9pxnZ4Kz3D1heZCVyAG
TdC0yxAqSYk9acN3RxPiMsomy5kcdUNtB5otYtnoy8ZI9rf7NVkf/m72gW0hLPZ6fNyYFcyJqrcr
7Q1iqGGqbOWeQvhqjRKl77xsErBLB0FkCvdFxKY0ybwby2IvsCSsCd1ml/NHIsqib+pCIMpNWW/u
QhcKAXRMDIYAk/N3bnXWDXyAuWdA34z1Jnqo3yL52y2m51538XbpeNBYbW4ynAg+QlUEqOWtu7ry
fsqx3/BnAeVi2icf9T7SCcgKINh2y5TThibDCHlrJzu514akYoQN4S+cxsUdHsuxyNW8GW47yBf7
OcQc8yOKB6WUx8e3oRr4EnJOWvdlpaElS8D6zSxqdI1ZWlkTz3abg9Wm9vSSvioGxL1ir3Vt4i9B
LRSj6ZqSjkSJmF8PBd4JkpVCTp1AE4RqhQXD/53BxdN4vgo80vZlChCFygmw+dJmhbcH2aREh+4o
KmZgc15wxW/Vqc2If3/ShymrxZcwjWFJ0wBU216bW3VgPXD9FEtH0P3wmfW7LRoT6L/wwdtug8TA
jy3uWRi9YvNcjqLox52ErD9d2GOeyRLpsnenyo7quU2e3x1yRDSR3ghtJlpIADf3pYaqbPpx/fGv
+Vqm6wU0hBOKhDsuQh0XkaxrgPLmx6LicSGfpqSIBVaVri1vTzpQ25XhRFWLltuSkacQA8tXn/F/
q1DfTwRGomkqzRrg2caLK7lCfn8gv2sTK4nGFBxkF3YVs5m1fSQ8BQBpmAc59PE6QXPrafbIZnhb
pDjxgHruOqs/6QDVcmGtWrBaFTRP/xpZHgdEDwgYWfNxDXMCnLdMRDxevjDYe7NIKX1vbsdqegNM
y4GzJUdVyJiHZeE75tJpos4EfZ9kcphIppQBqzenUvHFfgVMkKK+uYrpyu63uHkWvTxD2zf7cfCP
BwkIucx3W6gC6yjMD8Kr4kuVDtqWjBlYb/sGXmW3jIRxFqdzMPRf/xqeWSNpA9uUYTLmh8BScXD4
WlVzaLDZWlqc5txzu0IQeG7zOA7maV53WhncpEQZesKtt7YirGaZjxJWAk/7EJ3H3X/9KCd3h1Ij
C2jG2XgYKb7X51pGC4bxY09RxnEr+BqGM9Q5FHw1HyCW2zQuhBqyk6vy/++e66JGsHyWwuIsxCV0
tKF30BGUzlIei4qjPQk0epAYukyPSu8vPyts2xC1kWu4ZyKoXcbY+gvrHKV6v3e7yufDI/WSvL2k
evOoYRM2KPbugzL1b60AiDywHLxJ7zqSu2wkeDxp+w6OBCy9rzI+vXCCksN7iV4VnBMwDmNMjmwm
3AnqZBXUWpQKog6s6FYgefgUTqWiVvBNox6CXT6i71nLtIwoylS6EXOvCC/yMqC0OgiUokSQNxxN
ycmOHdjRdMYKmTsPgWdSkvXGwvXo6CpHiNxPR9f4pcfULnzU5FNnE4TPlJidtbuUVQ8/r+k4qdcC
Lk5C24ICQmVyx7B68E8yp0fZE4f/ztp/FWPQcyeKOgHOMglYUzkBRLOKnpU8NjOkxUB/PNzHVF0e
0OG/wdyf2HUHpcLYIH+K4uAHuiIpij/S6Xrq7FzEVrQgNVJhucj4auS0lky43i7SlirwUhjU7LrQ
SOex0+bxBJBwc+gfyG0J8wqwbtc36YdrCjhhbPQ0pt9yLkZMkRxhSRBasklCJhnUGycfcVj2gP0i
w/FDaM90AwjRaX1mzDSAMwMtFHTzGUr5Bh5BXqwtMk5MrCdicq7j9A1m/vhUgoFnIliyE++st3mQ
8YEjq2BFh1U8UZnlj51S814CBia8w8KC1qvdL+YpVwIpZQrPaFyPmD+a86RHeuenr9hGv2WKXQMV
L4lYEME5OGIvTsF5KwA7UQgECaoDdIwQOWEGMkrVpFSoc9IBVGROXeyj6cAmLiL/t2ndDmBVtuKZ
RebSpqKyS8zJXqG06v+a6jn4Yt7qzxDt9OKmGKgPXcIZxtyrY8QAbA60fT0+vZ7o7GXD1J9C1gJ3
nxF5fmxRqG7ZdhroolJrhMZSvOivGgjLIjKDabN4ZHkMTW8kcDyJSaDizPDbmR5cDTL13sTd8h6j
kDixWlY+W4stRkiJlhdB9iYgnlPTld5Ks2fQak6lzhS5QuunjfEP88o+viNVJ28rlhCtSZ26ywMb
j5bKIAItRcAGZpIQpKDhssmiUUjVT7M7qwZ/UooOJlO0twtXvh2J8zKei90Zo8jKxLMdNCB6JifS
/G8CyLxiMalBGeFp1rAPon6Q/9lxBpThsIo1Kdj6qD46FZzbqoIO9KU9UENYZtJLkFJDNtVj1NuD
SHpBLYC9RrbRUDGWclPFZsYJajSUwAbqkCKd+dLy/B0j+c99woryJp4TF0AVNzWtTh3imYC72fUg
PwN+syJehvwzusdNTqAII6b9XSfKIkg+MZ18S3HI/F4GZhaSCRINzET+dtHG2EFLRao5dIZskD+9
r2FPKvhsRhxiIE09yZWyBz0xmliGADxCa2plemQyDuxfLc8qlDcbT9wrc13/CtzW0riOu8JIw6Ss
oqEFQLJlCV3rMb5BGCxjP3dQBWOiEG4/ATd1oM/XBDmZW+vmW0xGg2cYv2sjWN/kMFuAP8iKJG/2
X4XWSqgwuLyNElFZeUaa15wNZe1msSgXFwKjSLGISZohrasADzdGBHq+Bhav/eifTJzG/lL04xck
/cMzvZvmwOtFFAqhTzCsC7wyRqzrALZsQkkazWst0ZJKJ5IjXBvxWkP2QrnrzN8KmalkoEexDgIg
rXIGf4nIMrOr9DW+bGS8Csf/p6RixqP9s9cE7gEJzNg6vZ6y74xfUTLgN/xwwuBhUcAlrRRHgM8c
WXFiXBH5OtD6+SrsWa/rrqxYb7lXMyU3/Z6ZubqbUK9eM2/yT0s4QyNMGh3wm8L+wagCuCPnNcK9
szsw1HtQ9X1b9e2+ubPLYzEB4aE7qwHs2fCevUFndTNhSubUWE9oKdArYPmEKVgFWgI6tVnncZsJ
tU+z4WJ4TPRYwGEKSBF7S8mwzePqPId5IupJopMvagETXNO6PATGBLFogh/kkCKVNe5s6fnZKUax
qKPfLHt6zNZtHYz5yGLv+kndoFEyEMOyc/nQjEozqcKIk/Otg/sC/2FwZITfHqvcDXsRLIdZd/d9
fEtwtxEGyN9BVsIu5Vlq2/MD/qgXRqjgYGFgg/LLYKyJltJ+mzKpc65fS20OwjAHRvTURpmHAZXq
i85hgM6D3uch/ScViEGgx22Y/l5tUgFV4SeLVATXU7o0qOutiKurYB5d1o+iwS3k6guIwP2hdLzA
2puPq1RHDSTGzljJG6z6JEA0/bH9lSyMWwtSrazyAaWVCuZ+eLCrkzx34qH6gaX7shO4scVYDyYX
YbR616DCSgsCJexeYslizlg2GylaWpAUbIBFbnVExlUAq6bU8xFtGXKOfIa/RZ1mJcUaeBcO1VWU
37lOvr3HnE+BhZIz6wE0yH0gkEb2rix6TEjsBlkOekMQ6IXhvYLeY1V/nexlX0yp+ScUEch6XACX
PTt6jP74xQLdf7APa/8BWYBaJzP6dr9ztm9a2QLULSgJ51KDRsmINkpMsoyws2S1V7e5uWm3crf+
zyz4DNbxSXW5KogO+olITySdZDsuzRvP0iIQMNHbTDU3Ohc+/c7Pjgt0+75o7VV4aJ4C9Tsph4Te
ZzbVBqKiWvNBhUDaXYRanlKdm3Kj+0qhMCBLeaAX4mtcoGsDHkf9/k6CmGRnhcBEDFqMc4ax03HG
uDb/+LpiIhz222GC+bYbQh5yIv8NZeup9ck9XkenUb3X1hCNmqhfTberA2Q4F1tMvfAIm0ThLfgu
9MVSfKiALpbOgXiXpU3JN6bJDmc7HBoL7byoDNtlFkilkVhL6PUUcnYkoE7LoBJSJ3rpGUHriXC2
AMnD9+ilno6LdESvoN0nVZUkmXpSAzNXU9AU7dP/3HEtlGJlBi2DfFnpKvntsjIeHzyOZWm9FMWb
Hz7OnTz3hxsHMmSZ3/CZJvRyWdHMpE9b/r2v7piKsvVLKJNSIPZRkJ9PxBaBh5ORX32zeEayD2Vs
SPphSfbhOxZ0UTaxEreHg8YU1kVQbrgWG19vNpYfjbLA0gow9p/tYWTZMpwamOJ1P6mQjiN2jHDJ
0L1HtP53YBtyfOtYShr8W1sFDP6JBEgWnxKYeo0wx+ZFBp+6nY+x4kaNmbut9rKPFl5hn2LgPzEf
ueshzJbnkecp/TY7iy3eGJKYuQwUTTyF0EPnRd/VkEt88KnWReX698rYj2hjnrmQriAy+CVoJ4+I
LRI/m4lDI0IfzijCnbU8JJ+DtOCu06lo0sTNS2OzU8y33sUNPTz/Dw63OSATHsIJWKaYy8ADuzFt
mIORi4XF1Wl5nduk8WoyTXN6e6m7Um/gMtyTWPJISeXcSIk2L1HIQOV8XTo7cC1b4bmalTu88UXA
+p2/ADKa6/jmKz+FropXnbeHjcnJor/jzAVr/VFB9M7qDbUQYnR4o6Eo3Qd2dJUViH7LXwlcDjrv
eI81hrBJK/yFAPr5JQScCNeiUlYo+DiIJuKzNtiZVWK9sJ7Hd1Gm+lvpJNA7czc9nchUKlbwDcZZ
MFllvZSRsqFPuaXbe6YXli8PlC1i7aV1u8MMvO1QwOhdtRjwWVMtqjeSQVsY+iNRFZ+s9JJUUAW3
RQShvEaqYiAhzTAuRpu7X42moyiXSSA6UZVvNLD+H/QadG8MoUZ9YqOBwdoqowWCd/bKkkxv03JZ
Ng7lyLBGEa6JzxKW7yhBKTazsowmO2/SWdBXS64pLQrGFCJihFdjuixyFwBQkTFxaDpyr6u+ESLW
tNdsz62M/tqTbLT8ykn3fZwAufh4vxZ+K9xfRfkEj7IhSktwBCxxYPLAhWCjkvT8Xa3A9iHQ0KTS
YDfwxXghUA6K+B3Ifh17Nwj7XOS1R8KHVG8TWcG+pms6+P4LAbGM4jkyG5Uk89o6lJ3CeDAzJ1Jn
tuQ5UtJ9ArtJCTQ7Bgdf0ljs09LlnML8d5CYLMofa8zs49JgYVkD211e0IjaZdWZ1OmNw1ScgOqZ
uiq8iUm5dO/olCjvHIvhOjWv+wymdsCMzkUsolV5rbTS6vhsueZilwwQrWr8OqBUm6UTIDUExwMV
C957sNa16TwboLLqg+hkuW2HU/wIlsu43u0rAc2G3gwDkCYBc+rcT25k9WsdEL6cSm4+5b/7sCQE
zsfXG5his8g8TSPzF55oKrYCO5wwQQr0q+F8tBBJGEmUBHw7UsKUq2kaTXqnpKXfDNcxh4h2XW3w
nUjudLOn+r6I2siLpynxmbbg0Pzz/6TEFTn3ny0pmKH9vbCEtZoX65rUEgykiDyHgZpCo5SKuhgB
5I+kooudDIi4bh3U9KvUz7g77GSeZZ0KQubgznaukpibOYALe/wrs+MocojxR/f8KFF7z99pVh/r
jezRcj6Z2/BOQW+SDI2RasPW4POY7Nn3S21CBa3nS7tTdO19DDZnFe9J/plT7V/VbwNnz8GDtjJA
uK6Bf7oRd7/rz6gL+6Sg1BB4q2RTBNYjnSa1x5bdnBND2EBVCqbH3f44FVqXodiCKFdzDAlZNWNq
O1jdE0/mkPn7y5D32dmPpz4AWzyS69vRQtqv2ogeEGdXZ/b5N99Igar8gnZg1xea7NC5wfj8zhM2
e+YEzObV0QXISufaeQM0iv6hxy+kAkkgvIyCj+vJ6cQCGBYr3ubUbGMzNxvoQ/ZA6QsnjjtXXtbz
t+8ljPRhxhT4or7eqViw3YGjzp/Yb6DLfYfcFHvSWGci14fuAgTjAT0qAdSYhHwRRYsXNimLTAlR
qOEUyp3H/mpE5Xpe+Pi62fQRsbcJnTEPkVVBdllOwvP8GRxpbVTzCOVYE1UAaNNwZg5WVCxS2FK6
z5RU77U9S+euUBScL0P5zNbUTLiSE36AFoeG0AaVR/GIXNnUmpxt22qIccOyP+dhfHStfMAuUay2
IxXwORbXKYaIsEFR9iQ0wzxMIxuxeblONShA5MNEg0bjOsTjjxpaYATWC65ANbPfJ/o85nn5oR+O
PH89WH5amh3plKiiojRSi35no2SLqBFBg2nYYMUTXVN0B5cK/NDA9nL0ewHaHPnyMz0lyEfb5U3j
KVR9B5WQOWadXx1Fx9vf+SmvFmEcIwIYI6RFQsm1/vaxT8I6jn06xfJb3zNpdKOWEHVoV1Kyheuq
oMpD5nUsVXf+6wCbi5Q0WsK/xjxe+nEhR7tVv6e8s8RfKLjRTYNNXP0rNa+T7fFk42BRaXmxOp8j
EG7uEvHftj9Uk74iEW1Bp17lAnPONwO36fHcO0yRXnQRzhH/yTxSt+CRY6gb+OU+7wG/20NQ9LrL
Zwp6q97PFX3LKEq6/m++f3dblxNUx9LOcelUK7G4HPCmIBM7z9MQGj4sT6gFU8fu0c8RGQFBL3UU
Tw5v/QSUhFIjyoGuTv6bCH7rZTkv1WyVCwePCSTVk8E8K2J73M8PefOb3W6YPOOec5xtzcSKpT7c
Tm00vkjNMr1oqQLrAIfVSn4v1Gzyi68GQEqd1PMDCfpu7SeU943mSP+6MfEna7Nmd/5pVfZ03tBu
MM7fQdpsNvLM566sRtVcaheaUWgTsQEbQrfaHtZBWvo9wTCBtLzOVCyajmRrF/7072XjdNu9yCDj
e2obfUyHBcVqz+v8M2WZnaGs9l0yJEUayRdF5KEdS9alPRI093uJuuThlHK+0+yTI+TIw2Ehxttf
VYVZnDOJu86fo4m1X5X0P+LwZ709wDUSR+CxUBkbk0cTqJl6cuTv1V6S5phbb+R7NoL1/RQcYiN5
2cXvqsbWh/Znna+VLPaXmATF5jeQEbo/RNdDEIr9GULUnP72PLEEBS9HXb8PWN5qg09gDi+OS5Pe
efYCjgXRzCrAiB+L8Luo1M7yL8lKzpEfp20D6db5xerik2xWCi0dpLPGtgHd/p0RMSKPypuNB+Mv
93fAHpVFW3D+d+oGNjjDeH3fhw12qqIaGoCSSm16zu+cLQb7kog1GcB29Am552GBXYHNj0MNwuFL
cixKzERKwSnmi1TXIhJQkVpsPsEMBHAwdYFm4M0LieWwMwljT2YRKwmpa7N4fOhf5BBLsSE27rIe
Nrs48m58vJI6qgNudeEiQGCKr9RXoqstkJ3B+k10xWVFdTnR8X7TDyUICmthMPYtnc3lr+diex83
QojIW3l15/y69bGYcQs8RSRKUWV/TAfGWu2mbU6Ry4az1bP75MITJCkt2J0DjfXK8osrh5R25FQJ
Ms993JxOOaJnIrzw8A1kyk3QrQuV/R1fKAz6b94RCJR+lKaIqiIDEGMClINDa73uWKEjvUCXx8Os
QnPXXTDuDROpQSy/O073/oB81vlW3nbesYRgsbWzRyNH8/5LWq5p9yE+wbdb4B4pV5VTOV7lpctq
luhm5QpG+DNU/B6npHynQu3P/uGRdPfRrBWwiwRe4CTi/EcOrJQzh2ROEsWjGHY+v2j6ODC84nN7
GElpbJwZoka5l0EuZQpKUu1r+vOppSxh5BYPykFIP6ceqsF33b/L0N4NTEFUDKRJGo596vCQ5eU0
gDjakteZqLZqLRXx3DZNlyYa+Ek4+eqG1ml8Xy0xSh+LthGCnYBkQgy/FbFx8KsYl9hMXY6E8ciM
1NfYzLMIBTn6/0r4rNxJqXRilC8q5ZUIk4St7F2ffXAc33ydfsuOpq1qAO/bLlqpyasj7wzuq4Na
RojVOW+qgRWatg2vlbwI4lQH8YkwXPTpOvYNn6Gcve1jcIGEWfx7M7/HzPU0Wn4tzYCnxBtmvM1a
AH1Tm0TIjfnr57WJlMMb2yf6oHp9njPD2XO1+MhY/1Aoxd4EL9MGrWn1KVkj1eKK6dxcvpoSok6G
KQcvvcNNGkaIjPRvakhpH8/sevjiVrhibrK5PVmGsIPJaMd69gUw0rfRyX3nWYxvEMhCguCANgk9
zfrC9nUl+iJnE77ZYQCpNQiU1xP/xy2Ge6Z9sZs7Y5aIsWvjaN2LLOYJDbtk347uWtN4vkg1ToeF
fupPGWjnVayUstSYn/W0m+TVUbBo6SxWM4fIq7zbTl4qBYRM01TlC9+aBdc4mNYx9c95tFD1r0Lw
vJpyUjKXmYnjWzHP6G5gLnsNdcKLRLb+pVbfvUp5mlw0kaYuLviKBzwNERxyCrlxvFJ0H4ZwVRo4
AT1N2bFo1umRbtg26SvACunSWTo0PFg5QpO2FNeHGGPicSpCGN2HY8Bc39a7NNzB9IJ0zhckhSEx
OA0bHm5/6ImuSiDnjjYObwWYEQYT48hqdA1nDGr9YbvcUOre3h5E4XNF051oqjUSsLQJn4jlKe3o
V7lRibkwU8CQu2g41/t9uhFoW6hr8XlSHGXfX7g0/Y82VtPiEn6n6f0PRJjWk3GuKYKlZ9TlW8GT
WUSQTMwMxqHSNLqaAIHVH1jqK27HRzL5w5OfshgJBxg6qvV8JnH7V6RH/JnAluZmoHFoo9dYhfOC
PMg0WGVtDA+ngUwSrG9YDf55AfAH8RdEFMV3x0SlTjcswyn6cr2PvqrVmx9pAGOoDxUZXncpZQqm
e0WD8wIjry2hZWwSwSIAwHrcVrILwnYGmgoBR4tXRwq0PtrmcNJ0OKDsUBk7NUB0dtb/GqP6DTyT
lFTLXou9p0U1jBsvRdXnronySijiVVpD+xXLiLmm9G1h9vOuACIxZn7m+harhl0WCEBaEcam4zEi
VcSCHWJtQp641MIu6kANNXA7I2qLxAkQBuBSNo7Bbh/g2I9fkbJPGkXxfNW4p+2Wua8vGFGeduWQ
ifts8eK5XqiutyViepcWQ7ZxJYhANbAcBzDVMqU+VCCCGY1o3b/53bR0+K9/TAO9qDdmv+P5COSD
jQbwZ42wapSd1bOCLmmTHxYUqKuuN4DoLwsrmHKIgkWgnqIzDTj6Rf6g61sZMcZVz6umhoL+myeL
5x8kc7agGdx8D8Ry38VUfn+oSXd56rZGWj2ytI827aDOKkSLbdGNjg8JHi1T/Z+66d/kjVrZLfy5
8zte0Dok/2GVHUCbpw2OkSU6lQvSXibngw9scnlHxDU0ZBA9khQ/RgiWlkeZxMTGNYywnKHPHrku
RWCbpRRX+yS45na/A2YejOSezoTSuyzsEOJO4i7ygu7hGhptN9p1dlH8kE7HSF76WfY02U0hSica
EetUatqYvXk+lDs4nSeM0MmYQufw8hHBgDWZMlavQwPcaNIs+ZwU8q+0nLTeKpms0wJhOmfKw2bI
Id40lKZMbRm49d1mr96AFvuPANnGOtGjSeWp8HP3F5Ob/hcDH4aDZomicIBfF+PMzZMk1YJK4QSb
QZduojmipgJbKK9KrjD3Q/cCbP2ZdhWQQaG5kA/GlDoKArPMlWOCybltWGFFDt8+HrCxSTWJivos
FPkM+ZOVp2CSY2USG+7YIwgzEiUosvB6cqpATmaQOoWRS/n6wVMrolAqV58zMVEVdXar83yU9eYX
T+FjpWsK9osjBQ+Ue4aFk+nioaEJy/ipG5HMtw3avnkTFlcdY0bVlzUnyrfBJUWmY/F5LD3F1KUP
tMkRzk3otnO1hrvyc2duGA7u+0ZokWfFfd0zh7vJZzIx4cWVMbM29PQDHDmSOXtSKWKD++1imA3b
Qfi7Qbikeivv+WKurdluoS/69VQDQ7LBaFk2KxMsId/S0+ne6fy6JG4cJJ501OdJdateU4ceZfcD
TkUimbsE9H1AEVp/K012702ZxkqydIJcPSAC/AmFMsUvdJvVdG1vEAb4awZddW6l61vSCNiiDqFE
/59Yx3eRpPtk+StI9Olqq9sZAyk+CcYvkQvQGM6iGbbl6kHqlt1CgCkjIAfkeQaeReaknoUTqS8t
ZM6d5TPJG0xwhsEpqJhOkwEkGUKgrl6cVJp4W72RE5Tgcz0GAV5wNgUadcPOi9kPqUEwRqEyZqP6
F90qg8+7dZzGGbkheQc2eZwVM3lTTjFtmA76d4MuC7n5du6ipZVm4Nd8d8IkZK2uV9QczyfNnMxj
4dmPJDUDoeYI3HkROBHlboJvc0ht8MOXiK+iqiDQx+NXRFKiWnvwl25hMlaMEVG6qUBhpMrAObR7
Yb61NFFc/KT0v9aSFhT4OZskczvWFXDLXHTHgjZPQuCl5YfV3L1GhtmmM9rXrYTzSDMaw8kDrL3M
RBMCkntSiZh09CPWb2MSHm7s/ofE/xXxzF/ynPYIA1oUjqpPvYqefbZMP7gqr59iFdrKz7Vnm1Cu
mIueuwnwpl2yip/UTy1reH9IEsAccBYmp5rzAHv6+XNl7EMeyACBMsJbxGIIuUTJYQnlziIeqb1T
xf9f8joje1BwUMoMwg3KhtY6NTojiE0DpCUVtCFqTqgr2vJ8ilNv+HrKrQGH8FWvFssljnvdoMiG
4zfPO7INtM5Jkw8Nh/N1lCINveSmAb+/avrChpXvQfXJFZCHOa4Q5jOUDxkH2ZFgBu1WvQRk2I7K
YVFPPRb3PvKbPD1F5KZBzwkjNMA34hoa9kNkO6/+JiQO5KR3mnC9jjX1dfVMxpfuz7F8vO231ysu
OS7d0dCOj3z5FiDg3s5aZB+3esuJqN2Ctp/2hdDU6fkpk7qEtoREC0CHCzNxuv9Jv+0rhn65dOFy
tbf5SAy30+173ho8bsIOXKIr60cQAz00ixMr1Eb2AQSPPpyG6qa1pRA/sz7VfCgqfjFZbOGOc0oY
SdMZzt6I6IO6iQ9W0M0pP2DkP+lFONs7DVeC5w+22Ys/1mG4NJcdL1qoLhjAoinAEYwN/8vGqM62
QT1xhNlRqxP4c0xjXimdWE8aaN0xgSlcA0byU2G3ogpuuLGlaCSFYwGXADm9uqqGhM+nEpGlqDsw
ZA5tpHUNCXGwPBBLw33Q9Z+qY2PDno0YyQKqpGIVyqXF6nVn7n6jG3wE5Txnn1pYsUXq5fTHfAg3
yJTfd+/DyeHOE5pm7fwZKqJH7FVKtIjjYSo6n8XdMnFrNclwY/tPJdAmIHsuwERVzVIwA9ILQePq
u+Tm8ZRKf6owvOolFGaVgHxK6v9XE9C3Zrkfuc0CVmtBBjcdNY6MZz58HalBNAbDZngEE1Wq1Eqn
ukA7MGEIpKDOdPwBFlMLK34UaV7onU1lMSsvhmX4E9eTRpaaF69h4+3x6X8Plrenpa01GL8W6O5E
4gg+ll+Dav7tdXuL+h3Kpe7TvQICy74EqUKHFkizPNzQLt+uPYossYkKZHf7cGYTIcnB+N105tA8
PPjpm6EPzJwyKSRyoPUYBbmupD3/eta4PmqlWw9fi1Y9P0U6iPR0syCNHeHqYRIUjbj1weGZkxYh
ySwfl+loajhvxJnPqqViUs2s8/D4q7rb5NwHAVZb0GFyLNg6D5T9GDdl6ONs00wWMLTO54P9t49r
ufX4L08yRd/VdQ3xqW4iD85Rt/vBcjQ6i14IT1BRKi0OdNkiER2PQDCFdKZnVz5o0ZnFnulA1LCU
Xi8wUMAtpyVf37l2rSQM0P0rlOB+l2xrfHyPgMsZ83f6j/ESxi7It2cHNRzCY3musNqyD6ycIwAf
m3QgTYqri8y70048B/svCMcPxmOmYwzONtWTfqfqsGMs2oUllTkbGzvkKerETzJm3m35mlT2cl7p
5JWMBD8QRDbuRtZBNYQUsO/7nT97vK42zKTAmsk9FfzplEg2sdkmUnp/ulspgfjdZcl/pxF2vIgS
v3dsMhDXnFCC9QadJktPc9+t5dsCIffkNxIPbbitAY0BG9tDhJo/RtZjcksvIn7qRkfh5GmD+aS1
zFPQIwMR2RINrz9b1TRicW6obcu0igcIeptKKveUQrga3lgzbHgznCa7hqbxrR7OhKT86Ay1cpqv
wYB8Oc9a8tKQhgZ1o6QjDM/CBo+X4rCYwNEw6fkNT4Am1A4hrSrqczOWGd0/mdKng3+B+LAwpEhj
0+Il/MVwS5XKr0SpHMW2ay1/WFVW+12BW2cvdzbZhEiQMpHMY3mEZzNmcITe7Q1TPMvgQ8Cp2znP
FPwQKJug16ip30BB/AAQ+6KZ4E0XvlqFhwMa9olkIynka0Q+oXo/8E0QK1OJB4nUvfUXYVxuO7IS
i4b5ZeXYiK2GHiZCKljQ9XSPi7xkK+6YaHShFAnscH+06IEjelylMHi8zQ1/xqew/CxbPX/GIE6K
xr+pAHZHESNg1y5kUIVq2xW9w7KJkrAKfFLX5gANKrNUGNk+mL47FW+DzO72bbm3TcK5ny/raH+W
KNOtYn20sKWlBJCNo9xykJgO75Jr1wuwP0jactqg9yHYisCmFRSMBF+2O3N9iAx9F/prvlUh8DEM
1b4cv3VGv9+JMD4aQ+yl6M47D1JJiaz6HgV8HJl2EVS+KcRsHE1w6DQPsgF2g7y23CS1kZ3NLRKy
CMmHsdR+tdZWgzYEacCt2LBx9iOEvPcvY32lqsY1u3nvhB4ojLDDLC+RdVvNJj9KGTDz4jklplUF
fFcoj8VGC2np6alwnNWwJhrNo1HDLyHaLutygYNl5xzgxLdkn94CV6uViNne1+cSB+GJzg2S7tw1
1QIUZxrK9Aw4VILJ+fpoAoAqfSMkG8urTSI/Y1Nr4P3B8/J8D++hsBhjmwlTa/mC4gBMf7ROMIP+
D59OxInvM3lDiK+zEXxp8h721iC2ZavOrjOn6Uy0H5xnfDew2OtBQe3jmgGMexyLCZNGshD5ysM4
0uwouSg4KxEhd+80nf4ay1+Zq6ICr0kSX8CBHbCspgyD8GwlO6kDSMgoJffGVIMlgpD+JyJrIgEZ
OX3dAdRW0uiblAL1Qj4pBVMrXahyvXLyWMr52QAtdU175yuqNdVk8qbjiU8SH4gwRSC1vf3ZWBR9
l1VsL1RulezvipKCe8zHwX1eIEPqMLarYXWW6cAUiq/6tzDYTw0gTHjLaQ95gR/e34EydOE7mIFC
QGb7CECr1IlSW1D4a0ImizvmElOaiWNkSp0Jc/5ZUnjNPW17UfQ64Mweo6wiBit5t9GQ/A+2ZVjP
Qhe1uHLJEcwtYy1lc5KO4HmX0oBOGVWHkZXvIAW+BR107YClba8oxmJyoiC4sG3Lh8Fj1iDXzEPg
YLu0bCQcxEIw0v8cNL0BQapzX84qoWN6QyqXwtdtPvap2BV3DKtCFWkHki18odGFW6XPEpvu5uE+
svGFI2WTVB0jYhW0xISEVEa+AZggwV4Pl/GppDsao9PIerFQl+siNvHY1x1CD8saNEOSV8wSinmE
NMIZfZ0+jidvlBFc+ck1XejuFjV2ovdD//xIjnmqZqjhp2e03c0S3DFoUwRyGaUxNGSKVIcrBcVf
Dd1I26+nnkx/SQUrkvfKGGb/0BxY3OUvvZp8+aykHFJY/TvkqNi79VqAUeVUlVrSgmSuw+Tfg223
jaY0rkrF6QjDZgtlxv/xAVNtqTkL+g6KWals/nF4+9ULvQbL/849QoAG7K7uTG64cEr7BSmhLlKi
NjC38RXSCaElKecTeSTNA3il5s+Sfpt9UXY7ICDcg+ts+zCvVgPfsy/vU8nEw0fQfz1CGeiFT2U5
HqFBjJaJCKB9SiW2fheuN5JFBdjFFzJBhG0SxJTx30uyKlBNxjzUW9JdniaX7CTv+pZ5cdgaMQbV
u8wu3XTxotVILNl7FNSe+WPhjtlm7NY5228E4prYRBdLZxCQyQIOQk239PqskN1FYMU+nZ7xQGNi
/xhkwVfAlYm9ByvpOQxVvRC8/X9Ua+u7wPLLUIFEnkxOOd74jj0NDajvUKdvNNjimLOTfeBLtBGT
g673vRn/B1N+VYloyICtpRWyMpjUxCNf2JhJeRwuEtyg7Fk6JWTQn3xFz2hv5vIQauU5n4r3TfEX
Z/z12oXQ1OepLC9DZobE0mo1SSAu/sLmiHeK9NkJWaivlrjAcepmSI/siqyd2LowEy9MXELFfEVi
GD+O+lhKFGXEh69Go3BsuQt1EWs0oTa/583epiVO1d6xBW3Qbn21qm1O/8ugwyUn65qUUXpW5+11
E1/T9HPZ5WoIjZJKRyVs5p5VWtPvCbFa3SEBkoCctYRSpVA+52yJhcSxQ1cSlagMO3l58SoOa6i5
TBUUr2DEKDnrVJ2E1Cnkr/GXTYRGplKMCDOG9+z3MbRyontJDU0Vbj8Nd7MLDapL1kcTowJGE2sv
q0L78sJ8RdNleW+53Okns/Ofiqv3UregvLvcNsfIFDHEk7Sxh94GBviMNLmkdGhZ4bSvLlh0P/kU
1fIDHH7YC9b591xqw+nzbtC51UdE9O/qebnAU96h2Xx4Msqy+URsdgZ+hhqDk+0ukhQ9EH6pd8WJ
JA2PZKJZNmjS/S21yU8aknt4+aXPGNKaFOPMYxXfYbSZf3nWZWXcGQNJiYEjtPVHahAEHGDnoS5x
Osad4UAI6IaNIe5SNZLdMrUItd5HqU/PKt1QdIKum1JdW8xElJ6Lg+Y3SFqSzqOUpq0zrMx9+hj4
tub/sy3/757QZQFg3vEwS/KNPqi5z0hRiFNPWQOibNVcR/oQHtWvLkU9gKDqZ7gjl4HuIGqSNBwk
i/U4SJ4cPssyddoe3RplMmT7fVHKVcniWlKRl6Z609Ug5fuvyZN7xzgYVwM4MHrlD/WVIQCXt+NA
JmfdKKJpaTOidaHrpp/6B8h/xJL+4/fPBkQPqxW9DSDvOEjF/W5l3uvotnhNtorhNk9PAtRNaPIc
OmFU/9zuQIZCYpbIQLPLdPDqbdJHe/pKZB9T9akPOc8aZ5L2pqxqjPdHgAASJoD04sbRb5LL/0s2
Xm9U5oeT7i5yAMW+yoYHQwf63ngDkKDk/IFPbUgUEgU1t5c6fIdirHAhfa5ZoHQNNW0qFs7H4Dhn
IV13NC8epRLqHEJq0VJpPWsgf1wi4N2gmiql7tHsSwq3OR5V/ldi21rkQeqOorD02kDaRdlH37f7
Kgz8r1RT5RNt3LcjmvsPirFxG0PuAn8SAfU7+TrCYwEgjpvsQ4rhJj+STEPsBbRxp+Z+tsDztSw9
ckykMmMBI0BIZfDNCea+fWewhnlSRcfRml6+XjkPTMP5+Hhvo4c6I7q8EJyYn7OSLDeEI/n6CqMt
uqNVlMghiyUs6ewBWxdiyclOowNkb1jcU1envaoCT8qWP0By8Py4dNtTPNudHX4iKkKmHPFUPOnB
gdblBWHKyBgpIa0Uhvfy1XeVW6PZT1WcX2EG+3mKKVIggt+olqJrl7OOosuS1iub53yBE/OijGWT
d8pW3rcS7DE4hptZWQdNuPDBqSpn+BVxHyvAiRMlY1oy2J6EacSISka3mkCG9MKaBXAqi6r2CtCP
n87nWJXrJRRq+mgl08qCYHLOVEqQQ1fLwD+5zGMMTCIGoMgjsP8nkSh7m5NKQDgrDg+ZF4EGifpy
lA4etbHVhComUolLLIfoEhy2kyMaggz3UzZsbF46mvSiV8ZM6hB1uUDZTkMfZgho6xuDwDGpOfAi
iFRoCyKx5vAFguufG5io5aJbqOEsd1JeyezYpmH4eaWBTDWeAm5q5st3PL2NunqOlpqzuRm7XoxY
p85ThK4unhbVxYPQfcx1cVWp9HT9ldT5sfSbXHbO65yK6TJk8wEdJrMbuYaef0Sh2dvwCkJqGBlS
qQdUMahxDa+C/tim4OoCHOLV0HzuI7v6U5FH5UtP20yWUlsM6JOHYL0AF3fzaRxa0a4cDr9UIW4c
DWJROLfT1LQbx3LMSqflBjcyFY3VGPttGOtQU47jK6EEpbJm/ffr3zfFEFodnZeBNP1bqW3FvcGe
XW7NzSVCYDF6ie2fPyufIorFrImCTIiH8yx1UEN0WDWcZi3M6XBv3RvijpZu9xP6QDttsjJAyBF/
b806SqmSmCzrla8QZ9Nqm9QT4BHNVeoGrviCMJ1raN0JUB3MKGsTHlAksOBYql2tdY0mogH6r1NX
0Fw+mJglfgJXfoe/WkKFhCE+NTH2Fp6IAhbDynMucKo3z3E0FALwoEMZodmXBI2UdDAvN78Kvf3y
0aobGcm8GDSd1mF0d0k9j+IRxWLQf3p7H484vJ/qKItjfpu2pFizVLleXJv7RLQXvZ0R1J/kobLV
Y0DZKhkwX4RgE1eRnnJKwuHiXhL3q8t1H3i+w61t8p4GtrEAMCSKGMajxJyOtsUpZk0xAP8an3vK
7ghfxZgmLPwrLPNhX2xXYmJVd4EKWuMgZrUOStco/0QZrGM1wn21WdW4N+9tGY2kIGBfnolQcY7Q
r+uQJgylxiK1uTbWo+SJtc6FOg1hfcNsLZCCjxzd+7ZSEIwXPLrQ+Qvq3WYgm5p+d+zZ5hg76GJF
A34dYHkpeNmLm78hs3BATjlzEEZx8265rMnOH+yasawmeN1rmQBzjsCdWi5afKc+62+6mtLA2K2X
7w//WCiv5BbKpU5QJFacaU9BGuaEQpPw3RFh/WilB7xs/XBb5bPxiQ6LutCgcMBdqOM/j62QuqZF
H82Cj+kIRQnNY5SMnrLV43/cgTlfkNWTTh5OUe4L8JhYUYodSTu3eLoM4kjmRFFhKy9USAGONd/Y
zm2prQI/FHOLW4fr5n2AdZF60uPueW3+8Y9zWod6J9HlApuhHVxHp1gWSK2vxwcFq7uF7gTO0R/b
lBb/Av7cHZEsKjtHn3tNcXgGpgeTVDKMIzpj1vSBanMUhbe5sIskoYHI7VHeP39HLtQ/jr9+5Lg5
hJo3dNk/g0kknjXrgMr0QctFR8/5UCycOSeYwY7VivCLAmyira81WkUQrzUYRkDCbYEuRtWlAczr
B1aUjyEvShrHNE+gc/CoEX2qjHZ2mLvmNR6DJBwAgYNIhAZp3QZStt6qU8Vm2BFAeJ9NH1o19qyL
Fnuivtt3r1L43ZuACoNnShdJyTgs3wpBm4eZjg/HhyTng34zvB7DUcx162lP8xRqKWdT6noFKdmr
yuxId5VjXTxaLUnI8I6WLoyRMCzvjOJv/GlSBS5Da16WxTVNf/fE8naEinH/3e0yUG2P+ZRk3kIx
OP6owTNsl9wmdFoE5qFX7vwM/ovvI8Wa4kQW03LWZnq82p7YDf8N8W6TIhmKSKA15BQsjNlD06Hf
3o+ZcQea34+epXzzYb4sGK/8/sUv5yaslosU5zruAC9mWjE3JVauq1kc1AoU+Sf41OSq3Ug58RAK
LuZqRp61M9Q0EcpjDf0LeYO330DqICxm1K1VDLj8zbhlDqXuIxbKc/z0EcpLF92VR/GPUCvc+uXm
eWlf7HCzWpUqVMThOJNHUUdZ+x5rtLanm9eyYfXI45x3NrQNqr2Tby6CZF/lNDOFOUbq5ONG5HfD
IcvgKIVZh9H4w9g3G/1SlXUzzL57uN1qWW1mmfFiHeXODouyd7GaT5kEI7G7p2Dpo7WeFmFtLsLe
T2SvnEzH6vRyYTKJWvf6JYWhH8kM9plxeNokeMA4nPrdpU1MXDIv4BIb5cea+uJ58yDEnaDrd5Tg
FQGcxh/E0d7C71j4YD+bxb77/v+R8lAOdJqBXytBmzaS5p3Be6tvWwvFydPJjgI24Xy8cUHRE+OZ
KrZ/VbiQMDE0iWfvvYhUI2ruOiKIfYdrFwrgULB8lBmpE5oEYf7bIJyRqEbPj5aW79YYWdWH1zrF
4OuW+zDL/ywtdbXpHIoMbigFzfvzSLYuYwxJrcA8GznECQoT9uh3OD7hrAi62wJdSjW4J9LDf/E2
/o7tQo3K8/nO2KnPPkF9W0ikcF+ItUjuxa3BCS9bOWWNVanYufNSixGquT2+5bfjNhYtcTM0U/E8
nF1EW7qG54EXrGZ/X+TmD97UdNOGrBTgXBPfCAO24lRzdT5xV83ddETFRCCBE9Vtqv5j4G+NOkNu
bYwhWeeGQIjxHuP3zGI9IAjmNhCCXIgo0HXZ5hIEVUe33A5UDCmoR5OoMCdeTb0G17WPpZHvAuaj
86/bdALdtE3ZW+efzxz4iLKiHWrKPdDN9WFPl2RFQkm5ex6LesknqmKY1E1hG6YY0Wwpxgj0xJrl
CwbRDqU5sVFG3Xg4pRHOe1koiQofXlnNjWtbmdyRsZEBVQb3DFrgduxEt551WgBLA6Asha8a9ezG
+UqBQSvC2UNQ/i3mS8MfkuIZ9Ikil/bMaCsdrrWFiWGkNExzYOL2mxLSRxinHvb3zv9/ybPQnxBg
eJC9obsAUP65cXJVADneHSU0QlSthQQnwVp1PNpD4xkVbzo3PmTWMTDAC837r9j+EoywbSWKDKrl
P3GlhIyAFeM7BP5M8c+tArRlLG7YUGQh38Yq2qLJqyofVzyuvzR+ijI0BOeIyVRySD1AfQ8PlzwC
uL5da9h8KD1anRNSyPSbPPkkhVgLdBU4MXMZb1nE4aGxytVJi6b35b1aCbHC4JRWWzlu8ZZuQgmc
NpgQ/NQHMBjDIE7hQy/FYvILq9wu+S7H3714ruAZH2Wy/s1G/eBHIKWD2N75/MDmmpys+FIThxtp
hX3T4ZNWUD94kKg3InZJXraMBgk+3Og/neW7GgW30ddnjrSF+XvdH2LB39P6wF+wFV77An3R8Ljv
rHZ/MZ5zPAGGkNXRBKAKwNA1jdPJOpWUoXI5TtcMIROE4/rKoytKRrgHq9RbJYnfATzBU4Ze8y0N
cwRywH6ka/MsmWXKYbmMXRHOdXHokewVx9R3A4uJHY5pUdLs6vXIR9Hi6Tpc2dmro19gVASEglDe
RGlpqjJAFLGvuFSU/aOkDgIiukvF1ktFhE8Wp2Um2z0U4JuuXZ96MArVmV1r6/8sq57X22Ye69ZW
EfhYGo6A2xTkDzLIiZeyhY6vChtF9nXSIVms4XIgmNRetKdXnjGAeUh9T2J0/mB+kELxBsokGOvG
ZbiSEPiXOLQ2d9BjT/dgsxNNWP/oMYs3UYNifwpSKKHcPnXGQkDxPdEUPo0ZaxS7ckoHcQ42xvCu
WfQemg4oPiRbynLL2HnVSwalezd2zyoRXSBK/QdwbTYWQ2LlGuAvaQoZbBAxKeXwujPa7PNkEhr+
rKkMZxxBx3fENo6HQikzyDUSeh7rAIPtkid47a3KYqLgA3wlIQdOpLI/evt858EcU8SKIsnRAt5y
EM/b+/3vkYHTclkBTeZ3LwC8gMuS6baUQ+talKb5dHwi03jXWjK6Sv8eaKf2aQu7y2a0FNphmKke
qM2m8AMQkW1LE3x+DBCxfhCgpb4XzkOq9LQim6MCfIlmnpt/tFa03viBgXPM9NAg/GxqaxJlDDlq
uJH8JLAok3pRWK8/V8LB12ZAe7Sh7HikmiHEuRqFExkebfXCqqZ+h6yDGac4q1UWXMNQaLCqCYlH
UmNJ6elk7jWAOyNZAWJVqeT6MhsFJGGrrm4rrtEw2gY4hnYn5yPnNnYd7bpAY8Q+9OVR/4GcCIvL
4dsCe/MDH/b5LmsYnEMTB9N/zZ7khoLW6xtzSnbX7fctVfb3TIrOiCTHglbRwGw/HRl/FSk/WArw
F78A6qY1jWNxVGLj2/hrlxvkbJ8y+4X+vohg69esc9+JwgufnvuC+86PQBYubK5g2y3IxA2qChjO
Y8rH6iYxDl/X3pSkfY4egwPnOCIeLcdhaclgzjRq/GnNwLk54SnLhTgxyBN5UbWOJoncsqxWrAoJ
ognBFYX6Z+gOJng/JToNp+TZuILaR+WFC5Wko+fy6o2X6finvWN+/+16/9kfSp9r85cC3wRWtpaB
XFF4b2FlWl0p9qx6OnEKhjDFaDi6NFOKyFY7rUefrKjvua76OmqUCwsaqgrsdHqbSlMwZOmJ8eur
g0n3ePxdkMrNOi2H58/MgBUynEaA5uFnilojN2z3IoN8aoDqPQV2Xj3AGQTW9nBQ42yW4b4zuDis
UnafGvXQEvQR4Ct8XQEujpYOOrodxQwUuqxSt27LpYl90IVkQvl0j95lNdMOGE/0m5npmZrIpovv
RI/UmV4RyeP/G5WA/Qz+MAcAuhvzuJ6eyM7sh155RDn6lgHZv3bAqptUxLoCdgqWPSRKYsfwgQlb
U45Ye1W2WpRSmGZXcKvArK68+hDYRYZNBgdhhWddOocrnhaZBLwiDhwdsffP0S5xSvM3E8zkL1cb
pEt2LSwuI8W9m5RxPjYBu8XkXkUSwvTt9KpjzxNYJGewZCups8FPsqpV4OlcIOqtNSYRlCgDohxN
Ahlza9C2rZnjhqPu95XUgcrF63uhkvR6vaFGsPCvFdx4koERUqvAwYUldjtK4VXGirNShCz/TOQv
ZFBp9ZKToihThGPNC+0KOh03szyd2vOxwmU6WCuTOpdPcQukBn74/dyQ6/33OTUBDRxy4ANtoSV5
7ObD3zo7YjEpFmKPqLhy+1KUof92qIQrhK2K5htSnE0+MokUWYHa2NAnMB9I0FdS4aDf4E46L1Ms
OOp5Vndhloege+FZAr4L2YfXKOXA5AR6/EKCA5agdFpsXNdbaMLiQufulwbGBVqTk4JAK7W33TT9
1hsbC34/nLzKjSfzwpz6Gn8zJ4nl+DVAy5JM+T4KCD7e1jqMDGgYDCnJCvzX7c5QZG/wBx9ycDsH
vfrvHdBJgG0h5VIfuCsCV60Q7AcMUZT1d3GvpjkiUBvm3iJWYGfFaMWAHilOSNeku5UWXYEEMN2n
SX7JEbTdiCu0VTv+NJGpzOiRI9vVrk1X+yCMcOQ/Um3Ae8iQ7EQodkbmFckdYWDYXPE3RnxF5Sc5
cB2XnudIQvSS0Gq2r+CoAQkQwYKN+NnpESOEPwSkGUuEGR4+n3aC22Q+75SE+FuF6KtKkgi8IAko
6o1C5WijBKGzZsLWXdb9sPbSAwJhid/D2odO8PAiqt/FD87d6nEuouf2LGwyphYHYPvg3ohH/EhB
HyW71hR2NICy3ivyXePUftA4UHTwjmHpo26ic4DriE6d3f6GpLjOyIKvEL5I4GqyvP70IEg3YQcE
UA//gH7/Q25xOKWPwjbjqEFBIQOlMyMI6EeRA5t2de47P1nXm9SP5rucjjZrwMe8Ftrj7AHBa/VR
fXM8kKZQUZJ4X/y/MmUuZ9DsS6VUgJX+9R/BonqTEDyWuGJYjx8A2LPAa+pJRk6pGhQTlQ8sR0dm
9T2jb059jfQaLDufpoVOuDKqK4429DB/wv8pE2QfjNnpftqP9u6C2vOqIa6BuV6twXwYMMddDfLH
VXWpSxKRCB+XfhBLbg3XMkeP15hkh/kcbnVvR+445W6lyOtKk1Hn7yBC5sdoISPJ4RyJGAlwK9QC
fd0WEb7h6ZmzAqCFybwHQDLIozC4U+66VdFBB86vrflZyRqRM+i5gY9uy+b8MLO3YfrlEDdCLNAq
zRjsnkDjQ/ArX7WeIQA9P9a4LIt3w3K5TFpq6/Dr8SvVUSBeZS6qRCkgwWDRBZk6RCUqJnSDqtBZ
ZljK/kjF0L/CFrdqeEW8s4dWgrkn1eYLoohBGgxPQ+WIRQmZDMzW/zanmiiOZeCqMBMMbRHztCqv
+5PtuEPOIweI86HSialVo+l0S1wfCaPs/urI6EUGcmirVqBLvQmgHwRomA69NuRRp3hPJDwPgQlI
3wnh5yMGhR4kqQBbfvIeYsOYpqQDvY5iMAYe2Mu9V0hW/YOviAOyfBM0M3YWbXwe/fPKm0WI+w8Z
UXWs19IK4UokUlWKj3nlGgVo5qFIF4v6HfcTkkxkY7MGv/i0L8k9uZv4x0wVTrQpy3hiWbdssFyq
x76CYPsAiAazlDENJ9jG+9cJgXcB7KzNOn9VFKBig2rQrJ86xNG3a5B/dBMkXzugIn4pMga7HDGU
KC7BoID1fedRw0ISE95AIFgETttKNAzeAg00X5RHFyAwaqI13AtgcLRXGq9lqyrHvL7skvG9HpfL
yTftm4/i2OM/OhIVl1MMyf0DItqlKAdQVqdR5kglJt7UDuHrXA/NM6ITRkSonIqsWrmT31L53uDy
x9uDXHfJv814pWc4WYf/F3JOU4sssyQ7Xx1LfabG5QLvwjVurzPI+y62dySrr7VplUbX/FrfqIy2
ugOMPQ6suDeJxvScYAZ032z2knvj8jzJbmhx4EmfgH2LYQGRucTxLPmAtMkjyBAuavmoFyNJOsiZ
U7SaER4MDYO4wfugtXjLAuBKa5CRgsDmOHj3Xlo/yEK3iWc8YcIyONErbhlNLqXsR6erUMV+xmX+
QucTf/hab8+2hlQZ3rglZnmLaZt2FPKp08SVv38BWepI7mNen4xTUovoVI0apo70XUjcHvv+2aWV
2ODiok2FOVQNQdg4EOsY5AUizrx8xRZMkwmz6aeU3FoIZpImQ5tt0DYakDoj+zk/dMYs4/aB4Axq
Je0iAsY05LonGtYuNWdjIt5iDt06JzqksZ7D/1MW8C6iP3l7P1H4gR2SX3Jlh73DOl1NKB+mp8Oe
ij6jRJpwtQzy0FAoxgGQv6hJEmeq6B5KMHPPlKHCoh+gwA+lJqZffOmRk+/Kda/Q/tjyHJo0bV/m
yDYByS7vP35Cxm9qw0RGLVym4MsqUXU8CieX35SXp+yV2QkGCUwNCpnn5BBdxzkO/VboQICy7IV7
ow9ocAFm55oX8831zlAH8X7Z55/6zdZGgXLESkpbYPzO3Il/MhcFa1mPz5s9qp0NwggrPhgImc+i
vKNhg85N9R2xZEG0RiegFQCd98nsQPiVSfDUpzUeXna23OlO4V6cnKBhtkLzAYzrPTIaY5LEL49Q
OaizvlDAHcyAbqqV98W5VR45JxZXicKzBafKERfCbuuoJYgrG31LMRCJ40beFCVIAoEUpbxH6CKx
yEjnfU/iczXvAIcSk/bnFfXX/xWe9bP7qLREQB6dKCL9ZTapHNGto2THbjejXzQOKvlvXgCd6E2w
AbxR+7Cfe9H4J2D0vjh6n6hgmEkwnTvOq+lWB0CPn+HGGlqujV/U0coOP6d4SMpdihHDNDdl+Yxg
sXXvF6bLKHCfyoQ7NWagkj6X1mAX/M8I1rPp6IBCQPOl1wzax2Ig2dvKLhsI3h4rg1nmjE8UTB89
uU5ejbrbrkCH70egKLY6A2L5Xsgg4zlAgd72/mMpR0i7VlwHeQ/EYIRr8x1ievJBmd0JBCk8SklV
SLAK/NJhB/9dSu2Mlp+KQT2EFTt+xQovfxvYeQI/WN8zNS3DVtazPtTh6+fYLaOaffQU9qaXIxIe
SfX9lComs8bIH9NsE/SiPF83APNjGxUjIk/qo3xUOv+BBmkAYa0QIf9KcmwvtXez9lIYWJkfjPvE
ax3IsfmlU/89HKzS7kDfYi/LbAmnDb0YMVzR6CEea7r0LYN/gZdHci2qMY9rQoq6cjJ3geuSpR27
/VIBUA+GRyAYz/+MIDiprlrSrQU8tKLENwk6cgRx6A0F5jXyLAR233zhiGJYRLsl8wpiLRpEIS5+
0Rr5zLDjHdZifoabQzZRF65PEjiLLYCaPJxEABpqHjqwH2um6jKgERioa1foQ0FYDhNa5s9wt+ra
rFK0YV4Y1+6UhuJ1ftkIu8g/50W/o2eXfPJu/a2HpN7mAj52SMJ1dmQhFMih6DIpPLadA4t0c4JL
A7Pq9MaixxA4opvDwE+RcibXbMJWcbiDgbqfRc6z89LPvZlOw+t9/d7o9sdM60egE1rcYG8H3Vy9
R71njh4ThsKyiTTq31BhwWq3w3jMgJMT57iHwKhFNfMROeiHvVQC9l0Iiz0XOiyy1e/VM5Hx/Ity
quBIPNhx1sSTEXDv6NK/0B9ewN/udRW9xpqEDuvE2y656IJbnAyc2iAowZzSDnPh9xGHCPhcjiYV
Nwo6psaGfcg0UIx0stjzidZkC+fWMCx1lEaz/AV6uslpHcBGNbBsNUPEzJettUMgcc0C0vvrhMnG
YIaag/UH+o/3UhFRF5iov37AOmAp8nUfxoVE2tq/HmWI9k6TPMvO7+SR8uzNe0d8D3O9KjYLJ6D/
pbb8cf6sFBFq1S1uahNoWCt9rU5+0veUdp9JN5z1LE0gH5Que1z3cVkuxQjn14SiTWUvvU/cr8g3
1JaTwQi117zsFlm8aDLovnJBqWJ4IJewwdZ9c7OCdSGi61FYxfM6Z2+0YaiErkfcAxdO/m4AI6i4
Sf4r8h5ov1VTjWRhX/elnPjuXpYti5C9zEGqX7TuhzeSUkK6PkTsn8PzwDAav8AUYJ5rSJsKActW
Vh7/Mcg3Oqyvy/jQl2u2PRWJ8x3pqwHGsH37yXfuE5f6sWTqF6FS1b+IcILsImn8lSBF8XVZCIO4
wa8xi54b1v6vx5cnCBoTA7ytxfImts9myZkCDg6LfhPBxQKIud+FVDHZKHWXVEC6d8PxBKEgub4L
yPo9mXYZIVhON1n2eXNvzti9aiUK1IKvQ+nSNDDQVorVzHQ0rOEcl+4dnOyTOjGZuNWqykzI1GRb
DY/6IKA0IY0SMS618SyrBBYPSVVumSryLz3ba3XWB1hfAskuHHMdxDDsx7Rsv2Ydx6KOAIe+lido
qm//QZnZ2SOPLIDpfjV9Gsv65QEfDHbjJdROQsKjAiCVVoMzoDuWu02kj24ZOSSm2v/+iV5IKaa3
Rwg9MqHgH7exT8FFmjVHxKDJnQe+zC1YU4BL2v6XldrpCuhxK4TDctwKnlY729I1HVOZLUg40YaX
zvAPpM2bwSEgXwshOlZUc7cycN+P0yUCivkntQxIawCtPOfdAnjMrcC5VGQ7SEeXRN1xVkPFJO8q
b1eWgerac/5myZa4QijNnunND9x1Dlc+/4kgyYpRk7itntNFwNwh+vFOMy4qbclYiTr0/MMRpnZz
/EpQqMfk+C8CtWVyuSblRG+gkV0EkCtQpSVcraoxfXFo/+tPwwBAzmDv07pVKbbnjABXw1pATYr/
o5MaaUMlDwbW4oD9SVNKDsc0q3o6QbTQjogFz1digX+FtZs5EWALmaIrcK5eVOanJ3+vusjEXrj/
FRsqXKlGGHZE/05iGURxdOTJdqPYACvOfYJ5N5HnWICNJ+Kr2IVNTF4cpKGoRErkGP0cPpV0TnBf
N6ya36pKwwzQlgThJFTPNFQbb/WnF4ZgNt03PoZCewRSxAKWrGc3x/imRl1W+E239n5bJvUHsDge
rdpnM2IPXUv8/BzErThw/W8ZMNS34FOqb9j9iozQY9/o6WI8i76Be46b1NrWkc8UCFSaAtIIEZng
9O+jJCQc5uu89ZuCl3cydav43OOp7xRzcVNeF+19YVMPhUvTxANPmKgDN5Qz3ntKcXyrcHDCcyKJ
5yxYXak6bIFtsm7A+aqXSef6MQ5d3s5APrM+jajuT3TNlrXCAu56yKErGFGkKvfrRI6G38vhjVaD
cSPAPF7dvjhChJI77k3Kwy3wwMySE4INEdhizBVLU/IyBL0LHrI/zTjqiiGr6A7ey8/QwufnPshh
rSVd/s5Nm3oFBxyRmxOw63yx8HD4n1UopFIu7nFP7FRbzj0poMmzykCb2FfaNhX3b+hTliHaQ/8o
PbyrTHGm2LMiEc1A7RTpigSsR+zL/MHqWKLIPNvMfhvNHppkyQxLJEnoGZvGWEloLgUlzNLnQUKv
57edZ7O5tVCyzZV2M2TIRo+axQ0YMnalupFPljFUpOIwxUwhtq7Y03cGm3KDON3v56rvivXddA29
1BLxMOgsmPtflgA/W/3RIFZh9ey6yi7Joaw9bg5jBnNnk9wZeJdIwi0ZwutiZPVM8V3PT33zS9KY
J9V8RwQdmz8s11BaWd9ZCAvFUuOOPovY4YfQcswttYY5a1SoVMk1M+tapFhDxJ+P90eewSwHQTKG
rtl1M+2TliOYYZAewliZzr2pxXS619co8Z5U+Dtv1/Qj/uA5Etlu2hf8KLB644u3oDPcdsGPHtb+
1ZIjgQABR17sh5U/JzOprfzAkat/RRa1BWo7TuMxX54f2y/DpW+EWGmSYAkNdspAy15ItRllW1rI
qvFBr6SNcptrVLZEyCoWdt6gTDKve9fOCwVeW8sztlzP3X3u7sZuQJs1m+LQPz+H5NOUOpEm8HSN
66NlWX0evkOiyM0YxHHFeMoqecBjATZo8jQaKxYTn8COBA0hNaI4hD66onAg0VKw1DXj8l/43fCS
2Ns+MVRQDIHvUWlVdwpU7mjOgS4sOxdu3bmoqlSFnRehyCrAWtiDUKVs/4Q/7xgA/ji36jCYNWap
naiV5K6+D6P2ezGENh75jmlji0wStgVvxmX8/Kdtyw7fHXlyha1s4UWn8PweLRO+VNk19SGPWC7Z
7/75nCm8FAmvyZkwxCmZ46GG/qsEGiFGZP+QXorMtWIPY8dKx0BuTVOBdEBKSsRZP6guw6VKg/cY
iSOfE8q05xQvEOoQDxNAI2MsfnZZedZhbBzJz2Oa5dOIUYfJG0omfrLO2tIzDIxyQfGi4An/7cKD
42wVvvcSZMnuEfHx3L5daALSxRgV/s//O6aCVpAth2ZbNrviylQBSGRUhVW2Ky1T438htCi5HaPu
CxztkLH09P1Arf0/pRQ1/S5e0vU39ootFBolsQDDwSXIIJwcoqPaaHCbMjao6AaPJFYc/NCXCuzT
84HewKsi+QR3OD1t/dLSFqsZvnhnrnCBgCtCLL/r1MAnPKKAL5xYMNJRznpWQ81n8qiHtMEUMYOv
2FKzZj8aEhReGPfFkgEZ/pkJAjq4mwky0oMvnDyXTedmmsPxKj41R6OO5ov/yGVuRHDiFdz2KtgJ
18a4K5J12zsViiuQ1+5q6t96n2i0BZCmvM1qvKVJNHwGOXByWN1Qu99WhTFEytSdYFm62x/aYmCF
ZfpkhZHYHmpuuLkXVSosKyQozCKFF0ZDstctP6PybHUbq3S/29G2SKW1kQEbW5+TZ5JFuh9JZryn
BCyp78Z4qtKUWfF0vUNZKwwmtdn6OsqHMhy7Tlgr+slViezM/as/RXhjLdQimunn/D6TAg+5tXVx
3lTvgbtCunjZzFJABiowh26A9Mmgln3VqJacw8VGEA9/s3LQxzaly8Lt1eeYPBBmm3PR1x2VuQuT
yP+yEFIuIKxiCts+P3GXrK/SE8nhNcOWWdT3QSsZKS82Lxc7+2v9aw6jQZQvmjwLc/IJGBNfFQPA
wbEaUrPmPC6pxYRCFTn2VftDUoSgJawAHCrcW98EGcH1KlX0Q611IghJJirS4o9rNhbYuOAMtkBL
2YnnpDJaBPqgPJ5o2IgQe0KbdDRk1nOQllIw6HZ8Fd1o/Nq4LTlAU++5e/WiVbQLfErSHalgrfcE
2i2cdgkBY6CNW/aAQiaOhQTAnULBwRUrMMfb8YPQaKbVK59AXUSXRj8Y7+fVHK6cXwkeRTjp6131
ydvLeklEAKTMAVI/INJ3MJyNUZQcgtR1am2EcJJpImWlPpkxeZlpBz3REFlGMtCzyNwys5wGwFjr
syjuki1iIYHnGEnbMXS6VfMCWiunvHElnF5JA2FyD3yHXC3lrkHc45EImXnGqjS9nsUNJxyT7o7D
KVeS5ejzEbtpQ3ChIIND5fY0BAs7QRYm5YJ66Halp3JDtrmhOmCUSmRKhWHd6Lf8rRYV5U640wQ9
bWxVGb7x89WiCMsjISGLr9ZLjs30Zp/U0jsckVAPy3YZoj1TplhVrcAW+OAMee/0OK+wrjeW2POx
3V3WDaGu//56968x1pgrW77HgGGCKVvIvwBU4fzNjeekCwp6rUp8/ADYred6Ug+/iNj8+d2Wat9l
Ba8x2QXTk490S2ruEtD5MJba6rGtnL3Ca/gH6rDHESxc3wYYsDLSWd+mmlqeQlCSSoG0A/700bGB
+aQ/IswsMmjNl3OA+qzGZ2O3EslKw/00n9/2PE6tR/ygZpRtHIIJV08EAKdYIFX5cp7xCVoa3U55
P/mylUeXJOxFUURRWdD4BoFGQrcq247u6YF6d1SCNMBtAWajj/n3mV1sjvsgQ0tXKVM3an+tF6C+
YW7B0TcuxrWTHhkn9qQkLVywEVqiESErubySyaF2tfxMSeV1vgM6xpLNI1X+I9WYTLh3ocvkFmlp
lD1yPMsiVxh114hJjAOSQrgPsysuPBgbmLioJSH9bmsA9ZDGiIzJt3rJJz8mIWadiiKGvyn5XjwB
/vHnOS7L3wTbH6yY+eqOX81l+iHIo3bChETVKC97Y64onONmchdqygocs+5ZMv5h9LDAYrHWthhe
RHA4+way+3O0ZVbvbg2J80Wpp9/5KaPUnUjCMs/eR34oPDLscW81aTlQ0VC5dEQdMykA1q/QOaLP
6zjIdehT887nXgu1q7ms1e3ZJcDUJb2VfbbMFXQlt326ABHRtOOzZYJ9jqb7qG1r77DOAAisprP+
oROuU7qQL29Xa6cc3NC3vaZWkCgdjGUcKpXU5wJ1+6icrgFCBkG9X0XDQw29ThEY8TCW+rRfqj1q
SwoIhUzzjjnC6LpsemWP+hpXb0SeWa0HlR6c9mYg0k2niQ73EYYWjOkt2QE77/mKG+Ubb+iKJKve
90/dtun2XCB9g2twrDTS36r51rtzPoXq6E6Sx5eUUMSDV0SwiKyFnHtmcWSwfG/ClKBhp8C7YP3h
4iExfdcXPcMo6R/spUX2szWTACk8IsojtpjLRpkKuK8NTxi5bJDbN2DPl4GgoA2N/xPmAb6+b9ff
gxSb4+F8Xk8KyBv/L4ZrDXTtphdeV3gDnOYJEAQs3+dGFwgoodgPGKlFh3SAY+fDh8k90POir5BN
Pi2tv/9Lt91i7Y2zboQ5B6NuGr7D3tz6Beubfy4oxwfZrb4ld7EjlmGu/O0S6sA45aJGGPkdAUzc
PN0F49mY/VIt8BxFYaMed9pnmxzAop9bRQK4R0KLsz0edHB82I78cBfYhZoX9VV5DWGwKvA436YH
rnx3gD4axS/SY1mJuQWD1o09JGTy73Xr20Ld1KQL/2cVOe33BPX2OmTb1Uru3mzDx8+qaiEUyZWS
4wXLvHYAiAcY6rH7YBwZqqZw0ork378CVC5YAj5TqipBomca0r8mlDyIVnk/fZnZjEduk7HT2tbc
RhLYKMLfOFCV7V/m3MWcjhp1e++3jJ8DGaJoVO/C9JepLZMNiGbTR86u0d1hqOExHNQjWwyKvZJ0
CeKrrWdf/yHm9BqyAYiVXhb3O6tJuw4d6Trf5xHOPYVJkHag6Fz8ey8H4OjguGwhLUuZIQcFJirn
ezT5aKCYm98tu24jwCqdIOTyVNFqlGHA0+UwEgSDckXgE99GVKeUNYt1X9TMPRnZU4ef215FTKJh
yvxY3kt3rL/wwe8XFiFqmWO0CGhbKNdVBEmULBN1saz9H6MOI0anGK3MKI9jlQJqz6XX3BXRKSfB
cd6uK2cQI1xSzRQ1dZ/UyTLIMBLdY55C/UO4oj2yoJk2FI2qfvwq6ux35fxceNs/7+ZJj9iNN5Gt
jkF8ExO5/qr5lp90ZlkkDZ+PRnnyawNBNKWhCL7rbZScoLRLWZ1Yov0n2bv2oOuHBp5O5cEUIzn6
SVGQUmivMOXw9fK+jLeBpAMl1yMEgk09lxTvVtZuAHKDqdM1gu06Q4TCH4s05/tWfs1oXJcWCZy9
woIEgFCVxxGDng2pVFA0QH5n1ZpsM6vAZwLtOTGjYFs7qTlNDTfTXGAFgO1EDjWhHSdwWZdUMg3D
pUf3OldYKOVo8XbtVQ3mpStSZKVANjj9swjb22gLU5pxhjx8rvYC7vvtw1dtb0oYL4p31KE/nObA
Xu8MdYKpz2OGV2u/uNoe34F69taZio9Ai5joazTtAXO11ZHDbtiKKOcn9tqOMzHklsP31ZqWXGzI
B9H3+HusFmtr0OoPu2deIZnMTH7Bx6nEQiKyEwpfT0hLl3keQUj++V66gW3ibCqA4W1c7ks+UArZ
y620yaH5unZfYq5DZzPYe1YG9HWlv0LEyyKi+I6W8VDkXR05uJF5lT9KWd3wNus3m/8jub741z9s
l3DLBKSS9x6wxKGhT3u7nj/QilT7/80wfctf7ZF0+nFUenou0DVfJ+RN+vHb1B5blevOrk0oEDyb
cnRe9KEKMXzdOzWsgEwBw70g+5ks8/uMFVUvukLPa0WJ0GvNTKkkXzaG2QJUmQwuGxrC0stzI6LB
ad7hTG8eJPyqaGijg/uNrZDnyW7KfCzkBN27mpa4LUtyZgg0Apv/CYmtjZRQ8cM5Hqc+F4Gy0NCv
DLZSU6kbDgiOBJzWBV+0NtfJ2BsLHeCfXTya5IsWjQT+qCSa4ejMJJjwz+6TvheBCaVuiiy/nxxZ
5jP8/uxNnlfVkg00SrNS52rM6aTTi5a9fXNr6N1/7aeZMISlnYwQtvaIoWFEG5R+CUe/K90novE+
PEoZnRBmGWbddiGRvLp0W7up2iel9IkEnc2kivIvjIo6rHiz6GG9PD7tn5fMXkm5SNRifeHmCVU0
R8uC6SB5lp/ZLKP55CSW8jKdr87R3EBLMgjDcqk9e98HE9MBKVWpRpFYQJF9p5Q6GmxukYOyslYf
PoZFbHj47M0c+vweLCHi68Cg93Jrf6VKs/nxYOfDbG82yntmh5PHji6n+4ZqdaBa7K3uw5JGR/7s
V/XacCpeWeuXP9MSGCrdph+c/Sd1m+UsuyAbztFrsER4SG6+hYGwLxvxavlovfsAFyerlIgLu5be
k26Wg3ZRS7U50o8nY8fjaw3gu1hstXpHTISIG4dryEfsATWM6VszvNw3+UGqQdHq6j54fAnqGo5a
j3haYQyBWvgqzwm0aeZ/USqW1jZJNKk7MLsb9WehPadYVhlxxFn6gDiBwfu3Sqdi2oBgyv6Q5XeL
TcYTvLozAIVW+CupWvfGmg+7QZLj9SCM49YJvLAVbifbeYBpjaa8OFHejLC6U3H4xpY37N1UCnJq
yG+/qsnYuC5HAsrcP401MsCReaR1z+OzmB6zHJaRZ5i+ShKFnE80MyX/DT9MbJRJiy9S3sU7qigJ
rsDN8DVadhvNNTj9xI0hNtR/h5jVS+9fD16SsKJhJ7rWEi3rhBiY0oCezHGFjw+mKfbX4z3/GPSo
ZZkMDyKSOy60/QdmlMJZQRSYq04+GXCXAOpyalPJsFLGrgHcGVLrKa9fw7U4eDbuaMlhk3Jj5RMu
CeKgbCOZZXI98wjA6SCE486mhhS7fllWgdA18TFRVB9V7D+jK9QYswTAS5KHIueUr0C77lI3KPUB
XtYXVWT5fyj0B0ZSphPQO86Dr6iQbIlFYCQiRwIk92dvAu1GttUee33u6CcWclKaj+rQi7lsgwTb
/jLEFosqpBI4AOySZNAqvos2wDDDXB3BmAuVjdqtAsolje3gTEvVdIRbTILO07S3wvi3wrFgdG/J
u6firUTweoPVZwQzoaGFARCXCYrVXa6+Ku9I1Irsj6O0s+TaZ9HZXCCjceAAarIRbmwKoqlsncHW
2Npar9aHKd01v1vrRHOT3V4aXAPgwz8ETgDavUOHAuWaqWOqJpke4cek61pGqYwe5Nd5G/mtgWZr
zM4/BlNePgG/gOqesWdgB/g8kF2o9SDPzc8EyVrddvIHFyhx4TGDUwnKTQTeQDUeghgCkCIrPyI5
tIi3dmkqVX0l2hFWUAijltYr2ZhfJta39kCazbgRj7hXTALZVM7KXpSg7f5et7N+VXXA9JJRxXXZ
s+izcnO/MwMzgFNHfUEYiYt6DppaMF+0Tk4uSS2lrmVJmAgsYduwCVOrh+la5bcdUjMLT80sQZu3
n2Q1upGo5unAURXgr6An23cQo4iE+Htv8MsmZ28pW4+D3pqJa/bqDnI/Pcs3Kd64mjtYD87VyJyc
pGHvxWczc3IAhlhO5cf6C3+DnExbB4Mu6hYP8zTNz9MRX7aAEHrCHQ2XlEev5CBzUrBfE7jq0HAc
SNhbScI1jOqd2VxcXDvVwlwJ33QqPafKuyWoEPN8i8m9TL5E/mvOkXmoTu5a2/11kAK1qLS2TRxA
sV8CeyvOO54zYpnoiSIVDsdEq6MyrVVJDRjU9wWugYP3eMdtb1rxFh1yjIcEJJePJRlghVaZoIYr
0dHcg3Xqj/3HtTxdo+RaTJ+OfKrCRuNy8Ckl8sTMhM0AD74t4XsxPvl7ZOO0eDcWaiEAZLF1fHYq
Yv+JET7IhVkSydRO0klsyWJMghn+cJOk2qvMIWbkuj2gixhPlQ6PJQpfxnkLuIc7M//hVGI4MqWo
bSjsRqYgWECcbtHk6qonThj3AWMZCwqSNigK5LSA80xoB/NSq/GdwRlBODgon7r182/BbsIze9sA
R46rSuJAUYLO0a+7sdiJUb7wULpKZAoMShKWPVkN7Ma8dFIIkrdTpJX3PFb8dcMmWtjX/hb5kckg
KWgB7Lzqu93EaFgH+vgnK/XGzaI3uZmcFMy/qXtvFhNJEung2UaPtoYVqtKiSjkC9wo0V7Mf1bUh
aPtDwOkln3tlOoVFw5DUgMRS8e+habKlrVSO7X7/1KklwUoq0zatCNhBjMIyPHuB+TsZKDmEvyib
ek8glwhi90C0rSHoaIuKomPVFpY6xqL89gzglvYTwgg+BmhxKcqdUuIAbB+2AAZn8pPXUIVWERYk
H4RFNCoWr6RxiJd0P9UzMnLU3ikicgJjsrQf2gQ8Rq5Sj3hQnzsWFjw9x3L/tQUDYQ4/K7VYdOVk
A1sLohLu4xkvfPHuzY+Paxq3WA5JSBR8McTPpsuNMZUFmqvWYgsFFlYKBdy7EZ8QxfpAUXb5JRgo
9p7U2XPwDfVk7q17HdZ/zP6pnHtcIH1IatZ6TacX9+qUPD/UWZAA4XnrFkIPgz0fz9mNKvh27Qeg
ivMAo8sTbMV30Iv7VNjdlHbX1ja5+0fg2h/R6/xrZcpuFL0LuRFe0xBfAQZe1Yv5WA/oGX8vg/WJ
m9szMLyP9x5lqMDalJa4KbCP1ikmOnZeOtEl75MXikknyAcJDOld8dR7S11X5qzWMKLt300Ho+N1
MbyqDb7snSh2aZe3QAC7YUqe88IbkL4kto7klTK0Oftsgko5ytRUHScx8afLfR6RBelhdqimkfdB
UAlIyq615L/V6LBdkDRhEoL+Q3VqRJCPiTdQ3LmXaK0vGZyzyYMCvIvT0ZGp/jPev/vHX1FtYSSX
ijhaYRFu+883bU6nmxGJh7KrqR2foLjUwQRXqDm+eBKps7lQdyt3dGO8lHuh8oXtETxduQWbQz58
ATqMQDWFgMSQOxB1PUtX18ZKQnhIPtHQLlr4DxsQBmdeJh9SyOEsA+3VaAJdCIbq0V4wgzlFlO5U
iSxZ2bnBH8R85mQwHhue5g7OGoUop+5adhv7V3XpwSoS455/zRKsGdmVRLrs0mzLZU1tYjubmTOK
8ZfqgXvr6e7A6asjo2mb8i8ncOjiTS8S3mFnnuLVQFhT+/4DIIlHJJ3aURfN/tLI50RQPi+J9XYv
fuA893binhOYyEo1xOCduMzhOh1Huj2pgcWPw4HCcXW8UuBy5WE2GTRJ9ZwiNO6E3ce/+5RvXQO0
I8+eFm5Pmbj8PE5VElJ49RnX1chMHzpywh0/LGn6cskNUvD/Sd/2kLcBRAFksK9+bze/LRA7wTee
rPd6x8hEAC/vsAtlBYaIB4sSiEmqd3W1dJ/gIKovsmEKUQotxi1e1sHIyuppV7NZxWCSgtWJHbA8
F9pSWUZdeiI7Pq58oftu80BHq/CyZQd22CflSAh3LSqnAF8eTCtknul912DXyKGKqaaHJLejguXY
v1CsDAXvsgQE0LE/Rx05q5ficeQurqFG1Ygyi8WoaiSj6UYPvaCAwvKl4QadvRIMCou86rFw2H68
P2VLn3XDVLfhz9jLMsMqE6vCOm5bt6sRF+su2thChQbvePTHSRa4JX5kgsWQQaKFsNGBTG+t2OAm
bpuAczuIA9yO94BRJTdzEDALnQj0qAY7BRag55CZUjPAGmroZaGSTSi0l+QteBAiRW8Hyo7Gd9za
oauGYDOBHRjD5Ya7E/fwoPYBjeJETHXbj7Dic8w7ZfeObYUTVHoj2qhfPwbZL9E7AaPti0hkYQT+
WyfPY3QyjrC9f4LzroWs22j6CN3+iHf9muSBgzaFCknfgO9M+cXx6v1hgHgKGlcZTUej3moWsIZz
8IKXp/APxOq8bBmCPw+CPfU/bBR8TEBZdWO10uygseEBHH6hytu0ZuZ8ENXTYJSUrleIeqdTPAUF
Y5rK5k2uYAwbSqEuc9h8rhbyCS5M9psTfQS3e1y7Xz8FalohNqSqh7rYr+EO9HJQ0LKFP+wH1CJ3
edAHQwne7Bfh4zgEo2txzBc22qvEQi9UrFqRXS8b8Q8FCEl6X61cpw29Ff9CSR+ZwkFhDIn1WVqq
0pf2N2k5+mX/QJj0IFer8yLCYUpt6K9bjPua4igjKQgaXZRgNbF8Viv1ghE+w2SXmN13K6/A7Sd4
wXlkOCaGCL+VI2gPpq9cYvc3EKrzOR/lD3QyIfZUgxTdLD8oWUNTqqT7bzVIrJxQBrBxUzo6eg/K
fbHMhLFoKQPfWxOFJuQVccKGXGMTdZ9enFNlTOrpnO1MMhpC+HaXjVKGOQGPNs5v11igEnJDKkGA
6gAUqg3KoUtLrG/Hd36tjTHaaZT6Fnh6BfdeGtWjIMTzvB6WQIvjS1TySQfADjC+7HCjln6vOvCj
Z9PbceS2KRPJ3lfSt3Ht5rSa8JJ18HbBdnUqbo/HaD5hheiXU5/WqRskZxnEO9yulTs1qdk2rMKr
ZUqlMXwZqE6Xkg7tbV09m7LJH8nS0HXFToPVCa8ZkcIemQQZ8NOq/U3so1fuv2OjBvjnviWXFtnt
7JWdLDXlpeIYUDccgc7mz86cQXXalmlKBAiYAyuM3J4yi7tTBGry749ixky4QPZI8lF8nHyngbGL
mqrq5G90eEfbf96UAYCl2fOTdlBdus9+tnWy9IRJAjuZG3kT1uJ3A2kyRDyA6XoDO7+O2g5VxEx8
CH5Lz8cMHDXfaAT98nUPukA22PxQnooVf+N9kY92z4V6L4jL+dYCJW/+w0JWPt5tDxcUvNnXcFfB
3KSdO5Ci1h+zgT1WYKieL5Zrg9VN8x/dQSUMNJR7vk7o0n2suy/8YGEb8GGZLvybdUb3/fYYHd+n
BdoDEkjVKHusPQrCL8A7K7iNKzzozONiDBeNkTxYhQXMLuM0YBDTxYKvPOGzTOJocUAZGFdrKZox
jkxTQeGw8zZbIOjRHL2iWqHuewOJMa788acB1BNW8XJ7t8tAbhsn/zdyRPjaB99hgdDMUUJDxB5z
H4Yb/WDIJNEnGP9aGhsQxMON/gqZFeY4ZjJ7jSOiiGpGN/hOInGkFFYIKH35dvypXigTqd5s+YAE
ct/WY/IWTNFDERiAI5KcrC3MzyEA1ElE2h97FQOrKuQ5DCK7ar1ZxiFYdzA4yRDR5LPyP7h3C5fc
awniDWNfNxRMoC9lHBmMJav0x5N+Vv39WwmmBuv8eDfbCwIgMgdCNlyJNOGKHziS3VBxz8hOUdeh
tBTdNKQxwOPR1ey7pjHWtGWfVN/obU/LoxQyZsaqIycGhcMTwr/Bpw5NxS56kzCIvqc3eTh1dDnW
vgfZ+O4QH9RlOXTS6ausQir44RZyayV7azSnhOpy8Qv9Js8/D1GsxuNq0UQl8HCOvt2OjIWxR9tN
Ar2XiWb7+eCSYSqTe/3Io5wcaoUKi5/Wb7+Wivu6JGvGQUMeeCCDitcXCkxNIgx0blGiyYu8pbRG
e1RD6TPckEiKV1pnWTW0ngomc1hMS36AvXjYlM4evQvO3xmnsr/aho0Lt/8htLtTEWeU51wJDR9l
bn/BiXfpW41neiuJYVN7ITP9LbJrEGocCjadEZA/uGhcXvvoBQ8ACIQDqVd0cYj+RSb9RUk2N36E
8qbe26lvAL/08zZskWcGBx/GyfMxJUMDqQkeoOG0HLsQIm2/fZ7ZhK4fWbfFYV4x+jooKIWIzgkU
VUM77G7m1UKyBMSUe13AnBUJXEKeFj2MtGouBIRdIr72uakVi2E7kT4J8RgtUB+NvfQm6rFdzcwy
iUx2kkogkHISM5LtRXThHDM1U/ZmzSoM+hpWZdo1fu3quSQPMttczIkx0eHzoaG5TZ0OixD6TXGN
6bJ5JwjE4AbpL//2YqwaAzK5ay+7iGvqN14CK+Mr5+PYZQ0/V8fSG4RfzyTKjWHu8+nrHN0y+aur
qLIZqizHvH0wEuCJtVyYK/NOF16gZOG8vgrKn/J7MH8Ag/S8wKUbAyEhJlIh2MZpPTxlbCoZBhaI
q7hSCaGLiT3ulWQVIsAvcbQhZ8LkmraHEo/6mI/aGmj0ljuooqGPaVpHI5nEoxRrN2zvyZnMSSek
V4HMQR1IJhquAkYmRcR+Jb2c0qZRB54xudcbOIHHxspK4XlqX1asUSDu0KVeMLJ2X2rgjEj6Xmzq
pvng1ZiTGq93FwUZgg1PCHfA2FJOq17yPWKKwm8apFM78w5vXXQ4XuLuj9eHEuicfiEULTggBOqF
Nn9/z70DTY6A7Y88fkKpkoKd6jHKhjrkGY07Wii4LPR08Xqmu7rVCH0D0FDtHY4dIkvfsKWg0wIO
QsvGu3qOJKc11oj6nDiNgBCbFdiTwr+SLdPJjTGG/in9sN+cGZ3FsCvlmhmduaqCFDD+o4QBAF7Q
L4A+yEP93StmG9g4pEU2PMpyj1O98GvpTgohW2cp9VnLK/USnl3jW6ag3OfvG//pSIuvzSEeBEck
4x58UypdmNvVwQhf52K0s4hUqVlcy76f75RQgX46Ynh2hBdNPVuIQTmNeKw3Mm6LHVN7szQtQvIt
MIbZPGklGD0hvdHmnekNa6lBIfkNee06X4AW8e7zIo6Ugz0Vt9KoNju5r4RkrMKz4XpUK8GVcuiJ
HYlawVdfo4lxJWvIx8D0m5uz2U63OMiTIfxnHpQbjQ73VAmaDnn2wt8CyiCGMU4Mm+uOGNB5ldhk
7YYgPgjMlSyY/YcGVSefigLigjHEmw+a55oRK+eCiLyyZfhovzkfR7sGnU+xAx/nwOVMek03zSNE
mvqIfYodFf/ojEwzWXwVkfaJA4tD9TvKzhCAgnZbkwGTiayNbqQWu6fOw0MKo8p3fyWTW0RPCKPj
XssbWnNLR6ridrT0lddBs0vcb5PR5l7VpmgXAbTvdTHYkDTrLgb/QF6eBgQC38R00Sf/7hhdTWur
6XsEi5KuLnf3FZdsNhgUs7Ixoi9xEbh8WCBmUprYdVNSU0NZlQhNrwGovpU4N1FWpCgQIlunz8OO
hcoZe8xMCpOBvdwAsnZCX6fKOk4o8pnUhHAjkLytSCb8iJu5YRTvl1GXaXCs6wZxSlBJptmHB96d
dKqXkLlErSydSwBGujgcwAPkKO/apMNxpwuhlW9+lO833FgVgYMqTflv44SzH428bg+atWTgDjCQ
OLO7cBfrQqwL8vkUsEf8+qVcVPzC2nDdwaI4YY5wUQhJCtRCekGYyCl4Gum02QJgrlqGtDPf0Xyd
5H9GJ8WOFC9KQU88iqJgem9OHB0HWu8zB4QdapOnYKBL5DDB5fEtmObNVB/gcjl1/t5CrSiSEyxH
+tflNdePvI9ADUOGWSlC8WXe9p8u+S8AH+Cpil2ZgUSm4fsP+uDkIk5dCuWUvGhCtTF//iTM5vFz
Z1QJTvJEAGpjmg9BjWFF2NG7+X8YHljFRmGhgbpc/KVq2LHfjHlxFGdDjaXJt9mMNGA5G3QL6cx+
WNzQmz/QE6rMpCK5QpVpJNrz0tfgmSbmCJBtvDnhPITF/hlapDMOqD7R6j3rANQTC8P8rsWZOvfY
9XLSN7id6v1vodNbux/XrP+Af98lZcPbzufgaiv4D+ZtpX26cjY5fx1Cjl/FjIVUD0GdagCcDoug
ak+JTvmFzYTo7fd6Zv1L5ReehxgzacEZxiwRm2aZT3aFkmzJh22iO7AgHPiT7CKC79PFSI2zqrCG
+rKqS4lLtRNhnYBeFAQSELWYFWSKyPM+CTOpcT+CXdIE/pyZg/AvN6ar0ktrSQBGBQgJYiAAFIeS
Xjo51ZEqD/qgE2Wyq65cW4Z6OnH4kDtib8Yn3HXfqtvgy09ASD401/1zxKZ0PNwbeQS0Wk+SE2Fk
4xKDNlxhdvYFp30iYQyNmZLZGtTh+fZQ9R9OXWgonzM0yw1mj+eoEzejQPRdb2P2x/RhIMgXn982
w5HjCQBbn0F1qRd7Co7q34e0zyv3+E3f+Zw/mdm6euqL5B7Oxrt/dmOTBnWic6R8OocwK8GfNHQW
Xc6fArXr3OqbNG3OzULz0m8E0k6N/2JAK5TrMb8gpC3iCDv85lQKr0xqcPhElDvrOsNMQgmLxCOk
XXKxW8gLfKqfPAExL9nixjBs5DeMP7FhxtW8tJL9r4A0EAupQJIkV3QrOMUxvvTjoXH8ypzdbEJX
pitPZzJakSMzjBiLXN2hDFDpTnEfSMzW/dhcsvzynKn75/Y22gRbUvwJNpb+GjgnPQD7nTabF6iz
d9s5MU+NV8a6Nw2czYeHAkSUs91FZV+9PphfGsnHp8zKHVZfTUrtWa9EZiNINGY3LS3xkTgKzVTz
WMjznlMrNU9f31pQB1yeb/eDMUv0LQi2rfviwmUmJKR4bJQtUixWeednCuSBTbPkTlVP9HJfGZFn
Xrx9S0uDo891ppxNvmk6ikEJWyCemsRbX1pBKMswnuUQ0FSJE4y/QQI+rtHJo9vpX0AvLtev8+Oc
aJWJhRh+CsveKw9JLq0wQ/ZXtmFNBLb8+62DgxPpwroV/rridL/N9CWn4qTPePlqCzyBklbEK3XO
NsbZM+OWL3nI50+ku3lE4QYkvpWgdRIGbt+OqkIHbLJ6KswqGfBFplucQYRxLlQXAZLFBnPbhvY7
S9q3tludKfQQeuxccqLPaK2JCTvioqIeUg4KabJumFK9cKofF8CusfzfDMBEWYfGFAI7MSMrgy2h
s6yMIMZfD1lYvBFyWHh9NzIzGeg3CQKb04c7jaG4eygbWBWyfBpA5+/NbU35dtsTS6RB6lUllpJm
nAc1eah4fTKVEuI/VSQ5vewlEeSHWC9RfQLMIfnOu9lvy4+AqeRsRawOUN+nDEikr089jPqTPXUI
Dq0lxShuuF8aLXzRGOMHyFUR8mmXR+1AOXG94S3leKYfyKILBl6tOMe9u4H3XTMyG0bupUAnsQ49
MhvpRu++5TipDGHqi6tuXsBLHrwUwsjZdbOqQLE3B4CrjtqA+j7c2xyZcGGSfMPBp16Fv6fin8F8
IqGnLr0JRbHqqo+j+VNAXlyuSPvkGXxKZ7Yhs/MyjPHC147nMGVMZlz6Q8oGQQZ79M/jfeJ9V/vs
M3oorkiGtqEK+wi0AR8Hw/0MfOTsNs9+L/avEftoHylTCvc6SP4he+35//IUMe66zjM+WebVR/hK
H+lIW8tHVwavNSJmZ1AOCu6O5AQ3t7cKqEv5IQTLfneffwFo0q2m5Nw0WqMdFbu9qKcS+9hFv/k5
Y9G5CeuddMcIZHkWiuSmY+oTIS90ILr8Y7JQoRFtoC/r1dixp1ny61olSmBPEyokjrKVx4V2tjix
hBe5oc93HNSB6H2e4PGiaoPEA/bx8DxHdiSQI1zg4rBgrbJIqKF4TBS5Wkdt83ivXjZPCXf72wYf
JMl3nB3/t3rlNYd79Yoouo4vUvGKU9783LD5U48SJfKGbm/TPGQ4kf7MMUjBRprCm2myQ3fBs3vw
QvMj7UQKANe5ExZ7KUIjR3StIL+YQH+wms6UcicKRecFumFeYDqBdrWhrSh4EhoLAKtuYx/pqeYJ
d32vI11TCXRonlF6CLNVa96Ge6FohLnRj5j8prt6BUIJ5fTqdHI5Ja3NSvcZkPxCXrrfEw+d7d5u
fBJEyoRIzCsMJqFyCXPfV2r7Xu05PbdxOs/vV7TTOg3lywdk8rR4jia0fu03rUY4yZmUF1Rj4V37
xMr3POdLLYJ6fZ9HNlxGX8DtilErPE8vKbNf4hNqb9/fwWJE57OGPIEX9GK+fY8GQACNxGeYlRLd
IVEZZnUIKY/CSKgdYG3mvjOwelmQfEJusZlPY2QOqKVfsCJulRqnFarm3vuOk4N/jjgFyZLn/x54
VvfLRtMTeYLbRfYHExvdWWwfkM8+8ywpstYn/SiTA/XOuXWUK6pYY+/gPxBB/Gcl6xbi7PajJNId
V/rTtgOyyZOkPpFGuC/0fpV/WRxYS15NvfzB/FRO8zA8njZEY5ibfESwl58t9PdCJIAACifq4auc
+gT3iNQVH9FNtjCxmucdCHephLSb8od6DPB/nhXcxQwk3EClm8N2JEKYXOCKiKPFyctylifMcKop
DDCqe0dapbRvJxv0KBE/kOEFPHFBf/UK3pE587cUJUz1sNK/2le3k0vC+D+RVbTBPDgkZHpHPbe+
6C3Py+4S4hZ0NmzB2Uo6j63YSfvev7MrOsYGLeNn3Sr9TD420HDy8RKDTGbgEPosQX7UQYSf4LVe
zkrW4gaRq6818rD/4sF13LEhu1wXhtAjmBKkduSojZruEOxVKdV84M4A/Bj0H9tgzCsNcIqL0Gfu
zUZU//1/5FWkjgw4NRzXWDp5M33X7Bd9eMRs3EHEUPyxTQCN58e/FNztgDSIaMvhPREV4F7eSJNK
/rcUjkFIW4dHNNeNj0OK9VsHJJBFk7X3OGQ9vavjzDPYLFwj+lz2xsun0JHtvr9NyfHK7b9rwT/B
QYdA6wxhPZYPVjy6RwKXhdQfKb/SBmu/43dir4u3wzSZPwUyaWTpv302wu4Eyj8fm44Qyqti5+lH
gHaZdJkDh1YZ53oihv/TSRPg6miL0Nv69OZ7d8OQXLJEackI3sMdwExtPQKioS1t5JK8tFxZkRNa
ruRanvVdeD1qVnxAJtS3ZKCzmvWFYsYXr1Cyc7SgsQyzkmHZ3jLzZWc9MtqSMyyYP2usfjlht52L
xSev58bqgig6bz8cfxWAldOV0PcHaHUBPRqcEPpWzs1q40cNOxxeHCCF/tr08qiF++Y95rvMqVJL
B50xC5ecRqrF90JLwJ5WZVrM2WUgCHKgr8B3PVBoFWAMKuHtvTuvKbi7aMIfPDRG3CFm+p6iLTl1
VUzPv4yUZGpG+TyIsuiRzgk72GgNj5cYMz3nI5BJMWFWd4kl0mDzDZ2WF3N9dh9jRhx0vvpZUUQG
s7IeJBSSWqvL9jbii9wWdkc5PS8+2tHaSe+gduHjWXJfDji0doLSsXimRp2uhZk19tvtyDjeyN4u
pGSVaSj++FDP3Y2VbC1TM7ILf3mGAxX0ONA0WWAr4f64mvACXiJui8T6mzXcyF2sgkHl7X66nzYw
23a09trzMu5ZRZH1nhbQaLwmqoibCbduwPDQDFvq+0Cbcjxv77+JmVueBvhkntZUYpSjiM6tD9e/
uA9jdt4eWyWinCXaCVZz05dJfd9TVtow3YBZug3briptAIF4pgS4K8jdGIyiJS0Odx7fxmwROpeo
pEWoBKrWowpd8IxeCv8QClZBFdcWtG3jA4OWMRwpITuG3/IMwLZtONEYELBWiP/4JtP6t3zjKfs5
aPg2XPzAR5XcErcxxy1a+Sp15BgnR0KY3AaOd1NM0SwPirpkj9iEIUhdL9ErXqKSE0qS88aIjJho
QEHAajCBQ8R9O/bK6KkPp1vNcSiabEYlWg1FnuQ663bk+r31rrQopZIEfu6nY6VL5wDwpPdlItwA
wnTG/0EaxY76vEQk+MvvJasrMp3p+7BZJ7vbPYmkp7MnBncMnE6/+aawMeXltbjID9/vVPB8mnDX
32p3Y4jc3uc1gktRlBceltvtpq2c77tzykMW4FQZvQMo24sqc29ETIztS+4QZLlJCpID52ci/73c
6NiagDii7fFticbIhanEtyi0SbEc9WoLX+yUxiiF6K4JdhOGN4St6kY7chZsQipW7uH1Vn50ciW+
O91KFJBzsfnPf8b8QnW7it4+VCBPAPosO+/E4Huz1jKcgg8Y4k4gKBBN0aEYeAs7v6mLR8dpAmiE
aQKoQxmDQkucfEuhEybjtezf0pJele2G8DO9eezS+HEDjSmHpakke3V1jI8GdlJsZPNJ+quwB+SH
PpEU1Ipio4LYmTC5J9VZfrshIoO/FcSE82/gwko16aa1AG9e3HwDhv28O/ZVtd2sB1cjUgYT1HWj
A1HdP9+XL7aQEHAFQTsPK6oMXcZJVqiluew/CmRl7f+3e9QJAPb32xiwJ+8gSuNYAXzIsfYcZuvl
0Rdzq9ewV4EYwmb9gUnlwEYU6ZkEoDIDlxgOIjXWUnog6bCHUOkWYH+mMAkTt4k23qZyoHqVRCwd
kxJ6WdOgAKzDj60tHY71y8ejTXr/5XxcmC4xy0OThYglm/Gpf1pWUcSZst+RJqTvnQQ/o0dhkm3G
jVRRvbGuoGwrBY2CDjuQnii2pmU7Tsl+y72X3kH8+nulNc5ye0pGzeDIISKVjWNHsHUkJRFgsXSH
47o0SGqkr5x+ajhlL5q+c+UEtIqcsd6dZJh6PGZ6YYogTNZ7TlWibK/CpH+0I+1EinQEFhlG0iqU
ygSed2ggemua7w6xDWS6upl4YNL+VR3MLcaNSF8zlCjkL30jfnxIO3kjtjpFa4x/Zvjc7MXu+eQN
7/JFgk8Qc9j+RUcnaYEAyI8bSKQdfqfA17yIYwRCnTSKfhEWWNOBsBeezQ0ACZaKKdNzIE3N49IY
5MQ2lG8TlJpRhFcnOKgoFLj95xe0WASDr6UaDjWbtbngRrj9/9yOp+nuEIh2B1Io8FwopExPiyFt
gq3/LbdB9puJMMiMi1eiYmcXNmmino4feLx39w9sBt9ozPq3ObzBV491Fux4kUDQufSGbhAG9a7O
qcdTLDh4SA9GluBZV0v2VskSvWYk81rdxGU6o+MdXIvICitFLNO0bs9SKVB+510O/GP37C5sS6NH
1XIWBbefjvtc1XAb+CUjTmLZP1vRdEUNsc74IkG185YQ/eO8KHqpNpSyzCpc98Qq4QIy45gHv2QH
LPmbU/VnrMWGzWQHHgqlQtyw7On+6Iabb77vRFo/ecKOVE54UVe7i6AY4ChY26zMlL7PZB6i19uu
GIxliN1fjCMSLVsfrRD+OCMx7bT/BW/Zb19N/CCZUY1V52rcUXV0WLRItq+mVk52DHwnKAdIqv65
TZywHZ+M7M80+s0wuqwITc9XKmuj7NjcFsV192NcEQVfZamyRDrWQaCJU4c8lyMZp8gPuyHN6G6c
+gCWXoC1JXqK17ktdHdWSbbMezQKawFeUnP4ZqjJgUqHCMICBwokDdES4pL9qry3V6vFS3ST96yy
qA0bZQPxKtjLMJXjKyPN1moItsT+bmiF5cG/3RlhUehvCx8OdlA2hs3hR+PujVI4Tl45qA9JOG6B
/97Ju+ymlEqe9j0y2XUwVgFHq21cou0zk/MQy4v7vXJ1zhvWZXiZz7PtX9zCq6ReihMFNVmw9/M+
bNyfQSmY8PWvxvw3tip6Re7eVNgiIwt29E5qy9mX62/1csOjwHqz4hX69viYSUNPlaJQXeQQF5ND
D5y4o3PxVmm5Uwv54aVoIxmYSZZjsGPbrFsFqe+XBwmofJSj4NUpEi5L43xq1z63Q4eWx0dD4GAM
DyJLAO9wOIYRoQR7jzItPhmHtWfPh/AjeI7d9ufVrV7T7LmKTCOmVnwgE4+UAkeBqN+CgDUxL42J
f5K/JOUtLtCS/wfWSfsNaI7IvAYlsOhO2SxFU3d+w/NIP6AChMYfuseUj+ugrKtST6oSP25+veGK
0nO+DjmTq8O4Ps44jXcaiHKuMiXP891CB6EEdYV7jsIlGHpFhKVCT5u9y/YQxLllL49DSQAXVv6c
wqRMYzBkGTs6JzkbrdH1fgTP24Ia5c0Ld1hs3gQZLcznSV7YNppXT/aK0sRWKawQzv3lPoLZ9ZTL
Z4haWXTEhHZNjOxl5vhzDB6A1UwcbcftI4Z8mOgQ4s9494son3AI7OaQ7o4CdSBqXYeGJQSj1md9
loKUC5Yd27BzEbriz4iy5fYWFQfKFtBgvNUxBRJMM8gEWZEGOdxsGNIYFMD/DvK/Y0gbbb+jndxn
zN7FVKl/hybJrTPUDWa4QTr93R9y/TQygmkVOKgj6vKRRVLhkPciaorD7dI2AfBHqIPn7dJf1/BR
dCPmqqBq6X5Aee9uIpj0GZADf486RzDdER0nQ1f5yWcWeaSwKkoBbrs9CaZo8tTtNe+lzrelpRBN
zIOUKbfw3WbEb/kzLYsBXzHnTS6TPLa+Yh6i1MnksNBdX02WhJtIUQXiXwnH9l+n15w2SQfyc7ZM
588XiCmqrVgnmBm4soRhntim47j0W9RkyRkErtrxP/bnBeYXseUgzAs5Eu/aSRIwkLR2q/HmAr+T
Lvi5eP9zcO7lesgvzcXoNIDB4CpWeuebDYU43nXvlAkddk0ykPsm5utsVaF26Cz8RmZaQ7wyKWkv
0dtDFBGm1XOUMJcFjeVVstS8YEzsExwhW8lFvd7tmzSjSmseNtl+UpVe2rdQK89VutFXwgSzZsc0
+8DItwo2Vupv9rAusqPMl9eJWC1SkLp2QwY12eTdKk3qrdgeXfbH5sD0frE+OGvyKgVWqer0cS8I
iLuiSV8YonW2j3oyuqO1grxpQloV1imtoAXoymv5zvgJVNNZxltv8i+/Zk8foYbtX+XpaPHZ5B3Z
qFScMdBya3aLj57cLtLlcDj79/h4gaW34gp2TbuJ2Rs+OEEvfEj8pVt+WzIUnp8i3cjQ6trNYV2U
1jAX5m6qlYCjfn5ne45/lPh1dsvYX8C7ym7tVDTS08gVL/E5AmREshm2Wp41lz0boLszD1AFMhZU
gABPwgkbuEx52jIno8RgFyWcweH3w/MOnUGESvlnzqoXz9CCGZ9uPsCW+BtEBTZOsELa6Qz8+Jrk
573ZwqGbS8XAfkHp+UmZ7sSCM4bPJq//Q6Xt/UAO9VSVp/59VvvXltQgA1M4kVx1K4VKAm1cOU05
+vbthRFmfS4ztjVT5QrJBmEq5Ns03w25m7ly3nuDgOuaqMH0S8SdB0Ydo6VL7Jk7Qrzuj+qXRZ/v
3P7cVKb1MP8EMCF16gfxlKENjL4sBxbmV+IEdPB4gH0cWGhCV79Kk8ZJvGCq+sMFnDEjpKBNSSwZ
EGvqfycZHCkJ0AzwJOrIqyW976eLSbSDNnqNzMpaZYRbj3knyuEv2SHrFR90xYOliwlCaEjJ5jsu
zuEQRkWSSd7YM76cNzzbdMk3PHTLYOdGbdKm4AyCwc4fTnUJn7hy80JM/UW8Ca8AembkkfsIOfP1
4KCuHHzand+zG0GeJE040oTcNQ5napnZTRSo/b1s2HIEY7E4uYeF/2c8fO2xw94NYin8F1zpxBUp
J4Q7syajY9sJNUiBx+OcVg3H2J57Frzif0P1flEkimgMaA6R9FQfAXmTzHL0n1NFN+MZLl8zUETW
WXC0cGBSVJLLxA0EuBeOjTt05Mx4hEhmU4zGqw1RZ7Xz7D3iGYSV1cdhJL22qxwuQM1r4qHw9onO
jsKsLF3vhKIDE8EgW1si/NQBMDc+wRdLVRdbpz7LQy/MvicYNwDEbumeIR3er2hzSVhHjYsHZL+o
+RiqzKTHRRfCR8abmrwWhYo0DxoN7FH59MnlEqXD5yWbqRymKdWpu6VABTa44alNeYTXngtkh20C
n2/xQICwm+X1hbwffLKMVTIsQN4sCZhaUKWHW3zSsSGJeHkYY8EFVJFAabtUzwWdzejzqJkAaZFv
008RaKDnY3A9OLNPd57z10/KEVe45E+LRM8o8wfqW2uiK9GXf9CE2MtmF42RfNkCauXeRZebdGy6
uzYQwlla9DBHsKr386NmoelRfU/DGEwDuoae+sjlkjJwffkXFCXrKA6KYqQT2Wsafzi9LMEvw+NH
BpoZ2LfLOkrAtothURVR+uGAcP+8EszSRkhgs+OeMRMZZqS/H0L32iAO/WWRjJEA9lwABhgJDJRp
rLIr41b8T438BaLIqtwhCXFAQNCQqeZiQiPewryk1J1hPi8hhBujwkHOKSqoUnLw5UexmIaypUe6
9z3aOMUn7XG17Fni7YLHbsLPo+XPat8kzQ/019jk00iPSAWX7f6xe9clrWDj1zYtM/pcX/qqtLTw
qCpDY7Gzh7uvkUN21nKocjJAKBcEB0rfoD5cWVxkr+EwY8/JUZVXuVAF71djm447McL2H9L95oU1
yVGDc9SNyeoUCpdcGrurK3/gpkAfI8CU4s0666B4rIzNV8XWec8R88T2I72j5jMK1G4RtlP+h7Ja
1JeHbrrf+FprAZ5WOfzePjBH1ZcbfRqMp6HGFuAa0bwiEwAUzVgJhGzB9Q7RAmqg210a5L0xqO6J
F/JNJbYCUF4qrGqADwAMJBnJxKm3YyAoCp6jZWzH8E4ZZmKLGy8VT5g70+9a1e6PdvoKbLVX/Jgj
fu2C6OS5yyAyd1EUcS7mqmgO1jOTpR4LzVt4MglQ2T9YZRxFqnRTGpS516SgociAex9WxX9qguiq
FO1ClzMU5nDIMySebHOJjI+f5dEt2Wr5cIa2+ZDrF1EHiAJ//PViPymNfGRiYXSNVu79rfr3p7oD
DEpl9xDD/5Zt+s37OHscjsh8PXMEplQv6kLDfoGTMLG3kwplvN/O2pP/nvaJBbPOiqDHpFQ5n12y
1NJ3L6oIMn6tnQvZ0MR4hDAzJn0Fjb92z88RJW9ZebUztNLlxv8u6tCULXw412NJYsEXie3QzkEu
wMvXx0YoGxZv9hmfJkonyOGKds+HpJ7mbialoFcHwM7g9qfxzy0QydpgLYSeuimo9PKp+FvwKaFW
c93rQQGpC+erBptWEoDM1wNa8rAQJQ8ySgfTr1T5Y+MxCFQkwX9YvnNa22mJNcCNwQRNGP/Dwf2D
WWMci6tY5MSFzf2vwrkvKsQvibDZrQ/2DbWMc6oF/i3lnJKS0dIKd72hvWJwnSfiqIvY84YHsppN
Fw+TvVwOlMy/DP2yjq9Ei1g0i7tiCJ4yhTuB9SfGsdcGpGsiquSUf+5iRRQ4JbiInw+ZQ2PjmKRw
gbMlBG2aXNRHi96WODbst8gCUvz5NDHxbouVlxmJY9rcwI3aT9pQBjZtJtDs7VoZibjKYP72aMDR
AXl8rbQFwP3NsAs/hfYh4cLVCeVAOQpQ3kJtfiCgwnLYXgtqT+AJS7+llmRg/x/cVjxZEquZSMaC
lFjhQ5SPNERZph3pSvTSZISJInzT6yH+870rNpYgW1I6m5qT04KNThqPpEn3mGS7KSNh5DibM6Yb
A55SEE/KchUi+lMXlBhgL1GsTrNJE/vg+VnewBojB9MlFc1BgvWewA1ntunLMiNfsi4XBMpSxeIT
WLXk/YHIV/MB+PP4wcw5k4fBPuUpRpPuxI5PTDVX/hq7m1PLFEyhStdTbuXrxGeMPHaOf04vkN0N
4cyTp9+4OeV4X/bHGg4A7cJsDE7R+ZbESvYVUS0pps8D65O5e6EmRnogTmT+4Bfq5e0lir6I1/Ur
DZNl0+mYYyWpCkix3EgntYjs+mn761+qks4iepNM+Xwni9YNxn290CMmpoMdrZQmuSBrBgp2nPR8
jYHWLZJ96OTtkXdl6E6kDuZ5P0RhbS1VM8w5Gz2gqJRnRWpe8XAVo/uFGbzHGhjzkZKDrjI8V0Cv
fSWxmeVvutA2lTUlrzjMEkDsDABRCXdBMyEti3N1WzP1duF5hDCY5rIpdxADPdS+ivSAMNypwOjM
CzOQtYfFovHV9kbdZn3ooEt9+Mb1d75gTXHQlgHdGnIiS9FK3X6QGhIXBztnbdJrb86dbaQZ3ozf
fof+z1f90s9FQ37tW++5aoNpjWEkkMiaGFJC+cZaGmxKWTIrAvkkT2W6z65KjMn6r2eg2YA4PUSo
k0PqkCoDno3Rx6offHFNGS997O/ELVXDBdJ1Ehspr8dxlhcJPo+qHP6vjXfyE4vVMgqdUe1D2/gV
d+Ea2FJsSZPEDUt6AhaWWf6BhL7o/t3+5lp7/ETUOvgYZaE1B5nQGWAOvkJqPFOmsQHAz9Oj0o6J
wCRo9VpODQ1sLMQyGu01GChGaPPjq06nQpRmEMAtrPE5zO/Re7L47LqyS0TTCMtufU1alp4Sdxni
oDp4TzG6LOKPoDRzV0jWNEa3b3CT5mciI8yAPdOXWQ0rocD56AV06KFtohVqoxX6qYcnGe6wSWL7
JGoSV7IDnOwqh/7/MpyVJ3ZKcrWDA2z2ZUCPioxKxSNvjQ1BiRkXLZIaZ8VXweP18H1q0TF5sV/+
ADzIM6OdQtB7cNfyMm+2SJHu5hrtga3WvOxQzwWFslJqZYksBLT+ld3Y4Q67pIXdi5C0A8ouGRlo
Vi8dwNuCvLfJpNWyNYeY6Pmpbne7wcga+cz4BHPVCbyNbNV3CoEB3A8dL7tYkrycwW79qi4TWD/S
1QwUUJ2bxfYnJSmynNEfr0P5fgVRPMnSCtUISbmHuWP0qy/re9HESb5gjkysFmic6noJ+HX/6BCT
kfG1klsYcH6CjNJ58VcnMU9CcIXGqSzndUUfSVW0TPnsnnfFDl1pku8MEv9cpmWrrbwk1WCYsYP5
gyrmkuVX5T9418K/QeCFgNbeGnauzynLpkgZuCz/qhp0gI7Y2sTYB0fz2hw6HYrkGHjgbBBjq9nz
FSapqQaqF27PR+W3u9jdspOddXxlMDYgncPcAn9iAZ3R4aOlXAnI28WBCaW+GyZ0Bjm82SmQLT7M
kXxiyd+fK+wwxuhrrtsrft73YrDUSjdRH2XM7qHTYNTNs8wc8LQQwsPiymaSqcts8Na/VOkUrNl4
5snX+DPytqwSJ3+DizFXT/akWXKAz7qZC9BC7/HrYQxByEjf3l4vTvVRfS8dpXfXYzhl5g+KCr9o
abJootS32EAM9icmhY5Ie562wOVD/TI8IpSv62kjQzpHQMHX/P3H1QUik/LQ+E3cxHwfW5nutGY+
gJgBRsIG28ZTFr3zqlFIvJSd8fbxHpA5lcH3xZwkhB29Iz3vZnf5Oqcb6AVD7b8S5upbbh7ZdhBv
G1h6E42g4f8EfNupsz1IsbiXDFn0dfnUu5i/c5AGA1FgdNdANijMzL/OHCthcJU6T+R7yWc4/3r8
UZsDnOGJEvgWQsZ9hBXBOYT7d253hnL861onRW2w/bOEBeCyg40fsGZo2oYPhNelAC6vhUb7RYks
os4z6IZC+AZT8XDwxbQsurAWQL9QQBZenUVGwXJf5msx7b2P3f2JtP3JWSeJ0Zxjg8Gt0h+vB3b6
9ewI3O5PCR6ORxYvH+w9B9E+gEptav/STL6jxdYrm4KUd27mVNti6tJ/ABPEujzsXQM7el4EmeQT
LDFw8WSvDhQpcVSEaVGo5ywoOL4Eu3MQw2osgZmKT+i999FP5RjLa8LwLgZ+aM/Fk/pmREnLNBXK
98DjM2PcraMXdBMZdvL6d7pHgSgB71siLuRTyb2o3ZLgTEl62jejmgEnHqg+Rbbx7CIW5tyUq9bt
pyZyJtSw19BWE829Z5SEyvNyLL8y3Leto7V+7ty2IR6stOZDHjz6kw3zqWaXcVPNl4BL4Dqgm8Qe
qGQSxAjank40lunur6BwKBzYTWQUBKoG0fPmOOE1ETAce5MMSH7sbLuOWxpA256TD3wc/LrsWJbM
NZXmw50PGA7lqE9IDdaSWf1qrUJnPCae1B70NaHZcOXFWVjenSOYHol9EWE3HucxckkGrCbfsLI0
2hZhHcyOF0Q5UCWyOeF7zkszddbDWifrA9yqw5w364OjbMUQu3M3j/aDG8eW90XK5xGi7C0X476o
DsVAvRbXOiapXNyWvGddDmXOTnCGFqmwTK9wZq6wX5eRdKstPV09zZQR8Sq2RLLPSJyXqVPiWx/n
TUjB1a+m3AJ1JvnWnkvUU5jYLfIjEBmzDnk+rHCag4FFgCUtMKsrpDKWTZqYJii+0p9cocA6bC1C
GwdnNr/xYaRPdNq/vfBzxaj2AFfDT6wCRphVJrk4G1TB73i3QBF8APkkg3YBPm0xd7oiUqaJGdMi
/H+thHFi7dWb0Rm3S0u0epSC6c5CcnbuQmN2QgH6W5du6ug8zlQyGevTtzgev2S+4n5t61eDiWC+
/c3+D+WMh9uF/oRAzCihfEuAbVFjgYGWU1Qbs1M6xSvCVm0K4QeZbRbRft2/1xXMruKeEy27XHQZ
TbKLmP+aRA3e+l90HrdoengfXPI5IWVb37+9EhMZZWNCKLmFzw4388/tnU4GSNh6IiL61bJjtPxB
yc3XLreZhSYgBNiSN8xJIeYt+iIzZvTp2lpW2nfkOj+k9mfzSHICPsHRcxk2qQR7Yz92pLhM725Q
DO4f6hRWBRqupUFXKuaaVSgimMGX9bhMj9k4ZT/fyDpAHyLXGJhtr0GhZVcHxuc98PhsusE8EnN6
GqL9pw3jVhrEgwMPqFA4jhz0tbwuO1ULOzRwR+v0ChUtjhAuX39yy8v9iIUN30b/O/fxjvDI/lh3
BYwgv6uG+sUtGx2N8yW2zVukKsnNmckaOGGHM8sRvNtfuFZ3+ov+PHgrzS/rDxOLQfCnkqcAs96g
k8vydJDD4l7rR60FOZHbVwuL/MaHzPf/2lHF9/W8Gsflepe+PmJNLbe7ZlDG18HTBF/B5Pkz/Ahk
bO1m5vs/5Dg61hTCBVwO538UKusHPfmFu8IpE4ED48kEhDSfdkMAnTThBoMbZQoDvP7ef+AsKblU
BSkqAkDMpt8iCioTYBwmsjVIVpoh0iI4arxAGixU2QcL1pfROe/CxPHUKo/xGa4r3Cy1BKXgK5dx
OVi7mmfvDmUl4/QXF+YdOPtEoxWuQOXcBLbE9AJfikbcTcV1c5IcEiUgs6k0EgN1EbkHiylB1av+
eQXx4OdDkpruF/GBaDGFXu1PqKnQlVp56Wc6tzYfKZjc1in4rz/3yLXJYSmR53Dh9ObIwOst4Qlc
YQk8HCYrRRMamuC6LTQQKv0mcL/3D6tnQ/+3NolcIrR0c+FE4b8p7N468v9H8pCKSrpJj5QsKBz2
HEAMIVlvLIOkfyMRMBUkiQX3POODyy36ZlhMYfduEBPg52+aF0EwBPi9B7qZNnDz0DKoh3fYMHK3
JkAlZzivLn+TFPmrQ/D62JAwIuWZmblu/1QPyztYFVXrjJ+KpoZ6i5E6uPiUmfdxqKxmfs+TSqny
gMK8g3Y6pnTeFXsePkXYJtnYsNkJELS1LhZF2ZC5QbGKMk33R+NFCsM+6zGOk2zh829Hjp2XPDWw
ZzslSg7iIl2HZ5LlDsUo6SkGuENe323byHDisO7IV86WVubP8rgUFWgaw6vlBIZ7rTmHQcRN5LVw
EN3+Y/GJjycgqbYwxyvmFANt4Z6Req8M/nIWnZ53M0df5bWTnicqi1/8IprYzbA2OdMxLgmkFbIE
3fq+g9AwIKXPwGC6zlMIbdAa+NLJAcCoSLhyDU37/EkRN43Nx9pR0npdeRuNziBaA/PjPxOMMSya
bzxfKuj34JAW5LiZb69jXy4x/4waR044uHswu55MttFcrXm4HjSmYk9Bbfs5O1GJCMzb1PGYlDCd
kwx/iV9s7t4ZDMRW/iBZ8iQtp9aCECixk/V9HBml66wKMCD3rmvnIGxlYBFOlSZUHuRE+a1lDKLu
UF8W3YSz/G+O8xMYxoKX7mzld/BP2eOJFZLp82i46aq3QZtdmO2afAH0QcLRAZOgtJK4Dsnt4oLt
FulX5tG9UzzXvZUT6GdTz/2QMZbfTzKk3ZuQMEc4PmeqDJn/Nl7L2SnyeQof0q85ZpOutcKWiMY3
iy0/7SjaPgUzx3DJ9hF5ozcJ49BTmU2qM7aGMvxP5e6sr26AGLXiCQV/YvXf/pjxMroBDpa/iwMq
jWpAHfOs+Ly53HxvA4FgfQh/inu5C+Sb2HBz5SsoIFAVwGkSDFfOvIX0fZ+cF+tUEHbc/0KBSqmG
0+zy06jvaeoO1DMGGoZO4WzhkR8lYrrJnCCADoWxoZm5fWnwBL/nUJRgtgPgdljvGhTJh0f6CG1q
liNnVhWmAdPJKkznes/AqB1BSTTRQtw2UlDyOVkHadQC7g2NrqmTYRqmeiyvq1WYozAVp7KIgbRW
F7ONvosynMcd9dk70Ga/+iKMih/gqptW4BeFHxvQyHiT4KeBoLebWceC1Rjz9aztxkxOrv+rLCLs
uO9uHpec+TWnHFWhKUWUDmcGWkBPXCGFxqrkcn21Llv+CmlMV3IVWIN/zfebnwL+dWHKt3nOZqlp
4/4H4YQUlR2tqHvOa+mMUw2X2dCWhWxHQzjbkGcxi7wODdSwFK6emvRwzxe3ZlAA1zq8fQLhICbs
4PQJVOio5bvDk/GM0BgHMJfdU7JZyojvsOagjNuCOuEGxSad4vafCAN1jlHfD+1gbTuxqx2kGIRE
ril9fg6YIcBtZ1YdZg/cpAeae/wz3eDxK8KhyOpa/6qiYML4VHb89nYlp3XufEdXaRBMHMBoyf5F
UrkVumVL1turoZhnYnKAJKTng0At4cFxsRWVbAspk6rUoRR+jIWUDcvKp1TcS77lS7pDiFoE39Bs
Q4PE6YOrxCNWhRFGnQtCu5JdLCVKo/WSj3T6UTdq/u/KVgg8Pzj6SOb6MN3fHdGrajdwQ3BSj1nc
aMMSJz83TJ/H+LWhZGzP/KchHGjS8RuALqD2h19rSEUzak/tfGOVpRQsWmo9KfRvTFYYdghl1AJs
H56zJNvsEqKzfusaCyLd3QC/OjaUXqCaNpuEZmwr0dNjZfAsQmjczHKCAdA/zAEL03Cw87/b8n97
kDqNN4f303dULYxXC8Egkg/L9D9HYetLRWf9uJu2PBvjKaP6MUy10bXa4yOivb7G49YKGlAjnoCL
045dArc6/8ydsLYR/JLBcTtQlg4rS8RPdADy7juHPu970Ei9IgdqkHxPQ0uUi6JNtKpulanSrSPy
aOuTnWE8AzGuCo1wj0hx2F/GG7Pxh9C+VjltVliRapIN0+hUbd1+CTkYaO0hg8HhUej7s9m9I8l/
jepy9ivPIQ3Ph5AaKz5Vmtp49TB/SKwnEAU2aOXtS9s0dMHuOfR47pKMjh5TRZvYUyWqlPpB/1Fb
mWvrRopde5Y8PpRQyUPVeyKf+SADz2l2K9RI/zDFEqwM92Pbnkd6RItA5iOWBMl8qC8Hca7NI/ku
d44TaxJxot2sKmku6ICSrP0kbEuYHUotEPaJkE4iKuG4muMexdlZMp0Nokje9EXG8HS565CRTKNz
otTbisFj0bzPs1D0jPEEqvzpP+448MDlxVne7qd99G+36XQwIGI+vUvMD+NnawarB7P/9CyNkMYJ
vi/NjnTZD3xBITEQSh25a69CVUOhoK57gbgIPuwh0TBG/Xw7/wXM8w+FkIDnWKlACEKEgybImTOP
bJNm0glb0Ko8O1mS0DLjlSRo8mZ239MAZ2jkT+tjDH8gcEetuvozHWg+knHW0iuB3nqWcFm3efqO
xKr56osDqNCULCl+2SEk6KQHIDAbCzliJqLl3XrE7sXAtlzCer0SaqfU2JIdT+aqxo2NCV9USMrj
bSXGHeOHSnoxGL392FRK7IO1sfNerIf8NBhuSYVwnCxcoZ9k3BSCqV1hVX28PuRKbOdfyvw7zDPl
S6mOT9pz59hEU/KyWgcYQs8pwO34+TPHEJEj4HCH+CHc8zBa7tBiKWXLQLRFonZvLhnBFDVN13x/
mkadpS9MsShLE9zo52baFU5XaaiNAddtEcnz4zFfsqLwTpcJzP8yUT0tv7AjOayS6QNrBeApsfot
xvuc/sVMxo8s8TfOOY9Z4SmcIwPRRYFsD4NwPODkWS7T+8gFySonxJjut/j7nNwU8NBYyqInSA8g
w7ZVD5x/iNX30dFbicD8uM+RviURIVA1JtLufs1KdvmTi7u8fsyOnROyxp/pFFTRZcevuO/xw91B
sco+/TsYksKg7TUXmUUAj5ZAuyB3OoQMr6WxlJQOL5HqWXQ/0/XMPmRhuTmjdo2xyWCNxMvK+zjl
nDsmGGm2Xvoj5ujd5OGjySVxlKlXxZTEPsiPPH5x4mrE3QlvME4yVkfadyo4jHTovDLV6kce57nF
TFAHjPyRzRYrXcaep2rkOzHYwUU5vUXbpNNkAWy8YNsArDC1v7igRyofZUqY+PkRpml7ZP57bvoa
4TKrHVlAP9CxuDRZdyK7afL3yXFdMQDXj4ilpv4igt87gQFxUwcv8cEIkflzf0ED9pn2sA/pIHpj
dNRdu353CAW+BItiQw5RBkzj9BuoCZPJREnv/4YduChfkQ5tR5GyNsnzwXmO7jt4dXkwI8bN9aaE
Fndw96h2oCDyW5HC4IEYdI/SU1jBq06e+CS96wl4c6ZzG9vm7npJolMeDuw9jkUdvjxv9dbtU8U7
dfCAV7eQHdE8nLaApAwLvdSPBWBGa/wQq0kYjnl8xewAcVmfOSYfBcemgQwPLbdztyL+dYJ+cCv8
nM6077sxah36EtEQiPbsCfNcFrAk9miGqQvUDXmNn1iPPqL+O8rO/aJOX+PWPBNok1z4PdEtoBf6
QwMxBWalGvEnZlHEHvlIWGW37R/aIUOUxOLIwIGpE9OvcpiLE3jmpcMjpQS+ZPshtdPz/FB1rhT+
ow3/OuMw5awBL8psI+d8rHyCWrgLZP3H+jhy1Y9C4Y5G12lC+yr6x8xwAsyAkVox9Qf7SpbeLpjX
A9CKCIXkwsyZ7DA0aadnjrZr64JKFTHUYgAFjx6XBxVWnv3yKujdNM/aP5BZAl3Xi21x4ttzk8TW
SaOUd+kZ/SlBdi24nmse5MIlOqADGKHRWUCJvxKhFFabPUi7F+JQgA1I6r/gwp/qkFWoY5s+TyGk
7KxpBMpUr6CCOT9OBHPqpBTkNNS7ipV8CqqMOHjjVuj9yZ15lAox+ipfz6JqfqiQHfNvsbHRBTN8
gd4XdXWQlhXG3crYK3M+NJCklLJdRTgNbahq3w0Q0wPhhza/UbwOYesz+art/5iNs61Yq6rlStGA
wzXSErrb7lup9Pt89JlfGSGVxo0Qb3h6XWQ8qqmBig8/pGqzPy7F9PRqQsG47WhHIX9CKTXeUW1Q
jAjreQoxMMkrwduBj3aKmiWedaXE2dSGoPKr7v8oMWotphGj2iGdJELV+cD2AFDyruH6T0Et9hBS
Aw7CgirPya8leTUgc1cAPcVXZUocI6ljreK7vJKjvj3+CTiFPrLqZjPURXX37n8F3CDdm0Pxv+Qb
jximUg5rDFJSFrlKvECyrY2PAHu2Wo7D/tf7mcdB+RRhJpCHwh8AVo+Yg7prvprC95Y9wIrkfy48
vTpAM5F/ErUddGtfiGQ1ftuDsVE7AYz+BPp4au/z7lSoSM6rC7OQ2KNr8KvF7UClD9UBkpsNHM1F
8+lnxVqko3t82QrMV9pTaXHufMZZfO/9yc4roZcUcC1je319MLr4rXqyOvC46K0LLyQ8T+P7vP57
woRMKdHU66eIMIHIdqvx262jbELoFWqCQ+s6MsPCJ35RdkgI8z4a4hOUfDLShtj8+/n6agW8Qe4F
TY7hEKDzV2dh2fVpJPogw9s259a2UBwLw2DgxhH14iZ8Rk4R4w53rdp6jtviP9OSz7qqPb/SiGpP
GaHJhvstPGVfARL927edwQyCNjRqd6eXqonHC3kD0ag7QhAWusbOpMiIVNM8Gix5xa2xFc57efhF
DNLKqm1QN/+EMr22DFuvpdYUchwONXEJjuq2DSNSMXGbRzDHxp6dcHKZuffDNzl+NRg7uRt0kNyf
B6kZ6i7IjXBoRNdbx/Umrrzk93NP4PVjPjmlCFJDaBs4RMZF1sLTxmjPnd6FuTaJh2T/rLaF4oYb
HeZ36vpqZlRxFo3EFjwos1pV5kcB5drj1KNpM3zYInpaYVQghHmnyLL+Su72zPPlULQOkXb32Obp
MFs3ZuUauzbqeo9trrZla8k+Eoz4B5snZ2m+rYfLbTryHF8hVdv3d4LbHmCLYnws++yfUI2NIogE
FQuul2Lw245fl4tBDGmw8UrOMUvroANLNDubZ55xTG9tfDgXdp4jCQgviDul8P1Z+IwF2dWU+kC8
JH5qwLRaOU+mWyp0KE2+S6OoD0pR6Sm9fbpr9MQqeqsXxSBJHmV9qlvYznl+ShBdKpSGIk9jQtCR
zZYyF4mxp1PLbid1A5RAkTMaH3OhT2zwLvJgDWWKCoqyPURB+lTVEb6rYNH5bWNxdPPHeO3IYlXX
fXDhBRCsiE+JotQEGf0UhN/o0N1xHz7D4gw+tTF6jiYuGy33ZbaM8WVIfB1sRo3TNkvi6KuzMdpC
w/DjY72MD3nQDpKgWQh3uDFMKx1T/Lzzy2Mr3ie6srwBrqq682njYeU8qd3PXcZJTEv9IPoJyoMd
pUylGAJP7WCWoeYDUTQQGU3tlGW6N6yGNpsZ7GGgHxqgJLHh2WyUl6m5OeGBkJZ17vFTNsnGyssl
1/wmOVh9Nkl+bTNyuD9bByRZDKRAidQ44TRjmyMaUMSXTyVI0ZQ7OOW0CH/sAFHWOflRNHniPrf7
Cish04DsWIN44hXU49lKEBQGsmLQW8l0asGfHAAHEb2AF2cKXf94/Dl12OVPxQVx+k3S44czKZiQ
FKflJq4JTbnxlu9LJ5FAZHDDqZyelg3iQx+N/9sWsfXQgwTnLNxNW0T3zlAQfjxstJ4vMaaMuPaE
2YEK34qZINWITuWeBULN/XQkFgs+XycxTHvC/ixjLriHSzcrwuqTxeoqIVO5sPMxc7pXa+fz63hO
Sjo+H4tq+K6lHxhYUAT2hhGA7S4FVZoW6iyCUpOBRq7auiGckWZn2RwevWZ4C3aLBaBHo8rdRc5m
XvZ85zWSKrwQv7s8L491rt+p8t4kWaIW/Os3ExZE50NamFAh6Q3R3EXaaVWPCHn3BOlraY/xxEDY
EZl8LvD3ZUEOeahUC5tH9jgKrXsRfnxJJP/cQeQe8/hX+4ScROiwu+WKXYE99otz7uGh5FRtQA1e
J5fEq2YE9PhTQPixzIxlIjDRawbZ9VaIxJzx2tV0Bahbp/EoIVedi1RLrZGfMNku2G5se6Y88OJj
V7NLGCReiqQIZhRKHpZiQ4edwofoAUZ/VvllBtsnYnXV7ksKSVCGokzNjUKgn7polsDe6U7nEKkm
dz2QNQo+xtY6CqvkLOfbYM+gCALFE1qOXADwuIiJ/469Mkp3Y+xnh3HAJI4RHtU7+amS2rfTJEyk
F40ybquvdJfVTFww7HLdE+9/WLmB2a7uuRxZEF3G9G7YcC2k3tA317+XGuZMgVVzllb1R/D8lXCS
zxAP9zHi/5/7J6RwICigM4L9yoFuRwV1vYqBEiQBB3AqO6tCMt+R1nFSyi2953KnWVcRAsKD2hHw
zbdl4R5sb3bVkpNp0FdCyh3eYnCH2cC0k3oicav+nB9H8dZR2F7+pE0O+Wwyrjn69s3VEdPhUpNH
BvZU5Z5GihzXt/yRjVUv9Lo4PVg1iyK0eSVt5a6KsgG6loLsDUnPGdME7AnkOybLsxfPb7b+sABO
lQzL6TxKRG0zlr+rfn3Fd7gkWJzqlM80rxHuSCMHVrlZtMLJRUzc09RWbvQLOF671DSc3BXyxOX7
a7bug8Z9r8grGuyvbGPipkcS/2VTpM5ug/9RNgVfUdyaLWYY+ioHTOmmOiw8VmrH1L7PjfXjigEu
xu6F+nEnbJMdTNm+QjDQpqJr2WZyyAknos5Tc3UP2KGEEtL6w2dF2svwEozt3VvudMKxydlu6Mtm
Dq7/sy5lECPmgfaJeHDwHYDT1PJikxPSgx4WMRrag13KuzwcpK+rHCiuRk+lOL7HU2erJUP3el26
xUD9fkbSyJno2YSj5p52lnNSQTZVzpomuk6ROJ5395Vfd5CPizU6lhoB8qqz3YPtcwDvTaAwDGQI
QF29UAvVUwXtzUHDDPgk/HVCTs5/DzIVQyiwp5yPdRqqMRRzOyd8Eb7UD3HBlf4ZPjYpQ/mAStUQ
m1Pix5806R2RvTG//Pmey4aGppf2uB81ztBNBCHQ6TnSK1MJcQuonKxBoFvqou9PFeS8EIwKE7bK
upP553liGIlIUKyLhFyAmK6q5QOXueo2E9vR7RaFLngfhC1OvnNtuSxBT1aajM1pRSGYaou6/YI8
+pGV+qzlZmciFmWK9kUt8ffPudz08ADD4XQBwNXbxPyMRyXLVAPWCr0dyVxrg4qwaMALkP0g/NaU
clcXFrP9koROTLbQV67q/Qx51VdGMB8qyyRslxrbImlaKVCMz9p54FehqJqwAwUb3K2z7gBsMmJK
vAglygyaIcHi709NCdN8RF44nqEJc7NWbyJd9gV++OWE3vXnh95VKkyfT2jHMPP1sBXlbvCpprlu
WVTUSJ1Ef/r6sx4zmEewfcufNIZ/JTdFYyPKvq7pcJNVOPjribKqIvDaXhwvpe7d4lPHQJfu+mO3
JvRexHlckialGxHIpSb3BJ4kXNC6CoQUi9dk8V/0V5wNZIKfYm3NNyzhd7/QOQTQ9QWV6r/Q0akb
lHoP8E+AA0i1pKhNbC00hqh+tbKrNgTF6vXtjQClSoErVVeXSvUnZZvkdtxR97sNEalQp8TTdq3j
IIhk9wfeWXGVFk49hPHhaKPmftAcL8hUeHkqLA5w53pYRImAMRQI12D5Cz6PvoZbqxswxCvk/Vcu
F2KJXZZFLNARc4QHaQN2tUpaSsLTUamjxJXGV7+qFfrLZnhy3q9DdXONz0OyOp1CZzOOjdsRp523
1XfMZZy9dnvaVKANLKuakCldYegR8GCWXiuefDIPbJeKQhab4c/xxxpgm8OiKG6xkwNCpa7uNI9Y
sSof1X1+DHEZtFVephQXHuUcgiuOpYk62sTbM+afjWZZhBPEDmT/U9sSQ6jyKIsavwqC2EGVcNpD
YO+PzKV/a/X9zsdHRabBTJ5Nc1iuBi248eqkjOQLBq7A/GhhFamIXiYdAamvSc2VvIIpn4pX/sRT
nN5zegwg7BQ6GWvykjyRXH6e1tA+tkgbVbXbEPNhs5sZIoFEyNwPqx7j4GyAJC2Wtmw/+415tv0b
3L1Lh/H32SAQDiYL+D3a+HQmfwVYwnTCI8lqPIUSYoiPPLr85lfZcp7cAXlsyWfWkhzkef6L7oKJ
xB1V/alJ5A3mZtFcyeqsFIm5Sk9B9FzhSECDlf7RHZQNOvp2mEZHWAKrGe7qcUV06xtCrrTM+qTI
241Th7K5f8gIyC3iCTVjoucmAVCLMa8QKEbDJYYmOrg0qBmk9pmJ25KbMmEiyoDJbJYygw0InFxM
/g1cxGrPQFzBIpiEMpDZx2HgJb+ZxCrASfJesBKHX9N9Gkb1jfYoVy9F9XSek6I+vAxviGCSsbWo
IFtq64SGbH89ljISnjKVA/D3+kTko2sKwToGILjroWTR3jqn6drzXSLwjT7H8TUyfuaxIr+sY+o9
WjV77elPzDTzMz1IfzdaDbU/W2F+yfJukzAfM5YJEdPkwSbSbHoyxVVT58a0ScoxIL+vl8ICGhYN
kU57VZ8tM5gqulKQqX0D/+jzoYU0wL07p3CH1r8xDf8ZMUr1l+1z+IxcxC24w5X/7aueAhYj/rmG
6VXz7/U87Hwmkc9ynTnSytzqqVjGqUqer2JMYsBLLNWPeHaIkZExV+sW5Kgr8dNNN9bTvT9KnzT0
jaJpyv8quZjEIOwHczr+bms1joOONd5YJOlyauAnLEjiZTByRgBq1lHtU73QxAe2fVNbOzLojvk/
ogXhKnbseemJ3+aWxiN10xNxIej3ed2mFdDRVBbzbSfsqNx59qPxbHWYwhuvpxbKI2TCoWs/bO60
EL3JbV5xzqr6x/tYsoh9SBTVs2OrR7/abBxyMmsXtf2bqfsxiBTORMZ/Z0sOvNql0NpOpmc2pTnB
jwCwxng/WG4acTz8dP5guqwCpfqAhAvYd8EJBQfTEBAfjVi+C2y70Jp8m4xuPE1rCV2xWRDHM7s/
0txhNff4MaNwyT0VNP7l+QSjFnoUmcTk70PrOu0G6iCVnvDZNJRloTWWDDf28jmpplUunWM9fBbq
hWP+eYXnOXRdOyDmBajW/CFKWaSkgQiDyN5GMidJ/mjnHLdduk303oVenZRjytL2qQh5KwR2HXi1
vmGvYJdO1budhzEVZDaum98pCg+0ZXlLYSVB/8N/rFMqRVGNJzwmHzqeWdgRTdQVHn9/zZCjEGeA
oMQ6zzj0ImgzjTMNH/e792/yBr94cI00EEB8eWBE36psZ+VMA4LV76g7MUtsTJgDOyZFJZzROTwU
e5Zs2Lmk7585si/J1hPVONAsZJ6sj0NugFYuvenBWIu1FL2vOrmJYEHBAMNu6NATVAQwXfAzkEnv
WxKVdGxcryHkbxy1de+jTdMu7EqXBecsGFSTHko6UdWor2af2bOl3A5OzFGAgqJQDHOc4y9I6jMH
zl+EzpNwCZphIrVI8ZxqRhNbmE+aDEZDfkRvMi6gLLHx3p1QMbEz0wk9+I81pxCkjKxR2JC6JHam
dAfBRn2xOu2wxOnD1A0pka9ZKajwOhgtsCkYWze8v/hZklpXoGsxGWZPOFB4sANZ5dTw6/p2RNEc
MzRcFTuQie6pyG5DHh+SX8YXy/BOdI6XJzWjgAy0WfxZaX/QPfoQAd7OVg7TWQbVMLbX88INgPCo
5zPuOuS4p5+7P/jqsK3sl2rNhIWnJc34D5/VF6O/9KApl7yDjwBZ1Ph6DPbJnA48vszQzQQ79oLf
0HuNTlWkloIHBVchAEQveRykkig8DELf5oFIdgrf5SUeBdDtsbLuqrhcpvk5noemTnpjyE89Bk2e
XEkYRHr2CxRBB64zm2iR2W/4DIAr5HV03Tvyh3SHf7mv/pU2+UiIY4cOgiiEcEhkcRGsGRsIg1oF
UzM08H9uY6OvCIMLgZIwM4IGY4uptRFMnPl1tZ4+rt2WYkgiUGMHCYFPsMPIEgumIgBDVu5uCik4
E+CZj+DKs7fZ0UixEmvMeC722eIp/L6JRf8YiXlwqK17GYGZCH8upoh3sGbvSX4KGJV9TnUs5ID0
O1Kd5HZ1EiyRlTpqx5m2VYfkE7BEIl8O0hgnlV3iR9kjb/Mhi6IYWH2K8XxAVdSUcN+1LSrZN8yx
+BmZRYjNBiuEfZrw9rGfWRtlYoAUk2BEM9L6XiiDa5UOm3HteOtT5bkhTlJp27wOp7YfASuPWLGE
XiJqFWvTvH/gDg5saa1XVwbHD+W1lIfvbRakeTc08y8D2srlOsQc6Eip0K8nIwapvsVaVEELgcI5
O+VbumEliNe4Oe6nW6o53z/qClmgWzGjUICKog5BFGTdsiTZh7AVF4cBqPlKURzcYqUy/oDduZVA
ff2ZBknMKB596JXSV7p/0ZeuFxz2EdY2y1ZGYC2RWGRLoDCx0meeTk4QjTVwJb76zrq4ZuBq8eUq
CD1tEMl4mXUuAuI9XNJhgrfMnBNvIC4PkqEoEvqleSDUtWESvdl1txpjG7mO9fgMfWEb6fIk8h0r
fXf7xSI8oN3+bn/AWOt2Ecvt/UQa48IOOzhDBSVfOIBhQw93Gm6bXH/ReDjoLv82Q6IvNid/5L8p
bAv4PITRGEvhhuTBXmVvYx0OyGNYCyPDXuw4cO+5v16VjilyQ0BDhESJHz1+CdBSgBr10HJpkJrE
0Pmo3CAAf18KVV3f4mWIePguhp+rL/dW06kBykJM+OdhC/ouENAM/gnSLZOn3YP+iu4o4gqKe+Hw
xh/ywNM7CpZU+HWRxPVggIvnpk13XIOEGgaMYcDLq2ymus9myrbQHvnK91nVvQykiA5OV+uHKiMQ
SxFDhX6mIaV+I/yer0GM8Mcn26BdlBCDPvT2gNrU2PZOmqj3BUpDUv/axSEZdxP8PWBqbfG2C9EG
ITXIp/3xR/+aF+bPdFC7hkcA1t09Y8lPa8QC3Q44/3oVU/VQN6yE5Debz48118tZNvhmYsVqIYy7
8wmQUUlTVsVOaiRNnajOUJtxcb/CeoaudB1b4S3s9ygBBOY3Q2SkGlHcRMJgdGSjptpH0nJaKi1E
51kQxmIY4ey6sF4zcDnyT/lYGBvraRKCsv5tE6je5GsDFqZo4JQl8l3aMA2Y/Gaxi7nK1jXfmof4
b2qlfXDIDm4L01Xl2nWM/i9NADmGiTximS57EjBZ8n4jftg0nPUtk666cgvSFHiUwYx4z9SfUCQn
0aF142aE3Lq+t//E+KKoU9qHO8F/8+FYkJEb1trylTBLW5Bc/aF4FixA/JXSLphBoKtqjgTaGoXo
+Rs+JbAR5IS4ecBIuXt948dvnsn3dXoRdD3zI+wmp/phqwM9Pzwrpg1nbQoTu87qj99ivxIbIWv+
DG8cra8y/yxVBscsSXVCsDsU9Z9oXS/vKa9/ToBfIwFx2sVnVmSw+KFvX1trP/1u78szSBhPFxH2
BLb1cZH7gA9111ir2a311g5Ry0Iemms6kSBWJsOuDaWQzfV5yyaw7s99JCOP+XjUtz9IfotUY8UG
5P3Nz5SruZYh5ZeeVPHBXNDIz7LhG7tLGKj5uZEIOUWpEEmWdi4E2XXiacGbf1Peo4yngs2Bke6v
S0VQ+sVT5AeMv9cievE7OkWMBxnszR8ax2woI+JLZUTjiOpsf882dqjqHJZibhvTh3Q8KIkXmfK9
AuWdW7fd79ZK3M6sSsabkIr3pbLWf4ErVDXfWCLVz6ftBCVnhosjWVwoMiUVuiL+2ZfrWolWWZqD
YRxrF1PPb3AaUex4u8sGeoNtgO21KGjrZ/rAUzQCtA9TKFlY87EZ4mO8nZ8c2DxlQLHIGMIyY6h5
zf0hYzG3IAhRPhhWMymRMkbuQBQZSgr5skZLlnRGLUCe524jGg2Rfdp1fdSfH4BvfJ1y9xjt/qpu
AVCb93+WD0+gQzil5H+UbiG1mW4YKxnvLIPXONlZIZ+H87bNJmTUWs1ew4Q56nRLOfdbXNvW9IiY
HCW3FuyMSCf36QNiuPVmbqqGxIaz7vMoyOr+ClK4KGFh0bTH15Zh7uWR7KU5Tm0EyJQEG6prEZpJ
f6lDgVFuTfMAgmYwHeRXLPdna9PzOYpQdRDryBNLY30kZ2Emnftyq80FRRjF5WikdQ+Eh/YPGpWV
Kq9dfxQ6IhKdv/uk/XjPf5PS59wVALhXN2y6dPvEv21XEIlSxISk+WoGYQ2D2tl+8+LKvZbREFLo
5TLibmIjMTliR5TG+fwY8j+sq1xVPOkGSKfLblsS3Iq8gFCQYAxsxGYKbQSPUPcbs7sq0NsrD0UN
Ezi83B176x/n1suahL/8VfK8ni5j6K2MUVyIWz3RI9W46QLGnHqmpHr5io88eNEf7iwb5uP1zNjl
v9s2LAPpajYhVh8XOn/aiF5hqS09rVV3/BPGsKVd7Y5JZgmFT4E/kO245ZdyLb27+SVwpP1sO6UI
G3yRst9iER7tXKdrUJiLlZziBknWDmZfeU7xypgOl+Bz68PFRWtnNqSsZEw2L/F+/sTOilBbKvI3
pm3uiQKqAFfKW7QSQsbB5c6hGvVDbKE292KdofgaB3pPrt10ddLxC/OLWW/DN/CaMAjWvDYx6LDs
peVv0/4J+ADDDK4UBhJarrvnESwzYAMieYJGbf8BIvBig4xYD4nQ2gsAmyVihnQM5Fh8+TMwB+5Z
HQZgAabYIlyDbJUXtlPIJYfzYeAGhoq3Sy24D1+KOtNq6ErDTp833LvQkxELbB+VEevAlrMP4e94
fVj3aZQI2qd3KeDWor62jSJfhj5OD7X3rODp50pqGhJ3efnKLh1TwN9vZiq2gU01CFbGZl9+cEi1
dT/r/MsG2FBE0wTIjebxTvVlLllGXeqbV0Pe472za6l4USrSEUT1+H4/HUD2rw0woF9e3cUaDPTf
KODqHt22z5g0JOG/z3A8q5hYC+VjSTEpYlxQdDiNvVsUuSlemSyR7fDew4MW+dX7aVV4BKr/R+WB
T6P8CBWVXgdC0JpOkHUjYFGczKgbQFGMomEQsn+XsIoKOnBkdmYbieTOIeBRFGxFqcGJ8okZ2gFU
pJErzLnAYSnXmZwmUzMqLjdPeiGcUnSnEXEO7s+9PoxhJlanJgeCK9yAqCujYz3eby22Z5vJsX5G
yVsUVQRyiyVonlAVjdxKAl8jhNiu1uGnjyAmv+p1Vw96SaWzV5ztgXKmtT7TSnTZsNfHvqTFI45C
PDP57mXs8BYLQVAfp3zpejj+HQs973d1xbYh0/2I2vhsghx5V2zWH37g0b1UYEc0miSgOGZDUMUr
yl/s4NB0EpWNtPYINOWZBgCtlTbxf2smE46zI+pT2XOwUu0ZlD13dTDoJ0TkSGOgcp8VoQ1ALoW8
U4K2KWie8TJIOjAs1QZ5T/dvrMq7emMq//k6yzzqW+SIgeuQznVmQPfubPtfuQ3JPg4Jz/yqOx5C
S2fi9/3fdGlEFEkxUNzH0Z4qeuHndfAL1BowwLjsWyRDFdeui8PBTH9P7e3VD+PxoENjCgmqUJiS
t9FNmUAWxX2qP77kK817hYTjUwzZFfmPoLUEkMKyQl5fUdDXBWG9hdHgegvwCVkBpQVR6WnDpPyY
z6w/THHoB28pk/PlbZwSqG3m5DZLI1dyqjKpXyV9/1uyc0vMXsTdDstG3CpUGz60pDrVtA2srACj
mVwoZClHRLNSQNl4kgY2Ofk3cZ50VpvPLhWkjR607yVjqn4Y401HzcvCpPM3GRn6DYn4dknbGxKi
fNRHGT024WHjDp62IFpf2c2r715BphIZmdl0CZcP4Fau7ZwQTTVkoV3tVuboR0IRaOhQxctDZam0
bKnzF8846KC4PgOoinYqzkPSXuX9r+iJyslC3kYZdham8gp93BzwShL1nwHrN1xCTxuAyIfzDMWI
BsX730B1QMEwgEKHxmDncwHKU/VfdmYgiE5XZZqgSEW+DiVn9Zwyi+IwFt4fmzgk5e6Vkq2tZwp3
WlNpKkLSzE+Odkk6DPd+lnwh/JvfIgQe7PKzJhGQtyDYQoxwHVMwExkNPHQdHpm7TQjIUqNlZ7CW
z3U1/CwsRCnLqyVIPoXYDbR1HQ+/TfJ4r1SJahLRaRZSmb5szRivxRcwQT1YZEFE/4ocEKj5I4gV
rv0nGycktfda+PU1nMrG/QxlkQqyBJYYHjapsK9rzQ+o8gLqdV4LzxfLiNKwupmSO8IipmGzo8/W
Jsw6vDLIu+ywwhuAOUdLZ+QVw0Eq+5RXFVPaqCN64BaUWlsABtnr/mSuqMviR6ewnGcfSA2OqQCK
KPPpbR8aoWbUgmN0fu2OG34aE91G9+5NUYo2RAnDo20O/lI8JAPx2y0or9+P9qsPu96dPG/2V0ok
f5AjKFXXob4AuuNyE2q51iOVZ73i23VGPiYGT2SXECiquW4PpOUraSueT/NVfe4p20JTUaKdp+sd
+Ks2BIexMbCDD85zNj4sXLrJwnvlvOmyTXA0QYEjSt9RsLHrxOOdi8ulDZEH2C15EXNnJNfPkJeG
9qh+fUx+xY2lytkGXnW5Gov0qiqa+W+TP6YfEu/n6yZ7jQaZZbtYUJ+j+LY9KhItfRU2ljbbnc6l
YxbJGPxSlGV2CcullPVEyMmbYmaggGWuR2n3Fb9uIxcnuGlDQMEnI/aA7N+/eTHbfHygpwQknWpI
4bolYeJRoRm2rliNH6xfC0KNYemsmU1eTpkf+9o/LKkgvyM2hHt/CRQn+h9vC88LYiTtj5fPJYoU
neB1trJI20kEtyBSTpoI76JwyY17Sw5/B6QeBllIg8T0EAuS5vxWlEj9WkKCnmCFaDeUNTz4xbk+
mmZgp4dkBbXCV5dHlh/ZxOHmtIE80GdOpg6rgnUik5oV2LfNOeLPx3G0HC3zs5gL/pUjGlUDD9UX
qz/ANz5ECdQzKOelBV8p1juIms4lC6BLJXPwAP1nRkT5UQ0tapSkKOehuvK4aS5S77eVFO1KEx11
rJEGrqQv4600jhJoldKD5Qmc6s5PSZzZ6ZziWGrZGxO1ywps0erLC4jT4eQwZFSM3FbopQOih1NP
HUyJ08aUD1Uam1Imhsot4LeZSIoIHLt+e4AGYeNwLE1pr0Lwh1W6jOnOgvO0tjIuW5Xh6j8yUGfC
1rIh7WtW3M8MYfrS9KMxbzJFV7YWoMdOfrcTenkeCMdR4/BpdmakPcPaaOjuFum/HXXGgypeBdni
vrXuHYHVIfP2lEjb/sd6oHrYS2q1WW1NYWYJCL7aapgvGEhDfUrp8wu377dFh4Wo6kkrz373qEKv
lJs+y6hP6tKLFaXtTVd+drZXBDEayyON07OTRKJU143qr80Bdph2U9awKt7yKdoRrMNTjvqfRMxp
9hGwnjFXPDDXuuX2DRceCgqcWJc4TQrstkeHDBVdjTfLBiucB/9liMkWuxStl8d6GPZTu+wvUz6C
k3aNA6q7Unmim+DiAJfZnXFHM2NHT6Pgm/2LfNJc2uNoC3D9VLIgRM5uIzXOC1dZCmob+TtzS7TJ
t35Xgk562sonZmtlUo24axqvgrluSZVQaX1WS9hGEU/L4nhKNRKOb+kxVs1I//NvqMvrfqSyfyKC
BSPp6glH+5iS8YSZ5xR1LOuCz7P7zSL58ET5ymfCTmJQ2CS0S9Or8f0lZbe1CZ3llMoID75jZMBn
mX1ABrvZp32ubKV8h1H64gy5J2hqEW52HwvdChVenDgduNTFRHMuZK1Ciji4Z1pw+2yOSoawu0PI
c0Kzdg8jk50WCtSkcYadPMKmv8WW6bcod9GN5e5k886rwlWpzuomtVjNAp4XZMIZFCakAd6C4KSk
wCs4WSqKzaVzIRn7t6AA8PNdkBtK4gYEl6xwselKuqF3zc3QC/wx35miZuZ1iiVcRHIjkLLIvX8I
Z11Ppz8XWl2YYR6am91ffCj0YCklh2RFA/+uHmN1XtbRVFQeiapJd88Tyh9uHNWtcj5Fel55QZdV
99hMv5bdLgjKcCtSFarmDzTTuT4BPkj7h/SCBePQmx/fgkiHRrqH69jEwNt52Qyt5YD6ljz14/iD
HlNyf3Isuxa1c6yb4irfTrbYLtxAh2v3glATsZ5LGYixlMIL+KyhhYlRZ5hq6MW/A206Dzm6kGB5
oF/9A3jid6TPmlsTQDN1T+p6pkhf2IC6EMO06fNiIMzvqLbs+lwBnmNxFrGhVTqOIHiOp/0RR0s+
Cz1vQ6YOI/iNDygANhIC4M2l3DEQG1fPPtxaO+LynUhhMguVNqIaxggraswNO+CfubS2EvuJNS7d
a3acjYFGvSN0nv9/F3xzGo4ZEj1KXvFtQKXf8J5dX+ohpXHX8mz7W/qcXquqQlY1zPEqBDktxpCF
sdUQgLcOBjPva5iFHPXPxl1uOcUNrw4SQ8pVgHgmmi6pouJM1359nWTr8rlLzBx+1FI9J82nhXQC
DHEiGNuuwNX0LygdMO+pilqfjPMxOiavCSmIaK+MGO+ZMqvh2wKhKTnMNDagCnGkQE/BpwiP5aEm
TxwZkPSJSUAlcMYi4m+IevsaUVOiJJxDwuWIXpQYlV7BxzcOHqJn1njUuaoU211lCAIg6e8PW2cc
4d5/DthR1W2dTc50KQJVePsQhSHZulqawNGMsjgpiVJAQkXpygcEfoVNfa/E1tmWCsUd5qZejVRz
C0UgQOBH18FRdaqQxIN5JOqMFHOD9CVfJ2JjEBKGT3qXYSgH2Q00YW+L8agDMhFLblLAw2EHCJt4
1T1LrrIEz5nPzw8/rMAq95XUZPHf4pXjdSx6DO41u4SAnMCpzHIWkkP8PNu6PrlHJbf8EpmfKrix
6pzbkhmPIDeNfJoIVSNeF888yLmtXEsqYIMSccsiKelIQXUW6HwmMkGcrMc35h6g+HVLvjNp7NVT
NFwR0nNnQ5aTN/q0Qbj0aQRyVh3XS93eOwfXqVJ/lh7rPGD7A4t7HAQoWfid9oUR8UH522+qlEbM
RZsR60+pnaVwzGbxnKF85CppPhut5zsYzzx5B19lYDBtgWwK91DTI/9WEOcnXlW/8gqxIIB8jWnJ
Y2TDTKetxwFt+qkOiFnkG8C0VSX8TfJ9AGVmbIyOB/pETJuaMZj5Zc3+H2aGTRiF2+TBD/JpKa1E
Y6HVN7In+GG3c9Wc9ud+dM1/7YLOhqjR9+O1m9XBp6pYnXAxC6LJFa8ud1u4ZXLqPuCMZc5Maxl0
u6zQbRZF4/UqQG714oK1WB3n1ayA8KsvmE6TlQ38TviapTJV/FSKYJpubWpehrMn/bRswO63eYxD
3eucp0e3cQ+jDWmM58JIYsNQgDXbvkmNg9nVH8SGQGZL2eU5b+vHE13roTgx1/roTGdkW6mQRRfo
S6qtT07E4FHB0Hs7af6alaGsd5/Kbh6rRVxqzmJeuYDT+rXAT2ZkR9TGY+BfBvO5hGOIf3BsoRLh
aYcOKEgSqAMIRrAy+aCbZyKsU29ZBUJvjGmN/yGCj828rfpjVkRH00MnT8hkqhNNC7FyGTBXr91S
u4PhkKZY4TFR/NKqdRI+ggL+7mQSaqRD139V/e08NYN8Ynl5aWDTRMQrOazWaZCJVAtYoWCY9JlJ
JrRRdnh8sU03uz9EaKoYF2IOSyzJrBpO9li4BY+JZLnpdRWwOPgA7JPVneS7Y4B4nouM1VINFiaH
wpMYRjRnxsaFpvX24FQ1Hlfp8hNCa8s4J9MhlIvoHYyFdbubztTxNeukys+z4he1R7ivRXK/75oP
7kmxkuQiGA8SkUx/FUrqGj6wgYq4vwDJe9sElJyyif4hNsCzWR33d/s+ZGOc2cWKs3iBRW4oY4xo
clkN29MgTkOe74eV5byid6ipkJd3cHfOSnGLcHQ3fOHG8P+euldHP9ahKwD/YEe6j5PdzEgI9yxX
r2fRWYDsVuKoATN3yXjFJndd1I0jWgrzjPODNs6TvML5sQjCKutuka/0xj5a/0pE+2Q6LKzVhqYI
VSqxGC3r3cdru+/p7h0Yy1eQ3mnrYiTlD204g6jCE6BHnW8r28ttdD2uhV38M2lBr+tc5HnxKNzB
VxFUeO7GIS3tLA1A8KbjeB+y7pzl0cEWoN0jBVwk6nCHGqe5/OLe4ZD/lUWXs1yak4LsKD/eUSst
PLgw9ejm7H2F53xTHjXNirU+2oBlz3O0VNlAZmz3zmCRfVhkGj36KErPpgP4O16/I4wHjzgkxJWj
YrgzyCNkUgVifPZ9VbqSuOwbsCBni4uj2I/hhNi2xk+cA7IrnQ3Jl2FZD+RqiX0sONZ49b+lVfgk
R4+npxAlYukwDQx5RDTxRrs/enWQcAkyTvQcCK7P8lPYyGzqqq+o1+I6Eps4KvMuyy6qeW+0xlrH
auaKX6kNknbBrioD/o5F+DmEa8h+Em2kXyJJn+Ikd+3P81G+4zph+Ofiwc5XK02Pzv3ofQSlkyQt
Vhm5z8GYXqwcAdGVUibWzcu4py//OvlJV4vipz0Z80Gm1hWtGHYblqFNYAsZOQOLpwHRxwa59V7f
IhHs1cogSFejidTU4A6iPJo4me/rsXavEa49597N0N+z36mwhR3pOmhgYQKPGVZKU/vDqKbUZMQf
EF8yfGWwfw1xM4RZBqTcLK6VKwkuKTs/RrqsU3mG6te13vO/JYPRqvZHUDzUImyXxyDYO6mNrn+L
tJKZH008SdK1T57m5Xt2CWKsZFQ4Q/YS6W+whIvrwou+9dqyYr9GX8kP5olJwuq6IPc/vwTUa5pe
mhkj6D5305cyess7Q6z5C0aF03zy/OxbiBGqGybmYF0VTohpZoyjx9jFffRljU2/yT7I0PVl94FB
UZqd9zGCLnGZvIrgXhGibwIuU8vSV474Dr1P3AhamTue0GdEFzzQSqSgCrJ3z0GL+rL2xY15AO7Z
WgXsnc+V4QIV4FXdFoYZdN8e7OqsnxGQvNJc5zI43NN0wtUKeSXVAgdbi+J8THmeInFVd2kKzLZw
2Az6XMPPr38+wnLV19D/4c2m+233lKxDIMKlrN+s6AVcYx02vVUAhciGwJqnsu7kzOFsMu5pfwRR
UNWVPKUXn8j6GNhLbPlya7nfrlNA9voXyPfVZX5Wv9YY4eQ76nENcOvc0sXPfKtfLXjLgo3v06oE
g3PP08hpP0yBsQkiKLf6VRABoxQsAxPbAEMIlroFjqLlz9NOMnIDx59j9VDLkPrxNj1EXdeTErK0
WNxtbU6MzNFxNKDa86JTruDKqekh9LwNMx/LFuF3UGuGbDdBJUCjnYDICdgT5LdMBEeP/EyiIgkv
e1MogmyiO2qBjurCkqsi2uTQ/8o2KrE6bCs/TQ+gTLI3cVhvMx0STkwkIaVG4xr8+yAoBKzjF+rx
JltGmkh4iGU5ufDyUtbytozGDXniWUleZlKOTtvTuUQj9+VgbOSXsui4I3qox+eEwH+eH53G1wzm
y+rIumB+HEn50qr4Km8jq8s3PcMR1shmrUERmYoESKeGLOOScKrWBXSJR73ZuqmhTZsQYZb3fqkl
Dv/wnqan+qBJ0cnTRQv4M4Qu+NX8AeZ/cc4I5xPAaGAlT7okFaeHOY6GLz2kFjnJ+EC7Qx2bup2Z
l7RmdGfbaLjA3CaL6UAGsIYNZToLYTclaqU27GFmNI4xA47TZ5YrA7gMtVQ9duU4Jjv4kNF3/uc6
vTQL0Mipa8tx7sYihQO8CU240SsxLZYvPqea2Kzo87dH9QDPc1wCLH4OzR2nBoU6ahXz2naXJf85
LLqgDEBlU3NzUR0tIEOC0tpB1NyIz8995Cu69rQ10zJpRMVRxHCwDfxX5BFp/M/SOD/Bbdc3FmiB
TvfBdVf58XRlhCejJMxgudCU0qkLMGQiHtKopbDV5T/3Y6lm2j5DVXiYCLv1f4oF4eU3zh2rSooP
9lvemcpQWX4hLUYMWw916DTSIMTfju6mgQczr5Q5it+9/x8R0JOlrkZigsXjtPZz3N2QeJ102/wC
bucYZoorMikbMZ9KzRS24EVuJlF3nyF6F4Wx3h3lj7eLGvzklaLhPTvyLWRweW5aKvZ/ebZ7qcz4
ZW/KxV8HZf9HcgxWTd+YDcDsGIWkP7FKT2vCvbJB9VW158o56miUPwSDMJpkyzOsvUtAqodIRX//
g5aGHTxqgSjsfLNMv60u5dom0OzDFW4lVzCL7I0/KgUoYkdXdaGSGODUuBxxyPjUlHua5bWX46Fn
uZYRxavUH+BdwqdTLdfh+6PtDwXsShFRrsa9O5osg+GdmTDnJii0sZKCu25B88+R6jkmZj7ytoYJ
6RaDTYRx5iyDqehfiRMQriE1iwvmX4TgyUmY/mkwpzMss2iTpldIf0CfVxXDJ6hGC7UUexRLYFP1
7D+/taRVE9oWng9vRxhD+n5VKNI/yShXWWVt3gMtWG3ptUYilkwlC7R+xkscoXH2xZfEHC69donC
htlqaQPMRKLAs670+9QMYZr77jrdrJJ3c0GIVpxnkzHXXk3jKwC1KbR0FoaN+maHiOM+oenPi3mx
Tjt6Yj/JCQgHoH6aH+2VEASJnAO8AkCIsQ8NcqK25ifG/XtpgmzmyKGbdBAUmnuvgShJC0UsSQ7s
spXlLQWs+N9KZJ6n9DuD+SW5foQEVlzSWI08tMC+83rQvm73Uhg6/D6e9gwS0QbIKSfuXvRPPnNL
2H7FQ7R97tNPdosMCHoMbRR3q0Fdr/BCghz2JHDfEVxPufldrVtjGNrsf14R3ZAD/bZZU41JFq1q
kTIgRcrkqo11ZDWjpNYDajejPsk7cx/i50H7v1HmH7W1zk8kaLI6+/h9COj7NTcGpVxrCBQ3eSgh
qUOJqR9VuXQBjKxxFyTSQ3BkE3mHG0c+VkuQTB6GTALQwBAOuYZfiByLewlVKU3cLSZ8GwfvryBf
I+6jZzJSykBi6muW2V2mguVTTutvofYngLJiZK2zrTwZnrqqhwgEeQno8/6z+FgMgrzV3VJlszAa
YOYIENsHrh+4DYPLsk86SnSGrSYHkf3KOfI0o1uktwJsMqHa6HcWr9ONQF4hSOypy0jGcmPYz3dU
TAh3OWscrAD5TssVTuiQL2H9tBXqkrm+MxWLH1Hs3h3U6agDRFz//gsFMwyTmuZu/zdnhpRExojZ
tiHU9FHYOW9lze5uVnJGR9ziebftqy0Zqt7/uzQTGxrYtNfcu0n6151cqbLkVwgs5SRkvUBDTdXp
NFMiHuljnh18o8PVtH0o8SZgWRh5klky6pzEUzsgVJyRCituPq3yd/bcgH4FSBwA2lEzuGHHQ5L0
k4MzD040ZCUSg3wYFgoiCIxtiSCnm0oqLxI+lg0DuHBoVTcBxIT6qyGn84sHvEv90h5yuDk3NLUP
tr2KUs9OHI1v05pGfASBoTDGokp7GD+S7LfK80ODdaLLjaRaih27B3Dz3XSVxsSAUGMmkIjJJ+O7
lDrPfco4wZFXvY/t1mekMoxPwDw8I3JF0bF+0l86QGIh1l1BqxkiJFKi2SxYelIJvaK+lh5cQbj7
g4d2+rTnnYQK5kV8LTAMT6d56aWH8/iP0EEiUgNnulpmy93asjQsncBFcPI2uj4vDVlu/lUQnHNt
VUk+LM/ea1am5BY0ZpUVmpkj0CcA7DdP2/ZmCmPQ5PmO2tboL2C0EbE47jw/BZgNFtwAFx7Lof2Z
ENRRxIi7xNE/Xw3e5kDtPwO/VAn7D07kty7Pm1aIq2em+6ayNh+S7x4SLA0y4AWgzCy5Ni27HcRM
QpMPtpywfx0/MgWqEhM4mqs0zgeQCQqJBA8N4cJgIbbLF1k+L0NWmpHpxGS5y3aqrNhboohf+GcI
W1jX94w8aV4o+xYKhr/dn6O053Qmp6uujPWY8V4yUymJpp50gmN0WKEQiy7++SQoBNt6DBHbRQmP
hEcjV2d+3ixmOQU9ubRxcwthwvjlwLkdRtTNCPTlfJau0ja2FEG4bWOjmYbEV7oc1e0JTbwvpXeC
OGXPqSLNOagryZ+6sLxF+8C+6uYqfnqPq+uQTmGVphFrsv9QfXBU6/Cun32dNRsilcTqwK5GIjN5
EVQxXUcAJQ5JEFilMR8dbFk7JrO4D+LTXDaUxoNlYB1UeZNrzqoP+K6C9EF8l+l007v8A0WiXYUL
9MVtU/zGYV2/r4mN/uEtnEcw3zO3+Ety8OPPRXE/Ul24ZoUCMcqfv722WB20JL+GTO/dpar87XRd
EUEzcW1fz6GeJX2y/ahsr6SJ2DcexhGsuLxfzAGbPwhyNe0s7AgOqVHk9I3AR4XkQrlcosMpfwMC
VoKT5l9UoyxF5aVqYC1ryeNLy9RUS+LMXS+EAT36PY1jfiNb+P5RMKE3NYA8iokx7pcSER16sRlX
it4wR3Pgk/crubMcrCORn0735uiMGwNDRgj/IXqtor4qfMLkyWAWltCZ4oEO6BbPVNNz7LeyZ7ZD
WqPHKpqoqcLccw1yGzVxjspDaLaX+SFaxxANuxG1TQYzwMiqXXclzyZ+E3nyE6/bb3uZ+egw5Hk6
ojhi0syKpBcQiak/a5+JEj+ret+BCbH3YjTOp/SBii0HP1LrRGGhiCyqXVZ1HkRQZhoyORQAoIo0
EX/ZLhqrJ9ecJpTIE5QjaSGISIUfjCVUv/vtrQYlckBsvKPOqm22/pIRvLaqO2odTd6QOPoG0Cxr
1ylVSGSj16fSYcTp9w0hQmcdTcgKD6mgIyXedIvCTCbRQywzAAqdUc0vSFEoTGUms40Zqpn7IOBb
VPcPsOSKE/Lxrc6Kn+XA64kjbw4L3+qHBpptjxBH44RfUTawlqKrK+5p4rDOYQ2jy9H3qIRW5iAN
LzrGlzVs0nEvWnDtHyvZgOFaKOLdvRpu1nGrqT7a0+NezVE+gvIyrNqHwCNRBHovMdADH6sD2VDP
NJZdkayRYg1EvDxoupSewF9rd3gel0ntgPbm0EpMSbS7omtdBhKONihNeQtUHHwURvOTqayW6lsV
UwbdvnNTt8Wu3/NPIY5uNjYQjORl0ZdIWx16dttKHDUVRoMO3nIfRp6eP1RkwxJyHGuAlJQ+6cXM
ox9fxr+9CePnr5PtVoUED0ZMcIRPqbNS8LHxiBxSv5M/azFFfoPPhDaXVz7zNTSAhjoz6LSwuriN
FCclcejc7SMTSoMFawQ6Gk4pAq8xhL9PvQApMnZtiJJnbTZzefqu3cEKazlcFtiFyKHU3n2gFGwm
pu7eOmoUeBmOUlFLiwub1oOOVfUsl/VbL8YcLbXOvIRpyK6zyMSif2pTWWpOEmm5i0eBWfRmLFQ0
6NYrsmWb4ElGEdHhSF6Q63Y1HhgZGxmcVKtiCmPmz4YF/mAXSUdb1uxHEmjglUf3qIrXK5h5eM+f
r82ojb7Q7LqpqUSC3TmL+UrIsRLALXbCoOXsolXYNPa637vVWJXnXUpsXW0h1dy2YdZw1Zao9naH
sg/gkzonXFUIrxbafkIdzZUleTS1Vq9KRax+uQxhafzvJvlrWSHdAjfKzsxgBCnD7Gr+WG1a/fW8
jm+8kD5tovAOHSjuoPvW7jWDFxpK4djPJW0Ex7XbzA3lyIIqDDFv+6hfcx8HgzNcK8SGdYMIeALi
XRIiP4MDLKhy8x/B7+mf/7+w4E0w1XRjx8yrR9AvGDxyYRM8Es/fi21f/QQI3EQRFP8VBbfEJD7T
quHdYhO2c+SfkOZeYF7P8qzcdKrdSLn4RMjXO95Uzyj5ImVMfCwxmVFVfgjMiepdBG9KZ9vsYH2q
b/UYPbcIbfdDm5XOMHgVfVN7QAEj02TOzo04ZGBnifWA4mTMiMNB/n3oydj9vXtLs0KbA82kI1/T
/RhO9EWWdiM33voO8A5NqSpL4t3tj2FfezV43naXobdce66OiZ66q7JE2THpyIIZBNfnZPoDUtZ3
oIWFdI7WzIURRuMxfZNIQUtcIPj78PilQ6CEquthZ7WZ390BFEM/+zT+ZqCBZVZiWtgcvlhBCdhD
JJc2gz4P/cdskTTBMECnIZo/jMjxtr1v0sAt9IVAMPM+gV/Lpw/heQLPYDqWqvFPVzL8PKdrhhEi
582wmpCCQzW53DRrORhPX+P0QMAaXp/mwtrzn1lt0Js6DXRMXMScZ26K8ExpOzq3slbnSJmoM1xh
5WGZRL8OtzHlwpjkkO1GKcPHohSRBQLI7WtRF8xcSZss0ndGMNGPQdlwHnBtXlFztxIlvfjwAdQN
Rt8qcNQc1FvkrArRcFkrZxOK4Mk4oL90dN6tvf1IVRJmxWmdQIcJ/iAqEcmpa/WEEUCW0GTfO97V
O9agCRAKRfV/Z9mMOxI/ts0kGMwNISXbpaNk6eFg6P7gq48SN1FhlaGj7Lnkxic3L7JT8mDT7Ro2
4LEnZLCXLDsnsrQTjhxsrTsI6T2qnrWSIgcMe/noyaXBtULvnPaOE9PK0WZF07DyMgoYG6vJZ14x
4N5awItGuH94vDmNx96iQnFYDXskxqrmviF+5zdilvGZUpNOa+p4H6a8BtJJBddguwVvSq1hqqef
Yai3kULYu7q5ZGOvFM+i9c6/IutSVKYa1yGsS0nFI4/G0tmORUoFInWaXzhZPTphHDeDReOiskqW
ClipkILGdo0BKmIuGBj/SVjcS6yS2yZzo5VFBGxH2AZwphCavQYELDeV+pNpeBHwOf0yshMGJHcd
+TMD6p16mszwq1TfWKr1ROF2IUW5HDqV982kpQJfN0XppGmVCN6pHGo4iwVv6Fuin/DOPDt67KQB
pWKKNONbEoXwD7g50E1UwhfS5BVGS/jWKGHJSN77HW9KCKqoyskkcoadH2uybulnQFYRT5ZGG/g+
j4UhlfMzz029wAUWe7lGUOYfeoYd4RDz44uaBm87WJ/y0BJ5OkeJ+zzFyoXT8/UXhcnYScGIMPf4
FLkLtXwtk6uX9oObEKjdaCdPqrk4/W7wruvAc1owbes4P/h3X0/3APBD6G+ZvntSgAnZFb/oSyKY
SUUUPdmKXowzsgiW0GdBTykWs7JRQmNyzm6kt9/2NI436y3oieR16azyAA58eToz5pyFhgXc0wDs
UlB1YByLKiEsic+t4n7GhkHfhrBSXp5qrj5GijjfHy17qwZWJEJGHI26OQ3hBaAukHdW+i5XeVgG
9GVm/UdsGGsWKSqXUl6+lGg4mbs9PsiPSOMYQ13rRltjpZc+tKf6xp1ThwBYqEDxTaAVhGY020Mz
Y+zgPetxx+o8GfXR7DZLrgjbfniK292FWA9SOrxJHjFmentzXxcn/xbdo7ZgXCCvb9BWG2dJxfjI
c7CEbkMt8NHETxm8GPkPIrAVI6FuqWKSR91Pglt4Q80q9Vos/vIB0L+w3hGhq9z7GOy8AoNcpk9u
weMbHzLtrpfmpO4FyvZSEK1ZfBZOfYKCSzVKfd8jEdDz6KWV78w8ncLtNOhLuBEzZhYzZkGomUjW
eeUbos90e40MjbkdVYt7egG/tRF+ng1wwxF8+IaGWx7CLRZ8bUyZlao++b9eFQioJylgyUAWecMv
50k6HCespdPESIS7AItGKoidtujcYOnYXSlzHJA/8gJaIuEwX2LLX5J2HuMFUM84RvUGTXEmNg28
TM+8FMjXrRXz5XfJh0mUIyHCOQ0FTnALumuxdGnU7Ov+a6YtRExlNPKpVSul2ZsEuD4UBhdBX4Dr
E/1NGmbTD1QVtzDOFoRExXLcoVAhgHiTUNa+LAd4P8TuQS+5MGeTPbl5Hr5k2yQUVblX//e+h2dv
XzwrnYxetqvtU0EYmqInpVeStgbYED1e+OXS45bf+uyllKCc8ap2GK3pSFtz+pki3pEIXj4MHIBM
q+YlCIKYDoKWE9SUQyJkfTtCygsBnOXiDbwkK2ZjRoHE6uFO4Vu6k7i8olVa7/PtuHaGelOg09lK
Eniy2bkgJ70XpUXSdhSf9ZrDrGDVJ7K9giJgOs/7QMF8joMncxpzEeXmI8KdztphV587Vb5jGXlw
KZON+FVseXburxJ3N+4FAtOjw7AVUjlP831qm5+PJ61C5M0rjzimVAXIn7jiFaoaSltDd/ZhNRqG
RXa7LSFQ/dunrQcp6A06+Xmj4IfAuGqBSPOa4gUuIsdq/8PtIDZ9dXSnqNTVz4KnHHPNU2WVVt1Z
14L4ob2c95MaKh1tT0L7hwhsYklheFsG4vEyvBvdaXmIvalixfkRqfo2wnAMlkyw7OgtwPl86RSW
+wTFglOWsuuIrUdeWgwm+bgHDuboGk1pRI/7+AqCA2LdYeWw5EwVnb8E39d8fYQ0cpH3FYLUPvcJ
nA/cHWjyjNzH5mydSRmhE/Zu7+mXjiQl5gzxNSKJaE+RPOYAvDAg74a2sMyhg4Eq1HfOVU/MMxIQ
0pIO9UoyYgy1JSP4PgiHqBXpnq56hvIlpPBFCLM62wTsBhlccN/0LuOgKI3u5Wh6wFo+y69UuMPT
DnEwD/ihxdzNMMQhVPZ5MHOy2GJvUGFZY0NgM3RDr02/p00jH3QD+6QOTinEEvAXGtajyBENR2ih
UTv+gXFDn13XIT5CthR2iXGDdv5hFXp4z98RO0zg+iDYnjlVJMqMe4KXJu6QWxaWJdvI3UUASftk
VvQ93Kh97D+S2WHmlPHWNNVE1VAi40AgZyVnaavurHUaX9lp+Y9MTr9fFB86ZbPqkrGd1h3k0lv1
AyXR7+mykjkqq4IarcvewQlK6sbb75SEDEJlmFu6PHaraXygVpNYU/lx/8/FtSYOlnlCklWXzo2o
1z77TXnZr+t90Ur4nRtdmuX7mm6z4i0cbXIqC5U3ue+ApyBhweZsfl9x9l8N5RDOw3241oilEW9O
QdrfWge6PwV6/er20YnehFWtEapAb+CwT/w1pJWBEc4A6Hza6yJ8M3OPRecR4mmRF2GkkbymVc8P
7RKcotRoqIUex/+0f7LFGlu1sCEcVgvH6OfvTR3+ZGeHRiOrdnkniGAcO6GSsCZElWq83dR54lGs
D/qYDPrQxydgxwqEO848mduYB3Bl/V0s9GQeJT8WBU7iqh1tGCJ7pxTx/blvjRFPkObCbAlUXVLw
8J+F61z6VCiTRKpFplh+b2eO4z4zhzC8GA9pmasHRjusOMlcn2B1YE6Jhs4uIoQor4Eu0hnDoRGs
VmKWLHzFbYrMx8/UCCF1P1v/YGjUFd+h2CYoROy3wbu22K6JS1NkM8HEh0p0gYbwM5UJMBMwqGU7
7t2jcoM63Tp8DZczoMgA79fDdWLZjTJN2heALxd60WaBaOuVdzhEFpdtC+cfS9BU/OA6didm4OIh
iI1IeJzRP+/8nl/7z9PD8+C+leJ8QlpSmX+sc3EHQkmoXP/I59/vfU6QH6zhNuprYejoIg0zMGT3
5Cq/vQQcZ9EJaNgUx095NjF0/XIfUpcH6QMLerEf7rep5hktb95NiQ7sYT3YHRr+Oi8IKSM6odMN
oSEP+4kTn85WOpWpDlclR7jXJ+SW82l37NEfN0Se/S2Agpsw39eojoJzR4AJyHpJWwHzzRudoWH+
xmbrzpX0IMUEPPvBW1cRrpUftCzw4D9FwYUktQJkKKkuL4CHJRMFt24znA1Zy3yDs5RpmlXz+vwF
C7jT3+eMe0ymUXENgZpdTPjxcmNvJ7vlFMB3o0xtqvQT90NdqgOoQjudYgKc6v6YJ3sHVxKn1BIL
dTsx0NYZwpwPyhh6nMrL1xraL0tXayMb+W0S2IvShl6Bj10eFBKvFr0gcUY2W8B3sxZR4J5mSEf2
dA3SmNGh1sesmOLt4FfNLdCt3desp3nJr5B26m1npbKTqt5oJPQCsdAZMmjtvDgMNQwOoCvlFZrO
gLEL82B7A6+PtxY+/D/YqkJET6X6wYuvD3PZ5Pvhj22SioKIGwn5bGIQbTqMJCpy1cqoT5nZw1hx
d19f0M8i90SKizdKMzQD5wru+mTmo/NLMhIkEu83FxXTkR+rhnesqNbyDn5Tr1T9goHYdbrpyQDR
4G8WDeZCukEAk1UFR5kyLNY/MlQqCopvfHcqs42VCG8+zdFDpeYWW7ART+bOLVb9/c9UBuKYrAXx
nLfPz5johrx4aUCi4nvSts+e6jNRBZjOuNh3RW2Sv2SArDi6CQnIl2goaV5EyDSrKKDKmqoikPJR
twUC8lpI8iSzHAdrP+AD/pOhriPh/tubeEu0T1I9Qg4gPldXds7LeYPXIw0FcTBZcYbfhNs4CPE8
oQNG3QrWiROOPgerAyRUnnNZanwpWo3uXWfPOvUS4AOXDsgEoghQ+OOEmiij8wQBa0TOHwKd9IPK
TMoRFDtlBH0n9JFBorqY8STA3CdDEEUDPknoIyscgt8IKqX0sySEem2OGBC8/qSiGF6CmJ59vtIn
impoJ7Yhxz1yrDtwIsLUriHvcvFjqbsi21Tin7P9psXEtYT5EwU5xN/CYHa7wwPrSjdrDQK6aRje
8YfTupnjWBys6K8FJnWjQRyZ3qXPFB7luLSRku9byp8snSS9k1cBrp1V/IzX/kqDk0FFGZ/TMpcr
V0ArKUv+AFPexIzSeUc2UFslVNDBcaJJWvj1I445M4bi9JBaU2IrHbWObzxZJCc9RCJ2WUZqup+g
ye/naEpGQE6NkvxZDUdAc2+V0mWVD6PMom/+Ln2JkeXC+YmlCjjg9vQjzy2msgGULQzR57cToafx
3TAPdDoBoLXf2oc/uSM+Bwp3qtp6hBkTIT7GLWGZacn1TbsfxFeKObET1vkCMSzrOrhFIosGj6eW
h0FK6mXUqqsv/B2TEpDVR7KBP8h0CwaOt/bOOjvlCYjLrEnx0v55WjH46xyZR8eNarMwbKU9+73u
/5wSK+o6+dSx1S07yFa0TILj+X8ewoIRfk3aHdvHEGNF3AiqfG4C+0V2cb6p+XaL47Zhh0X114bL
xQKF5vaElvad1TlHn5uLSFJ2v4DLy6z70O6QGUlMa8Ya97KJBuo5a7CprTs0rani4OhR7OoCBwPY
OHwM4TxBPb/nbwdshYJUwxn2U/jck7W8Hm9mXN2c9FoLKARcE0ms8J0Nmvt8eZCIkoa7nMuPzYnl
AnrgVWNbtCKa2wC/gWZiOW4FlI2onHk/zPVORttgPVNaVy8/Ivz8/Kr7zlyyn23TGCAZnn7sW7Df
uhC5hURub9ahwPWaXOliTr66nXhOrK406a/ZAJUzuAOfuzKbsmpun2jYMGkL33O4IjqJVugsZkSI
tqSZxsyET2ZLjnf3Po0WDDvyIFpp2Rj1QOP/8YSOwcIXw94Gb0MyzlwTnf+RjduWEzfALt462SCD
lAwnDWS4/Te02WqtEhsI9ZIX2rL0unp90utzqV4952cHHCet5w9fYcCXsp9AhipcTsaUAKiiAu0X
pCGstflfgmD5OGSQ5r3WvFeYcpAjqZZOykhl3mcrIEqKW94CZIoX9cTZr8usJXtujgO1pZ9HGd0O
AQZnzBEwytpjo1IQpxcRfJC6R9DkMu8ITvJkPdH2kkkHB/BQVt8XplvqHFGWAWvUGmyv/3Ej6eTo
aY/VY6PogcJAl9rInW/aacx9KjG78aQtczHr0Qhojjn1VsmGWowllikfGr3MsGvlbh/8PGiXueTh
3dj2XJRYDAGjlvwwtGHLr3G52SWa1DxOkeptMC92WCoBGtnIV68ICMGx/W96sMfRf9e1fdiAzuv3
zmDGANIpVsnAlmDNGFQZ5D5zQ/Pe+NmynfAHCZtVLnLOVPjSD49pXU01WGziMKnxY5aAoC+DqHRZ
RKyj2z4bb25o/KAPhMibB2N42bVolIHc1AC5giWX1MSyUgNxgs5WT++NshIZLeFzPJiiiY54qaVj
LN15k/EUJnnO2vDc5pfCinoUAFg1wiSx/q3QGPGbYQK9r653qjdgd8N/I9o7nPNWTan48BB4D+c4
LbPUIbc5qSHjfPGXA3G/8PEB5jteOBBgcCqX7rq0P7Fzbc44WLHc9roRlkWPVaEmefrMgIwrqrZi
CtDyHmwmW6V4gvmDXk5FngWI0wtSd8BcaZTr9aedJ/wxvTF62VpZZd3kuBvU3wutsY1UAXW2ceoI
6l4wSEloEOIoGvgnX6XzpYrhblladJGT4Gv8tEVbyZ6yeHvMF1MIM5RshKQETjv1TIibG+a6OzOG
AgUS03dKhqlZXGeeOqBA0jOUF7JdDt87EKrOsptHMhhazP71W1pkiq5mjmDwqMlJdQ2ReXys7jzM
/K5OBoMj5QYSq/mlc8TkTR2fYmEvXikBmW6FOEUklgu3RTxdY/xGKv8maKTkRXsZcqRKY4Y6KPUs
gG0qlpm/DQkI2cwWaDcIv9MjC4AmIDity5xmi9+G1fB13eY36gdBC1UBIdhI4m4T6LcajbmOlyYA
pkM5LMLPqqa1zIsfDxuVYy+8tOU09ZdYNPrGg0Iqk+Z/O/6UmbfXW3GL9T1bK1cbSQEPxcMxdTs+
ffwTta5wTVNmnMxe+3ni6FASLBal6UMAUK4mPYaa/9clu+9Ff+Dkf6jnm3WyxbTWcyhhkIp8OIuA
N7dPOEsS7k/QiTFVnz04tSHkRMLP399JlBI/pkiCVc4FtvTLViGyr99M5Vs6ygh4foN0sQAl8cii
oNrD2wn/lMnWfNvNofI7+BiMnZ6UpZ/9ItcvAFwYKkDST5kqbmrWWK/V+UxcdKSviJpAUw5BW7wA
rPb0M18wbkDDSMPdNqR4ueUZ35h0v572DfpUc52d5cRZDje/ZxGAe5u+KhEbyrjEwr3R20NtGu0+
4VtLBLqNsnuLiZmqHQ/BkmzFWYcnnvy4vobssVv4dah729bM8fq8JrwZwUZUWFKk4anWqekyTISm
9WOdgnuXcR0gUfSVb+cbtoiAj37NVZOZLgUTvLVvdLrKJpsS1Mom0RankoX12vYt0BHrvse0G2w3
6xCNqpMvg1had3hc7wdTWolVVctONX2tE2DPQRPSqBPknCAYpUE1RNke1osj+bMLDf5XBb0CtwKp
y74qf/1z5x+GfKlOJzjAcOxMv+QQcFVWYg15e1QmjMLcl/rxx2Vnfojb7Yh9dPlERFglnySQ5vi7
It604S/kJ+9Vvy0kdv7EF9SZunTnIAulWfwKCLAcrqiW4NtypE/AYxNNo05r4PCMlLXbLK1aRyXw
uXCGrRg/EkkBQDWy37YUGT0cL2oNvFR2efElbrY1VREn1uHq+H8lAsvfO/Xv0cekVLwrFSCvo3Ui
fcbeNX4/2DltcIwCCJRlxzEDXY75CC31hxutqGD4a22VH2qX8hj1jhPUQkSaN1Bw3MtsFPvPovzM
AWtG7gOcslzGxdI+xcDau8Dxp1rZQmAtAg1br8k7EJBNZVk8HlcVnM22S+mUoJNAm8tvLlyPv77J
qvRmLYIZXlzoOIwN3em1MshMcjT4yzU4lKOG86y8/kpHc8XsXgPJZJ+uw0DqJciXVKyoR+vUSmTQ
A2Q+e0GwFGpozD9om89G8I2OzH+i6sttbNV1LAMpsX2pdjWXXecrYT541+O1mYEi4CznSz3UL+of
H5X3qyKCMHWYFshp7EesOssZC1Y4svqvlL+83gKQZcQKwl8fj4xw633A5ujKRoZcuggMlJwtKxl5
LZ3S4V59TlM95QO9QegTPdB/A2hAMZ1dqVloKdlu+0lyNMsgATbfRTApn+OxBer5Gtf5pGyDd0bI
YRPA0FUv6vPu8scrCY2Ngz4Zy8oFpRmEFjquvvp8H4aIea96cquyINNblDG/xS2h0kGmtPwN0HNK
+qn0IX6jrslCpgNoRVABXpIbcI9WnmltYflTXEG8OiYOwjraV5XmkawK042zvqit5NAFu7wDynPw
JvQ8XKYV1qEnf+qgSFbrIldege4H92Zjb8xI00UBwFdchWyIsrOARQvOEiFlYz7rU1EF1kAbYP3I
5GvH3n2LbHIovXAwagg6USet9AhMQAd1hZLSRd95zrSL3fSFji3lxQoCiYFPSd1DCHC91+cV3dHU
m+qNxlcM45fE37RhzRlv0uZrlI+IPuOchHqHP42ro48f0H/ubbVQYmswO29mTs1g3P6HGtMUefUt
Hhrs+mrL9vZrn+tssGvqr44b6vyasc7Y0wQjl4hFudIiNgmx6oiNbxOfGf0dT+w+0s0jYGODBdWa
e/XLDo8ypBacbzZEiC8KI7h/0zHrlBFb2GkxdxHVE9SoKMB/i7y0+VtbFNW62PyKkn7LVjfa081a
7l/sTBY1q2JM5QHvYoDjJxI+JeCb6s7LVzivnno2eqF9ByePAsRyWYYdrMBxmUPlC9nzyZNVIvJR
q/+cKt0Eq5sO8V8bvpMDjycPEamgWQWG4dz9Aa3/AYnhALwC48P2bufTteu3P3c7VmkMEAKEmbte
PbrmdQbknRhlocQjjcryKS87g3BFk6jcZVwM09C3SZw1BZR/CYwc37FyU5j3bGm2EhAkHbJ4SDUj
DlFuy8ZxC77kJ3M2tyJPrPaoXIXlnjSLLnynpiK5d651FuGa6HOpZJtowJe9mAz3LhFKIXtb7n35
SvCkdhnjQGmRjbjRPP8B8mgVxor77gMlugKsTjhhpscnvWrQibmE9BEMZk7jQ8rmZHpFL/NsWcFg
b/P9SQRXDnAeEHuZ3CV5kvAr/0qvb08PSickd9qknv9BK4Kwnxt/lIk0Rul3XK4mNqp1rwLhRbMG
ou2R2vWBaWryJmpm0KNucELjWI7w7UADydZQbk60DZxLF8ojiqZHyAjCpHUekl7tw6rj2GYHp8Si
BF1sw4ElA36/pw4fklb9MM9u5FtV7dk9gzuCRNlclXTvgCJA3wEdC896gzl5UFMTuk2vPUPTnQgM
0e8BaXtWaYuNRfCnylfjSUSDttFqnSTbUdbO3+aJEyjku8B2yY8Gcrayc5YIVRevu+iaZUN7KvuK
fjwNPaO+EgDjEBN0I1GaqEoDjc+PRsLJoZ4NZ+llZSHWCcO0jTGVQlMOYj+piUCt9TkQGwKDPgCo
Cr6gC1sKdwyanRGcqU/viXtsFIrHwBpFM6PbjS8NIC7BVt9HMwroORqtfWf93zvc/bDD2KmAAYy2
NwOD5CURQKd3LNAk/2rew8sLgBsp5U4GTnY3PNIxp3mtB3e+zy8g+g+SAeQVutE2c0/t9bQezeka
/ppM7+g5zPi8YQtCdYkAu6gKNOEwE2CnyQQ3+8CH4e/leXGUBaQ/dnzuE0hTN8FkaQA/5gvVTdZf
JgWHQBdYo91CaTlSy7A8dCBXeq4iFPrkAmq+njVmIN3nr71/Db6Jiue/TUi4KtUyAsQIdoBi+TEh
S/ljqTgEtdr72kT5ADwvTKHDHyqGfHuIXGl9gfJ7JyAdx0yk0++er13sUMU6RrnKFbhcnmNEfR//
48vBaw0FC8u8KjX8HISke8kXyfTl96Ni9oRyvPtrqTmAuD2jSfK+EZ2lBj3dzLGsrCte6U/TvLws
sN2wLUZ/Ajj4xHJa5/Z/Hx+jYGKBAPtrHsmseuUdKTSGB7a/jk0gp3llipi7/RR4cRl1Y+XSUiAd
ZvSOJB/TvVPKGcYEkQgRJpFEf9v8RlFe/ql0YEB98FRenvaxfvEJCl/uwGoeh9LpqjmKYnDmRUSR
2wAstjzPXH4c07UQYF4QnW9jHWkayNQw5r3O4zdpXZNTg8olcVosoWecX+Ne+R+xwS8nE0mknmgn
bxJR2WsvavRFCYgqPgWroC1Lw4yBjN0+RTl0yYBIZskR3b6XIdDiSgNVBcsli5rdkaEDtDl4C4s4
dCF6/SIyqpKt0h2iZzKy/sJhISEEotL1+QQRkFI9v4l9e6SACHDScBeE/LDsbcgkLCFO0uIlTtKK
X8m9W3710+LIE8QEvaw1gH4Jvak9roWnlaggCiTvQd+PzQhuvv8dDEJp86W5T2NrsWvDwH6ziY9Q
XICNAXadEV2Oz62/ZNWqF1iBRCAz8XmdIyk7Y9p2KJBDHXkSkUX2vgfYeQb4Zsm8IcN6VlmvDCby
h7RysOg5aaNouLy/gg2hLfAwsyg8Tp2LQMTbsuFjbnunIdD8CUnhiiWg06VdQWRy3jNiJUdvqXZ8
H7xmhD8lEfThdycwnou7OhDyJzw6vU5qm0z/IpE49akujVo2zETFSnNy7By3SdoQcbRZHPK0bP+y
WK4wJMLEUL/ehVDMArBT+5yawVYLGeaSwE9Yr3vVt8GBIrEMWcXTOrk7TkSOuovyXqH5Co2VqEyX
va864v5KY9eujZR7VsW2wEI1+7F3pIqfC1rs8PfcOoYX/QjhYqGfvgz6LbqXdJ3Eit9IDZ4RHX2j
lLdlVdooKJbmsVXvKGefEYANAk0zxyRopJ8Z24BhNo8znfBRyFKkV8yRiB16E4O148rK/PiA7hW2
jN+vl7yad3r64pXvru6H2lwOf+4HYgD3BG+T73V1hfLgVlGuhLJevUaQ67Q0O6Al4DS02XcHu49N
6/2YvrpfkmZO74sSYWqD9uwvPMabMoGUXeL6yZPtB4A6h2XWU8r+qrsXFW4ImhPO4X7LzD+O7W3p
rQgwvggaVyUgZv5SPc0EC7H1LK8JqZPAV4uHuK4Jac0RQf66USwLb9wXor4d3A8ybmHMvWwSfd+V
eK5Z/2CeYQPcJ1ZeqmspYNwPEXh42Cd9HTijnlF77WsJDto/H2+ZM0XUqlJVvSPMJ2OSQwwugH+q
cVHEBuI0rpj5TxDZe2uiNur+Hi95YfhNN3XDeQNXUpH5SB85P5K2/AOhYuc9AyNcYxZ2gVoRR34b
btoyowBgiQgKMwhBGRfXJhBKscWVC5Qw368Bds6eUoZzx6rMdfz/0m9GxmRQlFBhDNXpUqlmN/WA
ZSyjRl8QT6e/uasjjv/unHYmX1JmqoR4ECqGEl5gHyjbwWFMfstXnDkBj6c5rnAgDzyRC387UVpM
S6gbwrAAF4yanlR0UwiD59Qk57pswhPFTHzz3KPFN4FOEY0DszQOYbtIEWHmpBo1rfPJLh1LJeGD
XhZxYCMwUHXny6GRYCEr74qO/GNgTlkHkx5UCSIv7sXljM/8MgjSI1f0AZ13W6jH45svSKwHgKIk
52izmzeiH4zOmjwS60auTokYOCz/j2xdHD8wlGZha63FcN/qdXUAmUnqCj72CpE9yWsXTK3MgiII
n9Yzh7E5uv1F/xRpsA2XXGdgyQmER0hU1fUcy0+T/XTcO56QCgxI2Dj8EEd3vND7rK2VkL5Tbfqf
/KKC5UGZJbx/jkf/1JarD6xWZFA+g9V7VPIgajAMjLeeWIUYQqnVyZpQ6ZXoM2B2CwfzWWihKEbr
/WlT95YFGPacysbUyN6QO8aJcPQ1vDZ5VsCcUTQZ/1cDqy9flMm5H5a/gezbgBNyivGpaDHzmBEG
ZnUOtc9WgTXX2omqUxWdcUdaaC4VkISUXfB8VL+ofitQ8/0fm1Hxq+JRzFpez5XuwE3lJ/fkeyqT
tpuB4vl7ElByaRUU7SbNUq5v9log+BqLr72s/tw9LvkTtE7g6LhsuZ/ELwvKpRzUSChkgz8fgesv
tZ8GEjc/5itfPzVQc8wMQXLl4chkvsptoEgpsI/R+vhy53oawdZqKI1wUCCZI3t5QNOWsJDlFqIh
AqmHxK61nEXpjuKrYX9dJgbwe4UL53KAqXhOQBImQlGVY7ZhY+t9yr+/JWZ2KHvWZo3ScVapFviX
3oZl9kQyD5v++YkS00SZ/hQxwVewn/dmfUdjCPsCF8EHTnEqnJwMPAFeD397V3J6VfjJks3mKYDe
5kzNiflxuADGapYEkV9Z4ZTcQFw3pusTZO0NIHBvPy3r5hXBfb+gRYytKxLoSkEzFQ9lWBs+/nzl
knOGjG3Hp8GKNO9ghryFMbyH1KNIxiSSb+8XIyZ8ngRcj51/7N7aSRgIYB409x0Ya7Iv+BEGTw3q
QX3QcvmKvpHasEFwvpxrhuX2yl8LBMBh6Mz2LnLEaFW9W422qcWev+BzEVn8Mgw0jAyDbkEl2+D8
wBNuww47k3iI5IqZiKOXGKvOYz2Br6aqGojMYKn7qQ3jYd9b1JxFGNgXRWK1UZtyTk9UjDxD2QBU
BsFRJdjPhHqAahDxdrTVjLninMU9BShnjs1unSNGMuKLvt6RxP+FrFfwPaMdJLSj5P9tUX2uonar
FpueZSCCjnQpZtDxTlvFTpDX7OOf+RclRlOaXuS96ZyzUFAebk3/mn+4ffIWBkLzWubO5knSazk6
CA+OIZA5+UAKKjO/yhZq6Q7kCn3Jk+FishAjRA/L32xa8R+GCZMl8zAuaUF1JR4CP5f5MCCmm1qG
3Dk0OP5lc+DfiwRseeVzSeWLecyBGo8Y9FBIcljGg/YOumIwlkxEPBnmrlExBdozu28MiJ4ZCitx
GNiMCOGDuA3AaRc0oBdwdWss/u5O2Ez587Lpq1YXIdnR+UkR73zTuEJiETDKAgp8V7VI8F3r41Rk
UER7qEuOgaWEs5fo83ryI+YBbDdSIh0sDgO/GmaoWJkgmHY6wF25s9qXd4qNVni+WEgQxV9hWqRd
o1wjpv6NHh8rtuOn7Fq8UTXvKjQcHupJ+YN6juyMloyRGrzKGzvDusa7gGCX+K3DQv9gi6cUw0In
KHuATun7xNqn05/iCrKNhpKsPsNjqJlHdFE8PkNMSCn1qHG4E7qzBo9AKQuD6/HHMH+c/ma0fpqs
R3vk2G0/CxIiCRic6Isr1HvsLT6aDrk2va0GDmfFTFrhsuAsstYq2ppqaggT/LIcHLjDEhcjYxLC
f96JT3ZJNHaHfbvcHoL09M2d5mfoEfEMSGrHN2t1yJXi1zOXYBCBI6QTH6UZOqC9059Ln5wgCls8
PFHet3nWSXngZm9IYmiVV7MTH4m0Qgne/ES3NHXcSSbHKqHE/n/1mZh9L01/CMkTgwMdKzuU/oCA
eJUsZDk8aWYiQTtHmm+Jl05k+pWvNtdNHs69Fo3U2jp9QhcTpAAOTSnS7Q60cy7XOz6Nlf6urCdU
nUlMcHeX7iaxTxhxaUP3U6HU16XO2ArsOZIWOcR+zdgqMxpQ+RCnG+/nna/Pvyz6TFWLF6OZ3laO
BMmkQtVuRkscF8CbQfBLtMJG5QWShPh9DAfSY1dKJxWoYZzDSmgDoWioMQ7NVUvvwzsNsRiwp7EL
odQxYh9HGrlIBcZjIkBmSBiTBCblPixVjThaeOM5av9gZnMTs5HcRwOxC259M+7a/amn39kot5oM
D3sJNJOLn4k2DF8apBAAsHpFseoxyQPPmk8o35PklIIt6kiDuaTKHtjw3O/6yF+DC5phrXyKibDJ
Ex8VhtRQnIA+SLbH7ZrPUbBgFY8CJMWDOHm8trF8/1vXdy2k9cz5X7cUWwdQKRA3tq9lkMCTd454
96Ghq5sgLsasEmRUjexZiYVepqwWkZ4Op/GX1HvSrzYcJ6J3HimruCBHm+ip8iP+KBDDQdLt1xsz
yl77mAblBS7W1d5LFhTvO8ppMJuC0xtun+oP/+G9D96y8ibMfb9yMU+ya+lh3ySSp3wS6TrO3YZj
zyXtilXL9EH1lT9BDs6Fws0wNlJevd0HnkttEAm9K9xs5RntspySH0LZwOH1fhtdmrTbUgGooly6
Jkf2Bk7z2b6TBRPo8ZJPD5vEli/+AWqDMuonCPwF9fwP+/tW/8LdNtkJZXu9Zn2ZpcY/9OWHx+T6
0WqoK69vZxYj6aWoVtl4i3vxpYHqZiRCm1wmCsNdJo9OOtvDpeze3bNbYCwraRfum8VeNUeC9zGK
BUKhiZ9gwfNFMnPeI5QH7dy9CpPLHmJYkjZ9sVdCMlCpPQ9TSwJPk3fxwRbV4jCSXZiedW4CWbTB
rqvh/wtfL05yrrD7KMV3nk9JvOD6azZLpLze2xcgYzcPhmgaD3ShTueacu/VrvRgswTYHgxuiz4M
aed8eu/5vCJwvhuSS0PHcL0uhHrT8PHoL4sfXRO1/HCRQl2j0aX0PW5sOtfhqdUxvzGBxI+SvfgI
Irw54iVxbj3x5aiVoN252NaO0BzVM4/xakNNMf92n36gzhQO1IUnLBHwRWvGpwLk3I1dL1RPEHx6
r+NSYXRMp9M/3/uUchhQazmESH2uADdjA6yEVYLGeia1TjjmRF+U2tBcMGHV/q17C34Z2y6IwbZl
trP/BJGjnuhkf5g+NrxeQfaMmKMWRrguV9ZWdmI7MPxNwthijSgcY9a/P1cpazYC6WBhYMysfeig
SGheWCoyTKm5AkG5MAyLgvvGOI9mz8twQW61YYnV4ZU4BrUthN9h2/Cv2T2IivQC/lhLyHmaWuEC
r1jIpEf1dQjyOYCuQIFIRnH6xp0aZRALD8B2j1OolVMxf5DIUeA4jXEk3Wu/2tNV7eq500njSMkm
ewqCX/BYAF50OjOgyBOhi8qHEj472K96b/rfTC2AZmzu0QrIW8gAU2fDYEhUa22exaDF8plqBKpN
0a12q9z3weo0ETd0mELjyuaLHDuSlcFnV0jKemCMNZYbWJE1V+6EyA4OifseOzIeoo3znTSyr/73
UzK1qmRCUNTpAbTPgXhUw6aYqB4sFRw7eYBn6OrXq2j6IKHIXbH+WXkfmGes6gs/F2AYa+ZQqLYd
sVgzvWurbyDR+Di+wjStgTEegK9PgcRY40h0ky56XFockMtsi6xCs06v78hUmHE3ZQiCHz86rp66
0/tScgwCTxizrqD5ht9mqqRhCyQ6+6KgMNqikg5wmh3QtS0lfxAQuzyajpkR7kOYAk0VGPFcAgH1
1wxIewNR3/g2Edb84IzI/ygFZw4IvNqPyythlGXVOmoaNJNiMbHdVXbAcMfPieIC/tWavlpalkJK
6O34uRVStvxR4i/SNfBx1elBuUFe8DvssLY8QTrrYND5SiWieqK2KJZhEmCpsW8fPhdA+PLPkB/g
LBfFGQ1j2AO8YoOVSexf56Rko2xxHSS3x/Qp9M2+Ei65yYbEV7cGjziZamQ/SeW66xrKKWc5iwTf
EZGYHz3OK8NmlQK+6kB49lBF1T6rOMalN3yOlr54XZIsdp/iV0gbuUtSEqg51/NHYgnp/0xYyndR
nE3kbM2dBMlmQLYBevCQZk5HU6VtVRu5PY8zOdw6Ubwxf1jLc9153zQHFFKRl2eA15EPLWGl3Kkg
3kf6AgFexKpoyU296enQwn/LSiUq3pWk64UL5J1n9DbohH0nimsSrRpvSG6/8NVTfc48jCMFViM7
KlDL4dzj+QY/Lr1JN0SeJEq6GnFyE0D9IVR/EzgCvLYYYKpIhzhL5uu5CdoDeBc1w4lEVuAezw9i
Ot1fWj2CsfdvHLha9N0Uiq0p4ZERDZfMxRALbLe+aLjyCZM23Yq/E4WzZfHOixlonMuFiIigwPGm
vHM1BLVXJt8A5dJCxyWDHFXexued4gMVn2PxVE+pLzF3V8GZ/1Cy7XoCWxKXgy/YJyUxO1Wv2E+Z
n8sLDGYdD+nXuElUxnw6di2bodOiy9DZHyZyBRb6lrUBm65y8kcoWQxzlJvqN/JK2cfn92r6eW+m
Qbp4ylRwgcNoCTtKAOqN+u2nYqnO0rMlkBil3IbIC3R5HNN9l296rnNrDzBTBC5Hl3YTxs2NmMY/
oNH0kQUP2RGo+KLMLYKmUsDDs2wei2wL+CecVxV2ihQ/QCKNLy0sbS+Bp/jI33MN1CNE76osaach
7oemWTjkc2WkDcM7igZDH3vViyQf6pwstZ3QZ0Y90DxFHuTd7DzbISyxaSmEPMf4ptgrt6hYALav
6ZwL0nx7ASFOczej38eyYIT2n/D/8uDan1CfNTLr/V1sCOtzZUG+uPl3YxyzbP6YkFFObeypcyJq
JRmmL/kGWYDkua1JwPoDpCFuhmB5jwOVorqH2j7FS0yyeai09dA7VsD5H/IM0w3oMSzQIOsS8PPh
wxNx11MQfcly0pYGT4K+CPuOiSovB6oEygOJGzXci0ts/USW5KsVvt/bNSve+djkosd2LciW9fPZ
UQFJ7CP66xMl2fe2bgqx1x6xE8UFI/l6vjkR21TCzyjJ/6LGpveFP6WTt5xEARCGGgNN5bjvhOkt
WZfnvvFzUADCGbH/yNoceHyx6tkE99kKcISpLcVn+954RDqIV0iQGbDvcEqFiLIq11KXpy5a1TyP
KglcdxjDgMTtP7LvxvVDiFvU2lSawKdRq6xcrPCnI0vaTtOpjEredy/m7C3wBevTJkSAxMKSu3Sp
MM/r3x4cXbHv5judn5vvifH1wEJMlOlV51VrC5zBt/IX7KEg85xZvNQA13J+8+PK3l7Z1ZspYJYL
cTcKLNCGrlar2hqpx04HZOwKADreBQyKBke0N+lu+V/63dOCOJzA7XAHYGfBFdQGNsnOy2OpEhUN
OGuUW2PiAEqKBFDR3uqGJbTEVv5V3+x106VsEtIeTwzVPpCS2FLbfYSi6aMzd4D9XeWnAjir8dUK
1lkSKv0ySBn9l3fbLTQNnO0V8E7KdHkmHJCugRc+WpBD5dPHqAB/7TfGL4N0nAbc34G1BPqBYmhk
MiFYb4fdwaDLZo42RRevCrZQEECDGBRUPxExxktPg4znWEo/+el5ZkAzWB7flQkovfhzAaGA0NkJ
G+W7/qa7lxz034zQOE4Vfq5xaUtopFoRrHrkf7TI6loUXr4Exw6Uyo1fGI2m4G56UG1nnaZcyEi9
JcszMNYUpM6W+bvVZrLpnZXOmpVybxRKsjPEWo7QMM4dIWgMX5WViTMe+PSMAzL22/2eiN+g1DtO
hznrAWsomXCfgw7stGB3/GhkMzVVchiYmz6Tm3comvucGWDWd/00h9k/4z+clfh1HaHpxF8gQ1H4
IyOcp22MDp4dBV67CPVJOkxOoRU36t2vbNsKsoq8zKNnitrIJX7X3agOwNkDaMVsL2xB1JmVaAmv
2QualGZGeKNyuxCIDYs4uooxV0CWyIJMgfoM/nLwIHBzybDijsp/nduQNyvs4t7yXsVc4lA9+jsu
Z1vobjE5mTR5PUwD35KVQfg603c0KHZV5h4K3H1JTJnSIQWo+H/a5qKrWZ8DXHdkLU9Wn2Fj35r+
CHD7rKEOZhK10B7h/he8HmgTPI1x8b00NuCVUKsmlx/aDR0r/uHdgjgw3tQxmZ6jbB1EPJRb/fGO
2OHBNxcQWUMnEWyK3x6fOXnnbtHPV+ZvSZFwVxmb+p2Hg2bgCpvoOaiEnQoySkGJGZBzL3Q318NT
LSjsAZizXGHoMBQ+lLKBGYFwznQafXqpWmFaYcU0DQuJjNb/qI66U1RQgiXewOJVC44jcEyRYJCV
KoFDHaqwuxVEl5mEmo2Sy+FdKz4nTRtaSDJlpKoF3Sxw1wJi1J+CGJoNdoUapPbwLHa36nug4tS3
l6wVpowPQpBIfGizHYAt2H8zsTMsjn/YVGouILDB2uxA3VdF5AoMH9uiY39aAkhm4NGM+Uce5oV2
HangSBF0zbHFxmeNgC7x4U3FvYJhdoxYv3S0XfeYuXiFTZSxto8QYeRQauc5KxfBGPn4a1KBacEL
TTi/fBHAh7c9BYy62xMT1ge/eGyYi1XKvJjWNVTa63IqFgoRadz+X3Y4vkvhE6aTk1TOZkPGA1bA
0xwdc9cH4ZUVOTFIHXu9bYM3iauSPGs4kTUgOp3LJfK/Mj2Wf2qCpyJpXcOKCVI2xUbYzFebUoED
TtqKexuL4su3Cm9PTHvg9s2QnUWRW2RU8TPCPMUEs+mpcmIqkmIByOJEzbqrpz4rsjdgrrOK8Zd+
ZjPWGyoTR3wCfyvtLv864jbuLLAMRylUd1wtIDB1kqm6vWDlBmWapc6o/ZEi0+wc6C5MOQUhMD2T
10lALzP8D4Vs/uZvrYpV69IRwz/jfJe2AfEJ6AHWBLlpcLtl29riVniC5wav48vfEsqrIRMZlapF
YIDOKkyUUPiRD98JcNMexZljyzXnImgME+ZkPk5FTd+Y6q7P/lD6Y82ReLKpn4trn+1wkmPupOgW
/Au6LLglOA7aOIPJNddsK9Fz2jwLXd2dBK4XXasJ0TdSHRc6iaY7Oc1GxKUsH3raH/91CPqXlfre
WOh+J4H+QPna5dd7gXgh/NVODy5xgDhHtCb6TLSCfP7Q/lbhs18zSYa+WI5yIu+06Upq5m0SzuOC
S60BBG7rWg3Cg6ttUW7ZAZyWWeguY8QppkRcbLUn398rJu7iixIyNEunFPP8u2pF7ymlsD6g2uVQ
YT3KuU5FS/tjrG0PYMLT9Ti5DZcljy0FanzwixCdWa0P1Eurkix7K4Xi8EF5OYGnk0YewvkTQ3Nx
CszpKeA3sSu1azxW95I3Rjs5+2wscsqI89bT99B6cIhO0YOBy0FfCft6C5DJr6ANkC5rB4QWWoyL
SEli/LGd70VYTQcNCdGqg42caLiBZVozkdEQQTXXXtz32HhTWOIlDCwr7nYrBw48Q3YyMDZamjbl
Ay8v4oQETvzTl0vo3JIjQ7B/Gevhv3xJ2C/0Unl0Kg90sLhWDzKeIpb7XxyAPjNA2G8d8RMJIUAn
Oqh6GUlrLSC4KRs3CVksRyA5nht0pSo71IBBOdicvkqVv5x6MgdHVjGwbbULZYdPTk4Fq5cBq4XD
GLohls0LIIfOYICNmetMIt9rUaeEwPRG45pr2Y+HSy+aN9BnMALTTiqSqgrbxNJXC7775aIhxYnF
mfS4RGeLCcwlr5BC6IRfzI0AWnkv+PUapZJlVK4V8egSczum/W76UBiYp474ozdjaXu7AE+K/l0x
3ZtD5574DhePSB8NO+2lFSN/3+6BHyCZ+y99uc8b5xyExpoKzg2zdF1VAHOeoqrUI2nfF7ofJM5k
lTjwHPRbp/zTx1oeUIArp0UZkf1l//QtI6vtc6AiOcEwP/LXUsGTGM6xL8H7q8XculnLOQNDBchy
X4w6r1Bv7NC17Ah37ZI10k4zhP8jIAypHAAZlvovakW+ucweBk1UYEGbJwXPf+/FWqRcIaamable
uYXwp5G2nwY17IrfVMb9YIfofl4v/+02+7MWXxHwuetWavybxlF4fZvhfqrnOBcmWVZuo01DCEhw
FE7PdXtgtLJfb2VosfrE26wd1VfQ7apM7XqCqD0EolkUIa113bpuFemXlIrYO5CLJM3NGMQycbEx
k4tXvWWl47HGr/q9U+i072CYfnZIc49ZIDvdT9Zjqoq3BxbF6cG3qfL6PWpUG1zUszgK2xUEQazY
0s4RbCKthwmi2alTaj4A3/7crZ5XE2pXNdKxmK94JWRLGPyyPwblOTE24jLdtk+zwMWEbZhekSmd
rKVcDci6FSXaloGy9ZxLMgRQouzyegelYAAz6hzfvw3JRSe1RQJ/WJFDc6N/AnAlZDxqxAIL8JNW
0mqUv9HQOIptMri1sUXDDoRN0gl3Fm1MSVadaPPVGcEI+Dn1gQ9w6wuecusPzZ59paWAF1jBhs0u
d+0GiM6JGjqHz0CPLCswSsQDfTpWTAkLJo2Voq9DK8qdoJjGXg3TwLu2Ac1TE7MBCgOqJa75l5a1
qBJn/8aD5T1z7BS36IaR4k9cpMhPPw/lHullmxyWTma2ZlGaW4Hehcxt5J5V9ytk6OFAuJOP0RDM
4cLRXj3rMb9NOa4EXzJh0FyhlTV0+GO4A8hcnQZzsW0jlGwDJFgaIvpN571jUB9KQZVcizAROGXh
nE5qaMq1l1aiT/H8M2G+V9SwOBvXjB1VZIh1QSL3XepISHKhzLGNtvxZuJhRibpwApRcT0c+oKWC
MJ2ldJSE5XTV54t9oaXO4t5VLb0VxbikX0w0X2O7jmdECxeGXLsyLjItWr58hYiSDu0mz2K+Lz4M
EUUR5hLmMci5yxq33VBNHoZIzYshBikeXTYwH/NQ14tH7PA2IlJgZZt7/zIAz9PkpxFlMWynL5xu
W4/jRvHm3F6kk5zlAemctiWaojryvnR3myJFneRJcaSUtpYE85NB3yHKAfM+M09JIpHYB/G66/mW
hW8R8gfu5LxM1dnbY+kDyWyolmPGnDG6SECUg/v+Un7cb9NYxfr/lCuCfO9T2ALyyVwJPttv1vvZ
HtuXHwAUusc+Bd4+yH7WMe+tiHZhkAv+8TKei793gH6axZH2EOEyWJ8yulyQ8FgS52vSjKJN+QdW
2dhtMKJrt+ymf+Nq1YLNBv5xkxLrng6wD2xwr5S+cCAvafGfGpZ/5FRuUaDPuP0izOKYC4OvFWJ2
d+bB5J8BnRXgbRoCipieb9kTMflRlcBve30Hx8iBelDFLxqRGcmqWEEfnbdYm/X7t7Iv3MrErlwV
Q97+JoUKzgwBRmo8cUvQ4FluJQVfH9tLO+O/fHHSUkRKagatn1iwuU7uStPfn6SHQL4NstQBxM6c
dI9jSQi4WAq9uasWH2L200iMX5TWGgGn1p9tgOW2XXWYgmtE8gn7qQz5sNu/wM5gcMQlutqUdvnw
l9fN0ZxRWN4gPeidTivlwNEr4nULbbbCysb9Ga4SVrXuRq8Zq0z1RDXmM6Bac3qd5XTaj7NTQVpj
aW5zKYgZl4J53FFAEYPKz9I2I1KTmCPMcIkRPpc+Q7vlXOCvlIezIk75h1P+pTsbNNEh3VJjkOBr
1HmMtP8+YofU31MrbKRihEUcI9BDCjBAT7zS8KLqM/8hn82L2azfPJ3m2hcG+EErf1USXWfFgcEE
tVkXfnNxIPsnZ9TTs5tDq8YK4brAheZxqFP3fPBDEyeLXEqkcI4wAu8IkSGAhz9mc1iKjS+e6/+m
2Uj4cqUp1xfnGqFKlUr9FXitbXrE6ORZtyDHL1ird510Wa+sr3XmWs7DPFer5/bjW/Qwjn/CG8Sc
1k/hUiAr1WxQOvGhSUb7WkSdFVIFjDCEkrgjLmC9kpSVuLu/H08aap39CRlUOZGgVstGhC2wIYFe
5R3r5OLnnsfkJjRmF0zbj7+Fum0Qg1foiPl2V0GE2XYrhBu03IOlGx4okbgjraU3aTuBW92yeCVH
RjBL/0nKUjarObq03MH0d7devOgdf+EyDtCgNBCkQDznwHjmJIxC2kJZYkZWu4MXYXp+uWe9/gd/
yP4sBUtAIrH6zBvIHayLI4aL44zsoIPtnXKsvEqsDjp/kSZFlmMtUSJ2gD+dYidNCX9EI61ecQFg
mT27d2OGuMC92Bkv/IqJvXEZkcbcqFRrE+Ip5V3H4IFTGeHwkAxtV0L4nL18pPnM9z5yMZD8EcNg
Jnp0NI4Wnn1sEUXzHlohYYMc15mKPJqc/9izsnFc6+jpV6wGDbWX0EitTZhc0oOk7YxPKoig/B3M
2LPrV1sIKnkE5UkDnmmcd3u0zx9wMLlYkZ+7U3kvmrvx7PWryVna+sNzI8Xc0Lzt10rlnNuFtCMQ
TCG19KSCdtqm7jNB4Z2y7t3wY9y641YdjLOm89HkUgJ9xA9gqR85O3TydoIyQuJ0PWkTzrnQPM8B
FeLmZeDQh7cpW6rEyL0qPZbRMxSuyq8z5KbMRJ/7SVWOLl3H9kYZwzONdaUtYNtgL6I105P4sy5e
GM8RF/G7LsbbwQFtGFUutI3cmt9JI50d/hxHrfOMKPd5OJajYxczu7GCIoIhpHIGJxPGMAPihGVk
iBLl/ntYeP6Acayyg+Oe9C34vUkcqYncL59Bf7oVKYdA4O2SMs4vHN1cVZPY3SGeh+aL09LjI12P
UagzaPpFSaeTwIAhrFYIzpeK8dGZlDQDjDKGh7cJStnYH2g2yq3ZEKSgqcBCPgDNGBX3VNW4R/er
zRGTuLNIDCgNr3Q9tv6incI297SeJ0wMu1UuIU0TMWkWydusMNWp1q5nwOr7iO+PBVAYL/W1d1S7
V3QXU/07GLYPS9YuPzMWMAMWdLlne+FrWvbZ+WFR0BJpnjZ3AJvDaFmIeBPabkD/04kBWT45WUdE
PvkurO+IC7VnWrxGwsVQ9NibB1w3zZWu81obLN66/Lf9mXz6fKn57ICtwdy1zJ7i6ejaw+Pp8t57
jitcuWhMObNPl56F7VZn/iXlda0s3iGZPBSZI4w/aQ67ZuSdMo1i8W4+G314wiuPHy4UuN6/mItF
psKB62uhbfgnAtixLKr3N5x3jRwFuF62m1/WFKOlOE2gM3UbQfb5BxQVHpUNtstGObp9gNEg0Vtj
zGkAGJhfgCTMLdZXaH0481s5J696zaZDOcLOvUiUgEIE16w9VdwqyJEEqF0YqnxxhVnyO7FkEvgu
4fXzrw+uS/uMBsF0/W+9cwJ7Yndx29cpv3ZEJ7nES4xOGj6VtIY29TKaMwKYUBQhshXooEBIXlV9
46aPd+0O6pcR70oxLafCcsxBLkUCWzSUORdMDlx9DrmVc++Ngne2sPlGjPZml+Td06Pa/p3IAdxT
a7rZoOIQ57okF1VQ58AU6FWBcEotdOf/i/CfmSpIXzdVyjp2iK2U00vZdwS0W3n1aGQN3+X2T7Bd
I4gqB0RC/Cmh7NpYWrpaRjMQBz+73Spq4IBNWVJTWjrZGlYiN/eXlD28jlFvK5c31yhJqvzFPMEL
fUeSYVBHxNK5tYyf/VZkx5RRTW9T6s4VLlpLOMj8UKN/CBMRh1/7JMrR0kjt0x/vqSH3qFPD47Of
Wayg7zdJmtf3ZTgr1jddsEhllqbySNoJ2gXnQl0czi9WFGCA1aWmX6FyUvoWXuOwXaGidsUfWNsz
0HPlMTfDDb0/My7awwLisNYIpeq/q5r1duW3OQ78i8a/nqP44WXj5CJms2J0KUlaT9vjva/mMhWM
60EhMT7RRJWVdG8XE4y5wWv8Kocbg5C/RFM8oRY1kL6BYd03rhKEk2IDYkG1GFNGzBMMNfEQuZ0T
Q7sMigkvEUBE3m94kSNbwXTYFZSd1yuRpxUJkA2NipueK/Aulu0PNarOviFth9EiDILkBz2B8wdH
pWhIBJr5oTRe0rECOdQwmBv7G7h223lgLLvA3WVyqWKMwZKzDirvpDC7xWkDHajDbeiHWeAkXjRv
y6XzY4xwhfvFGdd+CGGAAN1XgTs7PyXXa0PAu6im8WGROUj+ffFQRooh55OUFPzlin9v/oCIYNdf
HuKIiCSlSeTIlXaFsXM7rMT6fDuXpaprUgwyXHriyOavz8qszwSjWRwwT59i6xI6Nlhwly3cgctG
MIp+YSViA7TIvZ3reQO5G5AzroCbqrSug95A5WZV99qiCVkj1A3cF+8p9cTdYWGzrFYXFNhKs+y8
isGNmjHFJ+UBVO4SX58NiLArEq4K8Cm28xHx7cX3uoC+aWJ2tn+EmXKWpTmQgh+LSWCLvy2SUpMO
decOJRQyWngePco9HCAaPwiYWZ1V5mQfL0WFvfli8WWO9wF+N8BQvFVYQ3P0dAJ48f/yGdb06K5L
jZ3Y7cDR2QfIAoTVOoCWabz5Rb3SHffJ0htJwpK7u9wDI7BTU/l4H6uBL5RvTGsh6Yu6s5oiC7DW
XPCBx1EY/9UeFFc828XUzHGIAxI9uDYipa2cjGhLxQCtwfRSAhqemJXvCsMbm67tGh311rBYjza2
9ZMJqOb63z2jzNsavtEmMcrPxxyJnOHkAkLw1R5skDlp8iYVoBOh+9tGCR4761O+XeIrAH3KbdE1
eOX/M0lt7Gx8lbktvyABQ8qjPLD3LC1sWx/Rm37gVFi5MZUa7ztWW/PuU+S1GTfaDnageC/4Ih6F
akP6xTSikVhWUf3lCksurKd13dnWday2Q5iXo43hm44QD/B6LF9e4cw6xv2lVKv+xLkWR5PPx+7a
kfVZu1BCJU4qWLKnEvD8G/t3Bl5oLjMijoGQJqp/rlXgl46hUR+s6xRr5Us8OILzxhRD4nueCNgA
doUUFsKuQEgQESt8dc+xYLOAuGaPDQuKslCdkko/IS0NuBnllrbtVNvNo8pBtSevyscWJQWbZhqr
x+MNRrj4UsOyRIyQKsfK76BH8ojMZCiknv8K4bBeyFFPAteFaXBr2sFg0dO1CaxSGD1+YFHx8aJ5
nT4QnrbwmB6ykSXk3T/O2Qng9DQ3C1w9VB6E9dbq9A8arhji9KI2/14Fbg+XRapLzsS4d8zDVZ1w
qZexg6RcTOBRT/OWN3/0WCsokEZOpdC+LdEbYX/W1M77Gzvu+zQmQvBD8NJI5oOF9em4v63pwVeL
jipS5Id0yjgws+mZyKa2V3BCxITuohfmmP8RstT4ymCYsCva5njSh6JlDWyUawz+LhPF0MAfmG4u
Gl/77LM/YSLrfmw8kxgYCs7SwG38kfuXJCakfIy7yvJI7Rtw8QqeFvpBU5m+tztntwDP4sPUbsWS
cJWLEdU69tbJzEBs0M7TQcD/AWsLOvfN9o3y730XGFqh++ZYeWHeav+FUUr2QoSDka81ELaryUdT
LXcgHh04aE4INVnLOPOpYyCBL9e3xdvphD5Si7Xxgmu2chbamOvUp2cX863IO12xAxw8ikI53qiB
H6Dvr+jRINF1pySnM363oAfSL8JEQT1wfK6QzZfvJCx0K2CV+bHm0iIx/ppwfzAttlW7emI5ZdjY
FnJo8fHyfpn403yASZJbm0iukE9FjYPNYvRyQjYH9uAZc7/QeP+xhkY1ja3zdkYqp5ncGDA9Xsgq
DWdMXprA4nbvIwDm12PfQCVC1aqVhIFhGdjtYGCMZgOEqkLwQtVUVseHLRaKgdt2PBn/X4hT5fM0
9jmvt+mMgABrSxW6ChGy4utvwPx2FM/qBvoNN34TdM77hL+nsi5r60g+7zp/rkAgA3PD82b/dASC
3qFWQdZgaFPo4pVS1rCz+PIdn81yzcjyXl3KwgWNsdnnTsl1DD7PY6Es2Ezj1VW6+6lGoY75mqPf
G24h0z4l8maxrrNWrXZznCy/qatrN/puxC/aCi3CPTO5YeFbZcqAQEMFofnDXXXjnuNPnZeycbCC
oCGQedYrxWqF6L9ucolmc/G8aXzH0pY4QMc3sWhYpdZdcfpeqa6IMusXUeJSx+ACym7yvpx0KjlL
16YTT91Xeph5sY0ih/iaHNjDUwUxa8ppdwkLJtA0uCezvQ6Wjo/wA4g4FuW1K0sHRN/b/o+JktDA
ZyrY1LRn/0UVeDBiygAysAknupiQLZJE1HpzuLSZZZbI9IqCUkyKMRWaNw2MAxIbgXeDWd9V6Air
G6ydejdl1MNFLINW0FHwx4pkXz59ycx/Uc84B7b/m1fGGHh5zOqWEXdiYSBpQWJ3rKR/zXJBLVAu
xhVsJgw+ypMtSJOF9Lreb5+B3SqlzC53hy8pYNzrQEzcjnKdq5iOxy4yFeTrWJDHqM22SqU8OpeP
JWM3vrpNTsCnX96ER6kBRiB/OiyUu64S47GsuS+7LS+HvIl0rSHULgCmaJZW62wJJwFaX8QvRR0S
6sgLLgYldWno6KPuIy1WAa7a+pY/FMUF8nuVE0TsFbK8YpVG3v7fZP746JAg3kFa/VIlqNNHOkc0
1agEYk6PTNAqcOQFGIewlPab8GtwiaA5klOZyFXH4r/Wtc2tazmQdJbeLWvWQ5vEDw1CIPIIqrfo
ba6+peVRwxSL3UPHFgNimgeDFRti01UdfoVxM4xkrfuHxpvN5YZEeFxzmhCsfsVRjDG99Yq8oxdO
caK95Uj0c48iJTVs5Rr0Zu+ICc32gxoj5Y3wEyFdJEMZxREc6owHOkAiXyV3QB8+47aX974wr6QV
f4TJi944YHPrhi4IEnfAOdHcAc6aSZnykJX0jzaycOi723EyltQPcM4mOZO47Bpxu2Seuduaamfi
VZRIDYrKDJnrQ2Bg4YEygy1kpCmDNzYK02K8yMZsWsGtymU3cfEZ8BIDUrK37PPo4sLVa90+K1pq
lej3wbdyQCXb4dty15JWHnSlpStzIGZUheuayuJIWSsf2fE63RyK8PVbNGlaHtiRvsu1mkrN2hAK
9McxCGXy9cAPDVb99QXR96tlSJ43OXsBvo7NdrqCQUfRpg/KiCshmswEYW3XsciANUejOVAZ0fAW
pEJtA0OmOLSWbjWUX714dz1ReMKtY8sUAohKzgtfUVwzO0/imqTHb5O7N+XgzMQJDxLFWXOIOOdQ
jq4fEMKQA3816wmImD9nU+CXOv7Ryc6W09MLtArLzpQUK5450ijb1vOzJByFZZiGcUwG+q33Cawk
+LZE0jdBBhKqOTKmz6bm1zgk3dvaS6hvwbWy8lWp8mvj6DNQ7UuJHduTVEu8tSNKjNKShG3ufuaJ
cIQda9phS8/Lm55SXPVpa/zouSXDzTPxxbaVAjxzxRXkcF0d/HQln4l9g6VJrXzvUSNVORHK/9rJ
MmTtJ3Mbf+KNz9uKY5kNC07aGP2Q8EarhjMX6yHGzrX1mp/kj8S47/tWKa7sa5uBfoQPxihIOQqt
DNnDakWuHQoSKxK7gzQWzpmMSVQ5EfxQiIriv/68Z98zb4zgEi2zfs3A2YwnE7gg7+47BvMJH5HF
cCVCao/qO3CAfufrhS+x2FhDgVvT5sWtdNrQgbGNKnQ1IejqDiC0UQ69mUCl3NEJGULWl5T0g6zj
H/2Tj3L82242BVjxuoQB2uGZ1eTKI0J8MNESn71ItLKARCvOupIt7ES5/6pf/U1h/XJrDEVPIjQL
NA3mYKG4SUZVYEvQiHsvTdzUaYaHKwcMbACWPvwbQdGyiX5U0HQybuYlr1dyDZCIoUAYJzc90fW/
o6MRgulDDrpzEUuxFYBwwgZQC7g77h9ss70/8f+Y8GixWV7PkjlBYUF03Rnzk+jeYN38FW6w4ABf
ND2suoJjAsS/1Jl3PWZabJqRWiqPcJQ0Y+WeYF/HbyARMHwNY1DBtRVORfzpX2NVwPWPFGRvSenL
qfaEld6KjuexsQea7wda3jp5zsCWz/coPjjJfD4vQlNNb9AlBARI4op8Jwa7P/MwS60r4Wg9m12h
t1pii+dFu4MqesCb+AHt4N1j5NBDRG24FjCd65pzeQKyiIqRtBi7cuWWnOy9zGjdsymfiLIu+iE+
2VUZKRnyAMdVYyJldne2TxJrZNS+ZPW82BEHRyOiD3ll9wXMSBkcRVarFLErq7mPtrONR3LGOBWm
eiVNoksvkZCfIcXFmybt4axG7eZz42Zcv9ROfTY5VlzGlwHInf4l1VPXZrIQKDfNsitWWbdZwnWw
kzGqAP31R6lkC8n11eIgwo+z8N0jRmzl+rfxVaIo2ZWwmcCOM1hl5XnkOIsalRtn6i08fQO6fUOr
d00Ui3Z+UwHVlmZgP1vX+DXccezOX5zFdM4oM2AkfYfMTslo436WbTYWZIHx37p5z8eahl+bF+1i
2hfsS49xwoBEcKbl+m4z7crV3Nd7QSRKN6AFQEK73NCzFRNpkwd93bHEwBoEQ9R6TntoT9VyHmHl
/LVKnW9Kj9DXHLTS6BuKVCF8HEUMx7Q444XQ4aAadWCLWN6BMVjDKGEN87f6J9ek2sJdtsRC2SmI
kcwTcmENzHSrv98fBtfBI+CJGWS8iFCq3VMba8IPyQjKv9IOjOAwV9vTOZd6scVaTlVJQQi1/L8d
tJxDB4ZrMfkskR2YCD8G1dldy8zLopcSO7vGN5QawsrbTqUrNmkmNl8ifEUsYHpZC1L/fe/ysmdM
5ZkbS8S55kKZBXF12fZMxTSJ38xFFNTlLSByBpKIPW/4ssHLpkIflaHxmHnrvuhLFzqW36j1+DQO
WV3T/zAX/wKPt3+AkeI7ExJlmk0aVSZiDzUJQPLbPqQha8nxQrGhdrzzzQ1c4jOHh/c0izozBhOO
GqNOlRYQA00qmsbwDHug6lbxUeYUxa4s0XkDaXH0UFGSthjBhRAyUDtLdSOvgEjzLRDd186Uo1+X
tAqtAWubIGdzlcX3FMLPtLIj6pFO/RZNgFauWViZW5r/voyJ0ChTozfbcQmxiQTBxuLXmv0Mq1IM
7Faz5Ayfas3SDS9mX9lebkQbHIj4s+ycciEl4u+6KVosIztFUDAgIHoHGdB0z9msgrlXhw6t2NOz
OQLdB2uOgE03qeaYfDPqm5HcI5bJzJr2/ltX1Zioe6Vg7rd1g7djp4fHzbSaHkB8BSVpqyusouPv
1JAr8DkPy0FU6REBndn/BH3Xko4UEtiXWa9nieWA63WSSWPhHKr09nTD4y7qaSQvnuczbHiAQjO8
lNnwUbbeiRymvYFtA0OTV6J05AFvwQwNiU147ZVixlkfxvGh1vfSWtjnzcRP8BYF41BYeyjOGDxJ
Se5sGaBPq8ik7B6Lxsiuk1gwG4LmiEpWCsxeyrIRrjXJ+Rd3sKrsVu2iNnewRMzjzbGmwK/2Y6Xa
2I8tw7AY0FuIQchSKhbxAwAI3P4O/jtnbZx961JbAKWbiBz2m3ymcG/7ImRxWV70fZl6jzQzlrIN
DMqXHOy0rzVkSLjJvPbBBpAkt6vg7SzpUDqtxN9PJFtEGEEo1eMsaCL4RNcrFC5dSgzwS3wNq/Kz
B2smGgdw/3ERzWsoLi+GhNvXwPjxVCmxvd/ujEX32sMhcfUwzSfuCqNUMudSOgZK3yoGBYvNHeoc
GGiXcFB3qD7GAjRQaUM9V/a2A1caAETzXHmGjzuxisiX3j1vauI1JF3J9MQZiGZby7A0VLXjbHFL
UpswDKOnl2vK6dsYz2SrCNIi5H3G+CPDWG2l9geoCKCvUiIYOWSvOI2VGokMUqc2uHSCSYawA10P
hx35LLMcQzEy5YqZqQIJ5B1opOMmrliELVDrLIAJ3SPWciJZMV/zUFNirJZK6tje0FPF4fkd+akQ
eaYfkll8V/gc8/gxdIXeWu42h8hpo0aO+UL1m7sEX7fWKuhTLyUMhl0tSkHD3Q9yRloOri421L5g
/G+4t/Ha2CqfTQvHwsG4AiHiz6rPe4Hns9UZgsoY65h9JiITPOg2yAThy7vrNrzD9R+H1LooKjlC
GGDKB/1GP65oh0dCM/+S3AtfntAKAExkN//UnsSXwlWqnoAbRlYFxOtsNr0dMxUsKz5YlByMvui0
rP7WW7/xRfhTSns6m8M5v4Zg5jAGihD8/wEZ96jqTExjSx04+f2yhT9gjlQQRrqJysxi5nsxCiGR
4tV0DJgr4bfHTsJEw586na4yCuWL4lj2zqYZVD0HLlJEniPDFpE+3z0jGt7lSi6DlzYRZbyjnUbW
aYl0tdzcOB9aAOvzaNr8jUPhtgotC87kig3JaAHCXHRZpfHFYXCX/WlyCqsrsDReJu9IKP93ejlF
2tt0xKUdHSzgPDLMjEukoAsSA2f4uNITrw9GXXf6zr3LhHBXQrzhviOA5jwxj8t+fOKnldmNazKp
czNPxmArNYRDXWl5R1bhXNIpQU1uncJpLARmNa2+r4u8NKfdHx2F1EB78A43aJz8F5a5X82xyB6s
qHDaG9UheoHUgBbbVyuO27xS4kzhleBsh+jx6tjCX9o2aq8kMhTzyiuFJe5WpzTmlE2la+BhJ8pf
40cq2tCp/EIgoBml/ATSS3+l8HU3muNJKdWvOG2ESqM0Gt0ktw8uqRo0x/L9rRK2LbbBlwuIbnGI
jyjX+kpkn35fqfuEtHWhH56T1MtwP8YGTsI+IM9O3xfIQayukIW+3Q/U1beJtqt0c46cVbtaoZRY
fGIuv03DHmb+hKrCk2gCPhSHX6dsxglfbmhhE9RFi0QIfFgO1W3zGnHhry3D4oDruKoDH+4W5aU7
kNIDc70dTM54ZZU2YvZBMlqaHOeMJkeTqLpfnaPlIQ2d2WEsSKaqtEYpPdklREJDEy41DbP12hKz
PWgLAgGmr3LlwpC+wzL2tHH61mxOiv7ohgWdEp5u/gsa5xPE1RodPC0G8IPytuQ5fjCw1hyQpY03
Xn3CpojzUHz1myh2kYKKeaRkEwO3+FPNVXTmV3xiKjVyzl9Jlk5tmfprTTEuxn5TwxzjM/SI8C5Y
QyvKOVxyguk6neGevNZh41MzzNY84v1uDkl7RVFQiCZbuyqv6FpLyC39hiDzx7cSlxlbQIC78JN6
Kd/Z1myuvPQDDjoQfjEwV6gIvfcqQFg/LUJtYJbuxKqY4tbqDsWFlGsyW75UUgpDLt+YVu7P+/16
/Ctnba1orO0mVjluCmvWJmmWCGMRxKjODibMvnmdH0v9PgqORdMH430eshTB5x6qKBTEnI2BW95Q
+bH4JhZO94YP7dzf+Is7dcyD2nl5AK/2D5Cz4DV0dxOI2mbaZ2OylcIyymDCI/65j8N1V2PwttcA
UWZuyI1DYmmk+LXLF5tHpj0KqraLXKXnXZYfu4L7Jdpb0lv4NkSshu6yKHI0Ybbt4g6Q6PP1+v/I
bclvT0YirHNEAVz/YhiB64p+jxDEMWfnkaIcrU1ATdaFmdq5NiMhSXGhBdZ/dQhs/RqxMqhkDc04
52BkF3V0PGrY91hwBQ7OIgsHkupUs8Q1ak48ms4rOgzeDpKYxiaPnC+Cd3btnM8R4c05V8FbsEef
BGxd3kkTeusuRl8Tm6gFv/i19N/QLlblCFeJ7+1r/05iO2Xf/S/sK+1czyQctOwl+T1hAXpUa9VD
pLq/PhzSp/HVnZvqc9p9nc7P5ZX058vv26CF05H+faJOjdLA7hnzoxnj28jw6q+V5TeUrj8B7JwP
n4q6EVWn0uPTUenB0OjVJ3hTGX1O2fZmRaErGvt+vziqRtdw4kiowUbtXU59/psl9XLz4/lKpDwX
xSJg7vzI7g1O8RMWh7O6lMP5GjTjfzxZROr84YBQj3LJzDAlTohVKu5uTCk9RG0S/0TT3sCMKbnf
7fS8iZf3KcUiBzfzUG6Jt1zzVXG54jEgqULwOPg3Je+wqM7t54TeXy7H4hdxSpbxbVMP2Chd3rId
T2xqRcABfVf1M+k7abfnNrnlnyFjNXmHwvj5uw8Rzd+GzkSyHycU5mkmsbuxdQ2PUan8AZfTs4jj
RQ0pYb7+ij9Pa7l9DA9/XHBl5LkafEyDzvv+v3NvM4NYmbVeoiz4Pt3l9lWRtEwTOX1PZEh3KoAE
P9wjNyhvvPxb1LFz+bOaIT0gkKoztr5oUMijjgTIWqqQCS/bEjwfE7lAHpylPgw6kcoxXCo1picC
eagR4oQHjk3UiDwkfaMxuQ2UpO7BTqei8XhBKO5+a3NbDpNdvUbNT1YDIigISvjzNC5VceoDZBFm
6v0tmmUc2KvSnH5NTbeTJPMBqMMsU1mzSKPJIvR47jHgfY38XXf/OskgzeIYWl0mA+I3mtL7gfI1
3XDvzAsANPN9X1dbMiwKud0S9ZyLne+m/n5JKq+8aNNA4/2o7IeuPxCdVymV8WsWKUTeLeuZW9OH
KlMOJjqqkFwL+LHLmsPYPFXMUReuGvu3Oz6HPAChEk4StgHDadqIDyjy63aV/LTFwyQQixeYPSDN
FomuOjiuagNv7Y5n05+YNYMyxt2tv+gsAd1FNpc9C0yoM7QcqGLqras//C//TuVnUV/ej+G9740v
29D8mw0q33rwFwNiYDMOqxSQv05LvLEpsEK8vts+Ktuy+/ax6G6tB4P4Hjhffd3I1uIbffnivaEJ
HJqO9OFOmlL5FbVx1CVNXwMFbKzd87nvBMl9Dm87uteRhDhUA2eb1bUtOXg5kt2D0ktZtRIpQgRT
3Ztdy0ckPXWXvVVyqOo/WLlH28eT0zYXCLhTi5B1S9Z638ZK87ou6yCZSRG5HE0Myu9hLQJvQ5Su
mLkQMEa49orTrWG8es04MIwGVEcdMM8dpDnc2iDa7NzcZmNlISOrbk/PCHH/u5b3CsPveny3rNYc
EzDNWsvdODHyg2y7Q5DW+nnXhZgM8ROfGQiWgLscqxniBNYiqU9GZ7Yq5IdYt3N39goeUuzFfzKn
+DvjYJky+kUy0kwy8IsaqwtaLlU6H51FwqsjM9y1CycRiACOJDfMrdUiAZf5l+RYfcQuQhoC5+me
f8FmdxNxCxN89wH/tXiprF5dzVS1fWu7hBGVhZE7NzImWw2LicoP1YGL6Y+mMOR0HsXQZBNyESDq
jXgMWxtkISaV8N3alp5wpbraC24cux+n23Psg1TazPCNJ5EqXSHtadOTpCvjqh67OEzGPfJhrD8l
yJFcNd2PXVaIlsPwHQEsEgqmsMoCer8y4eC3Q2eZfQ0/rGEEgbcQTT0/Ft2lp+6R8oHWtdxvc/il
qCg05oNhR28DM/ydbZ7bXcIwumkjFcQWVS+D1eu5laow7fhsuJXWq1HD+vqIJ90R9Kp7hY3WkJVa
oahKx5zXCbBZw0TdU1w+RIm4V5s8zBdEruS3/T25YkRHSzAv8S2JZBlTkBjMjkeraGaR3RVnSlyq
kCZXTGylIndNV2N2+0ysWoovMTmrNT9Vyytf/1LUpLI0ewLfpEwOgYJuRVPzTTLdhogWeNRSzWcn
7HnkvH6QTbX1VLkz7oeDO9aETkm7sb7VbbQFCrMz9P4t0BTamfRa1IE6EbTc/4SdAhS1/bN/fSPj
Cp871q15OSrFqIgO4vXFTjU+9hJILHzGE0WdWUMmQlJHMZYEjO+hk5DelXgiO6wK26Ja4q8+eeZa
n6smK37UyxEUxZOUg4Q8HsgXoNY753pvGny8j/qx/fTyMVMmJr34K3EPuhiAgtJgQhM1dXtz2AQ0
Whpn5xYeTdZB0FeFoO108BlzPkajY9PwBwl7qzK+DEFEuzNB/i93xbdX1NXSPN0diLZ9AQbB9Yhc
JwWyWf9uODW5YwAODutWON0cV39Qm8RXB76a9qo4j5e55uEYUN/lPYvC06w73pkUsHOjqiP3qeWM
II3DLlM4C5sCA7+lJcGDYvK1FZ7n4JYwJKij5DqRAnYgk6WG5S8v05TArb8DhAitri/dJv2OKJh7
yrKIHFM80n/+fz/xqo2OGsjO6rW1HpVjwCY+XtXgwwIuidy+yIwm26u3DG5cJFfZdvwXooK7yT2t
ezHxiXxCsC4opn+1SGYZNjgjZC72LOuBPW+rJCS2KC/PaHzPB4vPw2+9d06XO67Q+a8CBckMzulP
5thUkUboETtnmMTq8CJjIt0ttiBB0i6grhZdW8G72jLk/N3Uq0X2V6JmGwGeL9Ipc+aPvoPtgaT2
fPekSMCJ6t62XzCrnbJqAmTKgVyjKfN8WMC5TcvsTaukergMJGGyjLzywi4Y10gANVjG/4BWn8G2
1K+TuqI57nkhu8v6ZGjGm7d6cxnARg0G5/sdfG5JAipQ+FYO6TCcRavCKAIgGmgNP1+CTxKBoyGO
afWiYkJW4D9lc2CQrtY9ANPs7jIcQ2nxywqS89Z15BoSVdgAqqwjdUtOuu8r6Jj8ssiysHeoVV6k
SLaOWe0OPZzGVQDrqXmqkCr3i6vk2n44Gs/ORRR97aIAtgSc79XThFA+JwwZp2LFTWsWLHozQGhv
I2lMiU0YV4fjtSXWfsmGSkTeuVD95janNyMLCCG8/38k8BFLdjdGZzO/6U6AP9KKltqAPXmHYxlT
y73ZAUqI6JP5vO+jWGt8FlN+QTBh0JVNci+xbtlGoJWEXYBKF8BoseI24dK552wBwQICBHz4uxTK
iCvnsOPaH3uEYwSQ6teXqfVtwPTHplKbiXGCCjI9/8N+2Emj8P0FB+7sEMDpS6ELIUDM/kB0DHde
gfejb3QSKhLm3yNvMhtxeVblZ/TIXZxGdAUYTP5qZqdPkhdV6rQDwCleUmJTvbTYJY9Huz/vb+L7
CzCGAyrO2bMkGy9XzyMDq2c9IqkZXTu1w8IWwfwswb7a7qqCYPTbY8GhqXCPMDg/UFo2p0cjc0ql
6PGiaQla2imr0rqebBBmFVWnqL3Iy9lnxH206NauvwUrtQATpePoIdPJDnv8D8LRe2hSDrpYuFtF
UoJTLMK30bQiBUvTPr0n+Tr8FGt/uwk4iU+Mf13FPtFgW6FBHAO4pp3hPN1vdoyBgiqb+Qs02oWp
TQo/DUzwPoymDLlj8r6/cRYxE8UOvshuv7Qle6kJ2/ObyAx5cnXPc4p254Qg0AbUOt98lC4f4Gb/
Juq5lSjkvAnnIYWxqOTktkI/tDmDsuZOHZSQktkltPRtWXQY8aB39BkAsspBrpqd0a7aRpZiFGZG
pRxaiAg4hn6QAD7z8YdD5BPxxqFvz4fYysQVWoD+CciQPz/2ZlKGUe2CRrHatAupGYhK2zVuoSlw
PF5zglkd13lmlGjErZ3pSwNytvhHBEQrhEL3T9R/MFIKtxbwqHwz6dRiXXCB9wQE5IevZfj9zUl8
i/SyYulkpu+4bDTs074Z2zCBjxmamfZyV5fef4xPsqaMVYxkEx4BZurMvZrFsmqe8Xm56AwPMA9z
735Dd9n3bAZFQYZ2OhC6ORIII2AHV3RH5HG06cU/W3OfsBeWxi2gFJYxZq/C8hmxWfGeRLf0cftx
oBXPh+ttXo2ixVbH+rN9WAhv4YSSFtxisUwDA4Tnuc+XtkbEGVWk4PPlEjoSc0SBTzPVjdQqg7K7
NsMPsFLR4JFWWfOUC2bcmgVOoeIxn32o/ZfaCP6FeZnrlbGHXIg2WqTNmihsJA51W9ivD8YLxL2L
ojqRpBQM/sQgskFSpLF9CaDa02QHMQIIv2i0P7kOzB16tyRrJAg272fdgR+hf31CsPpbTsww1wln
/xGcKdKfFXJXa42uQsbS6nIPDhazxqo4MaeFQg4O2qQjW68RD+inPgE+RBfzUOiH5sdSlXd5m7yS
1LsItCqy/ceVq64lkFCdt5OEHZEYNU9uIlN/7l3ODj96rLsqXqeYkZmsfDvOhLiSlJ6m4mpyCkPq
e9/8euiM9qN4YH5bK2PJV4gVPO+Ara22FChBmJKEw2aWAcwsXLv0nvv3kFlHTS1reSI53XnKZix6
Eki8r40ieO6NYuolMWUEPjNheXqCVB2iSoeT8s+7gGXNX7DHLb1RZlHHI6pSFvjZl5l6+iJD7oZ8
Zcgb+8vA+VGDKj/EPC8eVUCC6fprVMsa2LK5SGjFrH4c9EwIW+AMoE0m6P41cvD7cGuuMjgBJqhu
oLUon7mVGuS69JXyed7FtPSUlMFaJPgnlvmfOnbXwDWGcZ2gkp8kVTzRL6yTlo/xAyDXXf9r/ii9
HzYUKpwTDJUE1Ju8Dpy5kBXKnoZLSjVmRwStWx4UImApWowJYOLhXbNYZDtQORTgm1UwqiGjCy0o
PX/dEr0wyIfTWwcCe1Wa5VSmRKYP35f3denyAwhImQBmUs4tECGJi0Zi/prOxthWHjeUXikFY5Yi
jgBCCK8YdFipCnLN4T6R2GI9MPH1ZMcrSjnyEtkA/rxHHt2cUa+oqs9UVHCb1hQIIld1kmXCIGOj
n+Jdr8cbEKAXQHlsR8RDgmAd3GHUVA5tmG9z9tQO8+gw87kB8zjV3zUfFtkEsyJ2hrEMV4BhZr6B
Icu3IoErshTL4kCDTtKyLn+7EPaC4z4+vR+ZF4eGAXyBcwduNu8+wNgyreRSJjTRmRTX3hXJvx3u
RSzRxkQqujZ+aygmrYRVrVkQ3AVLr/nqMWQRjktsBYl82d2Ju9Y4GOMKRmCEtkhf4vJgdmmViuXm
DdnNcjgWdKnHLJ1hRuDnpsuw62Mz+xFZqzAoZboFsGGZgnjY5w5XNvLTZ51L2OBt6ItduZndYPYo
zyno0ktxdlw7rD/JPvE1cbsYBKwu8qwpmJecopsxK7/CZNoFxUgBxbQdklTGPsmKZHbRaOaHAbkn
FxzFOvCIWIe20+X9gNp7UVjMt6klyUJc4fyRRs8jbhlNBNbYZ4gRTwECtV7fWWUJ8h8iWRlQEBni
sRAtSpIGXtPgIhAJIoxJSu+3sSGmI2KTNz2Op2xNkXyU95pPB8pf21Rw2cIDHDiqDUTPjylyMK8D
S8u6L96mpBmVCMILhMVIW2pUaqzBSO6nKRGat+nlYo1lkjogy6oZ1FIvh4UAh+WDvMKMKXqb4ice
1WHV4kX3yk5z9r1jG7wDCFtoc/Q3JyYkMsybheYBGx4eN4jh6QoboKjB8DmLPWlk9hNA4usON5Xl
F5DaNXOakf2jYB4ZaNohlYJv2FKz99aIuTa266OX2ZlPFV47Tv8lGx/ZykO5V4fEvrT81oShMZBI
e9fhICfGm5YsomBb4bYtz+DvFZNDyD9jsTwQOD+szwAYMwlnAB0FH8vBlIOvMb6tjDg1OBfq4vD+
r5hFQZ1hkSYI4HsaIQjdZPUvSchODUJ3qYnsuv4zQpfB+R3vs0mtTXuVnTr9MRd+MhYMan/i4hVy
O9jkgFRGTByCaiGPmaX/6KK9Ct1Tjn9nW1Sh29EdltvfC7jfcfCnhnVimxFTna4ibowy9FbPu/3n
LYd3BWSYdpWiD1NrfUqxlZ0d75wZc/btKWAzqSiF5fRIZ673A6MV7e4mqKgyzNdB7IxZb6X/HWGh
sAI84lER+tV/Psg8j3LMgVcPlrODUHzoDy+uh01qNLLrF3W9ZvInsK15ROmiT17YQNHFFsCHbJjn
cINq9zcUuYjOe/lPdACOyc4G0cBjjnxwR+6BTXqpaxGJ6c2afTmMMPCdbJ0Rrv6ZVlgbzmGAMn/W
oX/FroDW/up7rUMIOnfgs35hnkd8XEiiPHIfEaTQaHkWTPyPrMOPz8O9Wti+LSOhXYKyxLhRPWzP
brcVS6d++ptNUa/VstgBfMxOZATsMEgy3EThfc7KFXQW/6dd+hbW1ikccuJuhtcmtUq4L/eHz6wL
4h2Eny5uEIGOizLeSfvlJe/wzr7Bkykhd6wLJIWunxOcXebJaALbGUIU2jH8DE6iJYcjsIzYdvVy
DAK84WiXkbph3HKW90HbQgVvSyFhCNcj8k0amm+GC8o/MbWfLfGyauPPJj+X4jGdivgtqpAWMFoi
dVpBfgsDBn6Rhn6IxbxTOpd8NoerJ5XNAAEaHgumMovjARpm477nQ52g0dX1ThyHCuGs6XFYRuN9
GZoPi7oNTkJHvYKsdHyc0N8vsPnJmZD6TMaPBPbI1BTmqEmrqEOS79fzyJd/zrAhhpAiYVBZFtE6
lP7aEcbPwL8HkoVn/HeAB96HLn8R9BpiDZh/ZD0AdwptMxwljYYfeME33VArQOUZSfXFsUUvMcLG
qqkk6OV8G5uYUtxyfKN4Se1LPSPbmx/XpVWJ3LCv+zQKAlGioUvQLSxeVX1j3aeCfNrj2/3WVMWf
TFtafsR81MR2oPGRuIm14wg9dJ/EG7IFrViWrkbh8FfjrYioxqyM/Wn3Na5Oi/CSiyC8TRMJ8IHQ
C71Ztx9l6dIzQFwRwJgJiEy6N6UZxD75yqRfd6qzQUgc8bD+23PdAH25oEVBwjvVj2xr+lqaZ6ty
4opNU4/0vZsJZQ51cpzLnUyN5bBVG1PA8eQThTF72ygOO5mDaJ/A7pdcXiQWMaL2sZvAmrblFmkl
YkYc/MpU9ftg4rA/ZPV9dlzY61iixuqFaI8V83bn955IMdKJyV3FDM+CEkzicYHKdZYUS+Z94OR6
DlJhSprSvtDdTe0YsTIreWPj4d2klGXPSWessaLLLOJWjSuSRKddt+8d6IO8rsDdo1TNWxe4LSXR
8L2Kzl5K4hcOLl2xZAnXnyVZD8jKOTA5/hEcw3s6IpKzP0WXDUw5d86H76iho4chUrB9T2idk9Cb
2nDEP6adLVVSMFPwXOSa/aMEM8Be2cMZIwunrfY11TXLLku+krGXq4tRUm7a7HRXthpo0bjo4TJg
IA3rS/tn0L8U2u5IO7cl7JspbISR4U3+KP73wCQH72ppjMGwpIkt2A51Ul2viuEVpf6Ycc/qofS7
jFdTdqs1Iw8nr0neZGrTfnLLxnd+fHkNsu/XL0aowLfpV+QPZpkPJOU1Fi/gXh1BThVT6ae7mtPc
Ce6nNjPcgwvG9xXp5sFmOfPg/Uk2tJaTPCh2yKMjdJV+BvEHR/nRu9VnwEMZmri25FCYJhpT3fBq
T2BiA9BqkVjvgFUNZq8MG1vVOA6BqOERYs1p+eozPzS+tVDSD1DzJo6HwMR+JNDc+sG8RCHpLg20
JJlC8eish02lz7ZG529YhpWiCeBl+dRSMUBaUiuhWqtqDhGpsDWGITtaIJPr2dzgaJoOPsnDV6Ay
sKfG1nYLlI57zOu0tXQjIliCg/msHbtRO87zHn6JwhW9GDh0nuTw1u6H4HXCg4Xn/2mftGVCVkYQ
xTBBioCbvfBD39aKImLl2wm66Db1Xd8RenYu//V4kCBKEXJJre4iculMzBEoFJ21eSuazDNic7N3
D3EkNzaDSW8Qmucshr+J2azD7jRT1+V2ZSn8qw0+4Ez5KxMTrB/T6zFVfndm9OEW+ruGPucY9UHA
/azdTrZmprgqLM3NDdCoFeBUbpQYAhosjmIj5nrzT3UgT1D82jhOAORRQwMGgkrUnrnoID30cIos
V9tFIpgtFGMJIwj1zrgyu1Gzj4vhfW6Xx4LeqEY5v6xPWk3HeXHq4AiB62N4qNOAXsgiJy5v126H
58LVO9dE7sxOV97LPe+Xe2k/kwtO+Rja5nNF3Shl7glACY2x3bw0o06W2xhe7IhzU22b3uqiuL/i
3uH+WLQPD15Gu2/Nqhz5RuIxcF1dl+e328YviPuM03ZJKrLdI9D/VaRwLjLYgnPa7XLGLCeq77Rv
bhWZ0eTpnbSJ5Uzgi79vZzMW8vRbTsb1y4H1uz3Qc/oKRKG9PNTHk6NgInEfI+FApJmsax8z4xln
vaQ9rNujKZfETlF2d7ezrfcHZNOy2tnTViU3s4AXxo5oXQ4KgtV2WM6FJSh2GukwhC8aT7DSBfQX
uY8es2QvrWXaao/Phky5f0DZJVYHmR4yr8C2fMR3CbUfRzw38fO4IbsymocBG4JuDj7/4D6Felq1
0EsQ7lTlq7Kqpr/kcPWSzIi0wY4vvzT0QAhfXinH+oGV1wfi8Ak/Cwbr9JcszkhEm+v04QLI4USF
mZg8TSTPAPu8VjG/UaUcOs+8QltaGk5r/5OrVKoWwEY+DGWhsdKHqy25cQgBymX036iLQNKoOHdF
SFasOBj6ObsVmIpciFxVnFfS1gwLWySW3A5tCwiCvkKkMi20lSaVI9k/jR8s9+EWiuuUh2FcP6hd
FHQHB0ywaC1Wa8v4lTcwni5vCsFqfT/9Ga8HViIcBv+BsIr3XT2bexOkNw5PZ2Z9SC3MGIMTF8zr
sPuOndPEjZgx6StVXrdfuIZdKesWet3+7Ho7JjAt9/G5qNQ4Tos7Uydd4W8tjFzU4a5/R3xE0oX1
vYFmI4l8QMopS4XoBeR5pAJezp/Z2lV8Uxsb7i7zv7VsQSzryuPsvATevkeGVNbsVgrc+1gtFuIB
DJACKH8OKUlvPitjnBf6M8B6izbxYOySI63ED3E10s/a7F97FaIafny8usvIRqrgU62siP213gk9
W1LozL1+44bHPzx8SH6d+MMYAx8ahtKvLoWRraMY+X5JBq8TnwsZ3mKoKjK983YATT8723hiPvZu
xvOgtc7IFv/AefTyDdRJ77tbpOu7Buk6ZiwT0BF1eIZWgzCsT8y6esoRg9sSdz+UMV74+ifVHgSY
Q6iP8uKwBEAeUD3RfCkZy9bdmS2KoJ6LyxmUvnziOvvq/OG72P2roUI1Ze6Uoh7UBG8ZaFK+4VdZ
E5+6CZZv51KHze48zPvY1COZii4TpJXK0nW6GoEOTqAj68IgfYtt5AU46bogg2x+DFszpn4I1v2h
4svsgZFSxpiqU2u0GFiQVgBBsgZkcNy+j7XSFkPQjlBZ9MNBM5q5DsAAQazjwsq33oghdJzE5/bO
TLsDyNJrEd7Vjcz6lhuFhR7UESmsL/kx5rkcmFLhlKdodyb7eSkYF3M/gGqAtHIvsQJz5KaMMIp2
0nhs1JTRKvJY4VSMZsOh9O8RZGqGZoBoeRRpnrz6GompW6tsz4vePBLk+yYFjXV9T7Ggi7uARhOh
8OTlXlE28k7fY4tEMVIWtOMXhiPiGsJjz6A5maH7BaCMWbllGbYQ2ze/cXE3fUQLZSrKvQb5iH17
OvGDNoWZIVJeDCBJ0Mb/5QySjCf9jThgOx5qeZx7EPlD0dmUIp3sXJXuV3RXGN57BRA6OE1bnl5D
ctgobCZu+Z0nQYcmr3srYuwuv/vO6snNECJLOxiIMVq5BaLqmPCQCtbj+imiQtd5omwNXjymNiFd
tIBcOSlx0TtUG46d4ptR4ZFsJrr9/WiHTxthnmCiTKUx0MG9cQfBGU7gyKPwPhZPN+7cbTnxVtyQ
dCU+yIjQYyMhEJTYB8Xz14sH6Q1JVN1YyDW0Vpr7EVBArKpV8CVD8q/zhUZAh4VWBspmVmpgTUoc
H0hGmB9sU4gUlE1RxO6sE6eDggBtQ9AZbAHOvAGeK6NPt/ci9pKlqEaRJlyKdfQ4/hG/rl7BpqIP
JU+3sPXnooNpWLvc1rbBOFuaH4X20JnezTY/V8cu0R27q2yDXFihqAkyFcyUXpjrsj6VSik4RGQI
QMP4HgQpW58gJk7jxhrPz4UYsYTw6lNFfXihgeJLOBqs03n+ASmNF36bTtPsH+REEujUd9M1u5q4
xPyfBC75NHWoVi/rGdNqv4yYoybhfSn7ohYWhVCBmrqYVNJu0O2pQptBS0Ks6TDM7Bf8rIddPt07
3qlu+1PxC2QVgg81zBD2UwA+AKmdovsNZhUnkI4B0DdPtqUdxweKKeUjdmUVv06try++gWu7lCrT
VgMi3/zd5eBRh/R7arWsaqfuCoqZLaPolLGxdhDEuo/DIephqJ0vZLRVjtEQ8pQPpz2XYR01xCQP
qjJYbNnWPkXegTMptPXwGwbe+4a0G+tjcVYDpXqRdvlnMNJ+h6s0pniImJEmhq7ZD9FRVCaSxbM9
rmBM6Qdc1MUv+Csd1bEDVwfkO/Ti1mVU0t2++UeSK1XjLY9RZpM41knFXjQlptnYL2mInJGZeQWs
jlaeBNwDlB/b164pfyVK5ZrYqubarG8lPbtXPyW8MMG1IP3csYl7E1S0gP9NSYbhxuJOYx3YrqUZ
k3hcSIAjWy7qf/wcSvNk0aKey5UB7nHWSnld1mfjty1cs9i5xENmrDadlqpSEbrXR/k2Oczi5fMv
SShVkJ5G45I0RUFE2jxU9tTnfZbD1Plxx0xy9Mg3GAMMBnXcmUPBhC2fQaHcCUTv2JcQNhSTBQo9
wj/rYM9ujs6zXx7iAWLQrc6PaOu3zB+SZXZ0TZHBfCzgmAGhbLOZsKgh5Iiue1p1L1xfXtfTUlut
13BgKE8sRuUu0kLhIn6J9O7NBptsI0cK7E79P/XUzvctQ3p4UTeSOjrVV01pLwaCOdlb9IQQuJ3D
XtdkVgKEIVkB01L1jGk7/u3craSfYzdWmJcwmCdzJHgK+vFRrsReyMeRQnXEJafojxZ0zFPGB7jT
zxDAze091qT/DB2ecSJ6sAhp6/ro8gfwI9llIjR6AJPQeyErc8yGblvMtf7qwV5hKKx3corHg+Jj
KsIdEcPrakIc2rtGMnRfOx49EeRwWr1MsQX91OXm4N3ABV/dm2Ymv/eCO6rUm4fM43dzrELwmoLg
YTpQLccMqwmN4Ddp5vz6ykPmOek28nj/8anOTyK+CmR39s2bVJDdJjkZ4PANsqud/treIibQK0U4
8A3XGhHL3C4xs8caLONeFGDY7dMnh9MNpxL27uPnAcAfdAs7HTJnXDxVh5t4SKfv5gXF1XfBQMJL
H1x6G3CcTFjnixW3kFYJnaje9xlNwp+4HmIl7m5cPGSAIJhND+WAiGplNB/2RtByiOT+jFBEFdZm
C+r43npzV+fTFf9WI8j2Qp3DT0XYkh8p5u2jTYbRmEtHevOrVZHMh6xwPDQnNdHxf41Z6Lr1xuV1
wr7mJf5/wpupRTTc0z84gtS54lXybxD9Wsq5Prqbba3gNac+8TSSEDhnn1nQgzo1gZt6BI0TupGd
qm8Lwnt4uliZOHHGy1iNAWQDdOnNR3DWnmPJm0uk0hxsEunHeBefiuR1kPrhettt3PvLJ2DwoZ6q
+k9+A2xbrF05/Qr66h4pRsuGaj4TROi+re64UeEiPCgQd46vZZR4524uZ59+eCKFU03TgvfOMPXk
vIAGUSJGHRIxCSCVGKyFMZHjquWd+E2IgKwlfB2txnXc6YZbQf5r2gSCywOeNcv0P2Jy4BJtprkS
zYVrmYNjdqgv4fvlfUiwdEGgXl0G6/w8ywIkzSQYbyAyNdgY040LRZLHY2/9UGXgogSNfL7VP2Y8
BH0M6OXkgEvBHJiLc4i9drW43Y/VrTMZb7SHMiy0hhXY+x3QDIn92u7FHj+Lv2uWxCDOa3ezxLGY
XwF64xdyCFeV7QdKaPcvyk1r8hXcf4UeB76if7/ULmj2874TpEWQLWUbSocCjoVS81XHuwdiZr2K
NkLuQ9Zy0b+HKJEyu5TeWhy3yPHxxzNgE7HLXZEUS9940uFc+kJ+IhMrcOtj22UTH5KKV83cI8tL
YSs9B8XxrtVEeGRRjHQhxnWPfnxmIaC3rkie2ozyxIExR7H7pPjLcV+ScT5nJn5x1/FsQAEAdTF8
wCQpSpsTrdfhHucJm3S0FGq+7w7vXiXEfganrNnLKTplYQAgGyQM07sOXP1y4fY3un2Vvh0/6Kpz
ZQVDqD8V2FQ6DdNDB7z+nbab3b5mad+9nXayxXoZZcfmUbm1XGdDZ8o//ddPChaubWo2/Kj6wvRL
FxnVqu2tvmoeUR+p6x3tnTWuyt4KvH9zDbvC8mDAeOexS52cK5ecSlPpVSVSwGZYck5KlFE6a3D7
5UYZXmMbygFy9roFuKwJhHRKcVkHPH4Kgt+hBN4R0M7CRwhdZCzsQ9gXjaY+OiBfH3uvWQ5+zkSH
/N6R/zKUq8tohj9MBNrXx2gfJW0UW2o9x6BibHaI3VRoOtSw0oVVh1dUyf7TMwpOTuUDx9gFuwak
vi6UAg/reOzJHw6LSRwjn7YqzPW6t1MzbMR9S0kiwm0E98IOX272GtEMN1DMkyAhQJgbrzrbMtE0
jlEkFPYc4us0akxHPxRWCDr/bErqzp/dHuRf0tTFQkrDxWS446IQOLY7PiT8nPcQSzv1QnF9TY+q
bwYpWUAofhrWLsM+EgtreIckPPSABiIiek1w6oc+ubYEDxpn4LMjJseXCTcHfBKBMAavsF2H/5u4
1PJWDl5htvD2J4Zdaxtkg6BBUqThHxFc6XIlYcOCbv9/toDrfXt1KvTCbILfssRxjij9up6QvMf2
dKL8sJmwZ28PETfi1Yp0QuTXooeOeBzXxc0SSqvg1kHcarH2r9MU274QzDI21Zi3wi/Kdki7y4Xr
Pt3YupzGosVVjPnZMHzmqdzTa/18oS2mkj2LAdvaM9409XWhMAbIsYSuQYmM9Ka0GKa5hDImDRzV
g8gnD7KoW4ymdRojJn/UbuhnEqB+fV70piFLn3Z3BHzQCqmvmul39otEmGUY4/g1muxhjpFKCWDw
91bys49UE9fVo+BYJY3pRuM9+bf5ZaRo38vCWbLtCOFrvV0VhsNKDjaa4YF7v3HyXCfIg1uS0Bsy
YyKp6twx2zu2qryxuwJSfO54GE+8sgTvNZs1dzHgOnCr20U63r3I5j2ZEjvxcTdysTtZnQeJUuZ1
MQHtfbnZqzqLBa/ycFFH3ZGcuAnMaSilCzFkFKZ9Y8ZSY24cO1Y6Zc28H6ubE6GbBWRcPmcohLiF
ZwhwSIQkjFmx5o/mH2te+MRL46jhOlxguIzd1knEEbAgMu+LQ+PeJvguTxggJqUB+ZMas5kvA6Ah
qMNlUg7tri8DHlbLtwJ/03p0TGM0tUI/ToLHceMvv5lRqsMZEefqIO+hd23PHfaSPpNomXBJwn80
pXPLFgzWjM87lABwxqdhpAitlu30E6Df82CN01LGi5J/zyM3nZrqIPd+TpmZs+3Qo8yeJOS8FXo+
wpX5vGQxXQNqLZewzjC/l3Bu5SO+CNYCnHoWm7oykG1pjNmbn4ywL59MoDMDGgf2J+SMlImjaXJf
tu2lRJd6WYTEsWVn/kALjsKARqLaK3K6zMLnQDb6qxNsN2BWGXYqlTlSenEsZdbFULCuUhZf6k9w
Zqp2/9IfqQkH1kKGH320ydIdJ6iCAUp4k8kWs9Xy/EgTp3rvXwdd4lUxg1HRMvdDD11dQymgrKYo
gBWQ2Q/jg5Ui36N3Av3GPePW0tnAuxVu1MUTvm1phxsFauYuGKMvvgYthfigwRPWlXdDfpEjVGBb
Ej+FcRQhSeN8ugHLN3hVnci3xwejXEMPl80yD1lDm9X1UykZIK2Qe+/9+3/J5l1nLoZWtnpKqq04
WlCcJzNgrN9lLpYuS2wQIClWdbE/otgM5mJ60ey3mFgH3WBHSgttHMYmIZ9CvEOTWULt6lUJk+58
v72FP6tAxDEQGnIUE30k3tQY+Pp9Ncttm9Vb+F9AbsI/csKFwY18I6bCR8rKgAzPrhvhGk47/hiJ
t1SgrBMu2pQ65kKIHQn31yGKm3ql5uPi20uPrXxTZZqW8EgCXuQYgbNByZazHm2ofb9uIwz1vfms
nUlSiGs720pnZmLsLF8kwUdvvkXtQVwetUhIHHGf6ZwQxcKXGMJfEAitX4bKilVAV9qxhLfZuafo
TybILg4D9Ajm6BFzovfNDy+M3xgxNn4QxPDTZiCuRTOwnpG+k/1Puv2K0sqNM/YEP2Pl20fzw/rD
ZG3ojpQI9O+nGcxlqDfcfIG/oEU3kHfpXsgcOSwzMCP8wqqzXU6zG8tC2+fEvWZNJ4xueDZp8OAq
ZAfVWobfyvA307lCyMGfyF9Hjp577DPU1DHBl6iE/cnoFU8wuLTpt2qyWZR5Y+8czbx96bEDsHSA
tZ8H/9pfksAcQY9OkPvdYwfUXiQYNcZ4E2UxxTZ+md6TPw+YomV+pOFlFj1C8qt58EFfhuBTIhyb
DTldZyu6zpqjmghG+vUvXsd27w7lAm748MTfA78l9bhU0XCExdWxRtyBvKLma0qKwvwZulCGIImM
RGiBmWEAMYnjJTTxbW+w7NiRKaf3nx/CJ3LG/dk9v2RvLRw4VxGn+soAceCOztdT+soEFpZ0zjBI
hcgqfiTEyaeMiORQCZsKszccicwcCTLF+O4TN5iIslv3Udwv3hf2ANookvpKZnFgOgv4UiThKjPc
GwUt0nwxLHnkP4L3KJh9XicfBm9lI4cyOEBt5gBvvC2aI2xcXuFl+Hb+jXW5uKhxvA5YCaFJD0jo
cKimDG9vhYvI32s1kIZTs8xP5Zxducwf8RqbB9lquiY1e7cKf+72AicAtS2K8beNufp6Hl/K49E3
wUfZS91IW1QqcK1iuQu8R7flsoECICM1kJf9P7/6KTO/33f+S10/MIBMKg9gUvkPyw/WpxWrRW5G
5WapewnSYtW6Qd8+qklImDNtUFFeyFM9F7gkD827LFHXVQoqszWxGCjUfxRdwyaVElMqeONSaOBf
Rf54+nDBPTrN+opDZ2VSs2NHZwVa11v+OXgyqeoPuQcQHc/vLDkymdwBFtvSHHbD6syOs0nHel4f
ur2G2lDQ3akNmM12Ee/oIqbhOrKqi92r4SYWHV3NMNDZUS9qDnQEXiRmu24uNsYdJ6x4m+wMJI0D
Xm7IuvRgPtfmOGBalZ1Yd6VXm72LqlGO+AhuOdRQVZy2n+IRXkwHsihYDw8OY+/YnukyL0HoGUGV
wcZlu94B0rqBrCkvV+6/ycW/LwXEpo0RBWX1IIy9WeorwzeDxjoCy8dnjWCczKfnLuT5IFBnIj76
BURbRyAIfKrQPxzzUGkYl6cIxJgkph23sGYHcTtvhIWXYm9HyvLwPZUP8ks3IFtV82v4/LnReG3C
afxNmXzKJhQMsSBfP4j3iDfGwwviiu4zVCpP3IknDmAz7PQEn8izMpX/PCROlvpZlaKdU3zYpejH
CxbFafVP3yjcF1c8TDlgDr7VmrdnU/RIt5gYSbqh1CRgFZsPJtrP3pbShHRxN+3QKBuo1UWv9zu1
Dow8s0sacSMlRbO0ex/TwEh3Pw4WqwmkpAddWyr1J94tOsWKi9VMmMlSQdyjDSNqNc7FAQ5o4YvK
AwB+Kr8TD46b1xdaYSJpzbOcADRMEmcdHMIDTMAkM4FgP8+0cUGmSrejZMJJiHwBhxy+1TBiIrmX
Qu+sTcIiQNStcUx/og2kSj6aZh4/Uh0OY80uomlPkelOeOxDfXb5UyjsYwl7e0ih5wg3kTTTup1U
RCohzdVvLxWSO5xfQ/4TM2Ak5awI3XloBlu3i2M1C53O7QtJAopZOgsjOFWSHZPE3dkMTa0Zefbq
lqyyik7tU55BsaDhCBS9JvRuR/0BuubnDNwOUfQX8UHUdfb68/oNJ3L+OeffWBjKWLoMeQUQPv0l
4ECqwKGGDvT68IxqMFFLKo7HgItOj6S49zLzxP9jyKufdCcggp8Gr7/w4oCq1BA1dvv9E2TA6/6O
ATFWrj4ekc3ruQPTOUWF9a0/A61Pq0de8BCHII+RcrktBTIpXaulg8DmrBHT+0QMiarIREmxtEWJ
vAufVBVSCWIGPz4/IIt3Pz+42wRi6MxtNK3SDW5+bEg+Wr7oYoizFec/Ob40r2xAxRc/SBuhy9Qg
1iEHe6bC+UpXjlW2Fw9rnQE+cYup3gTZPsGOAQAHzeG1AuYuUDvbfx7c3SgxAR9xueNkLGJc26ng
TRnNTlp+q/59bXusxBeSx/a51x3hLTxvbVblNuX+QAmbiAS5t5vBM5dYZyKal3AptyM8/QNFeXrG
nkbm/7JU/yfFYC3w0/c3cvJTPp2cedBAvNboF/tU548w+A3LpAR5oM7Tlv/EfaVzuJCrhm/CABPI
NVmasEYaT27ttLu3Q8N68NELayCm63Alkxgs3QY4i6Yo1/5HQ0iJYxwHZGHiqiQJIlAiTn7DNEwi
YJbBNPGC3zNsuHYKddcOXxQfTH78v8gsSpQHvNaPd3Vi9fHe8+spnybeTVkZnrCCVdUK5Wen5r6M
k5B4WGgv9jwhufqtg3BcL4PuAafZ7o1FoTabVNzVZbw7pSTb0RmN0RZT7ldJgPa9qL9/CEh0k+0S
etpgY6hedko0l89Y8W7Q+A9gIBExzYKTBYzMWtmBNlSvojKRpl1kAgkLUiKbJJMVqWHR36yxRMRM
fknVS7XuTV/EKYOkTF9BpMLYGk1CRKNLTAzmjv9lyRRbH4HK9tDy5FKBn1EamI5Zj7EqZN3FEM2k
TTWDdOLoTrH+LFqyBz08rYngB13c0cqwlNbC/Q741/oCaqaKNC/t5rXe29W0NOIpHkome8+6FRCD
hkolL4SgNgPbyqOoRccnbjMt4BG0d0X7MxRm0huSkNozC3ALv29XDFyioRNyYpoSwOwsSNp1wurD
fTQPCncpo/Jqx3O3m1sKiWZV3orzcaVu4OPeyFbW6hmAVCeoD0+UOMfcBBypJUP5nqI0nmHDviMY
ITg/BS9Ubp9N8Q+I0GANFO9X3dsTvGWdg+WTXh8UYedYpXifQpjHT2yVYn4ynkitvbqIgzCatDS6
gDnaI0lM2eyyf5nBbwaxtZhblk4PP1zas+H5J12YkDE5P/ewj34hWgbg14A0b8bOUMG0CN0mEPdr
5cseN5UQtMrv5mdnEnWxZODvUjk4X/RLQn2qNdTybsD5zdKgwEQam0nIefXuS673MQIMySEcy2TU
4yMgGO5tnzBJ8braLcs8p/3c56I3pYTIsi4OHSvxsvmMXSZwfgw1ES57MqfE5mOVpM6kmtR6jPjI
fXAqhhU4HX/L5G+KGwKmyhpou65G97Pf9bp81nnPWQ1J3o7EVJwlOn+SYIge6YBPpGV9+OowMk2P
go/rK969GctgWWyrIcoYDy9UmbwTvFvBqgUVOK0B0laTYjSbKChec1Hxe7Uf6AIjGOD3hpOn8jOF
kKFo9uKfRYjD1hppSJ68U9X6nQqR7wCSOkBwUX8nRehXg6+19JAJPqBnhviEgTWZS15ReqbBtkSf
QAK45O2Enjb8PLJ6GM+7bgiecVllt4jJyQvygK5E0QsgbbF6uKoErhsogf3P0ETJoAWBcV+gz/fQ
v2TbiHgG6gbvbJhBadUzzqmsh5b5bNEZKE8znd5/TmDF9kDV2brJs6fHBHOud/cPnkKH9mKeh+7g
ZYdDah2byzHV7j0AywuwRaDjw2/m4Wvj0uWGPCsg0PziKoGZfn23XsYQrafa8yEK4+2ccr1LKGzO
Gfuq9nseN+AgSQ/VgdbwD72UibcweS63y+lRLc1MCG4zNCK9pjYoUGERsksFKn61F2OiprWo++dH
BplQACzU5J8MFhYyLxO9hZwsU55ucZ6sdZ1fmPu+zPDUuKyd4bMaAjdRlBhdjZc7LhcR8eTIfq7J
u0Izv98hs1EyaBfcu01cIPaPCScOKXj8HOR3YLJbbiCLDkqeGdwwKSgo+ZMKsoUsteTo1oTMa+Zw
s1cnMflutKEDmg5sIIMaOx9N7qmDeWDlsFlUrFvVGv9/75IVOBqH8XIeEgcT0tht3g6EaUTWiLGx
p33MImeHvcy1dYZtYK0cc+gCcittQ3gXBg0/ohLhbXNN+Do43cIzuQb+w3GKvl436LaPAK7sKJmH
CfZ+caR6xXKIZXwSTiLRsmdHY+Myo34b19/hNfYJ/oeHbxx8/khSy/jWrfZL0W5OgxyFnZ+5jVms
F/RZy5tiwkODq/PK72qS2od2katmzyCM/wLHU/djuLz9fHPhSDufrPVDvSfgmN3QxPAWk6y4UpWI
6eMJzHMexegXaKOBq/aW3Of9YCaOxr16GCaf31b05BvWWkQ1p3Y9mTyPKHrkqZGgo7zVPUM9x0tr
PNBZfAo58SWV8TLQkBih8/A7Bw8vTNLQGsMcd0Iob/mxEMIP77V1Bt/KOPK5vm/qmX+mzWYyTc4C
MXTXPCGz4OK6yVKVCmJre7uRf8VPi27fG6B2M7c3HMdylzPcms6U98hWtEodyMTbHeG149cXZ6dV
bRjI8Mdr4p2c8JcdRUnIoJmSHRbqrfDnHThUWy4oXjVdC0nfkprW0TZg+0lY26y8c1DEakP45yy0
KrDYMQZkyPMGoZEidMVHK2kg5LHa1YLqyGooEi1HiCIyJ9bmrVHbm0tVi3TFH1VOmJ8utKpB7DgO
qEpd8b12Y6cdsigNK9wgMa1xGZW0n0ourZ80uRV3tyr64agnpUMEIX42mK6bYzhcGufsXSPLPHgu
lQomhBOiALcQyL2INWEqD6g4dgXESy/oOYT3+1PP1P4ReOreV/81YaQafJ3EDNEMeBU9Bn8MtST7
eOZPKn/kD+b49hiNGKzD+OKutk2JASNuTlEjivdL3LrBTJtx7Wx6cVG49EBORneTTYQluYyYgkAz
+i1752l/1iNT4QeN079BM3Gi1jxNP0YrFINSUscC3sGfdQATFHRnk/3GUXekd+GTD3E1YRAVgtN8
fnRXw75m6tXcHGTSZXH5bcAQlkLHRvaHSwpTxB33g0Oafc80FTsm+7xmEuBYJldUmiER8042avux
YEPpn+Mhd5ABA1n0Ygvo87YFhjx4b49Ru+h4XPUPNtNRkqk6bonRKiaqNukcwRjxfG+opp8HgI8J
W7KWkgjcTCEJXk6D6Umnxdqd5+CzJz9MwI3g4nXbkOIn4ddBD0GIx8px0jeg6tPwKYGas1HvyOM1
CVKPaMixjy4HgHSbA+PbXHWVUcQrh2t7AdS+sph4qYBcEl2mNoa/Q10IVPjzkS+tdXXw0BwVFsMB
yl+6naF97MlurjYGTe5j2al1HLX0c0g13TUBCRGU09uzvskstP93XK4WXPbyIpNA6b0EVtFXqZce
2ObqY4CwkliX0AcUN1H5e7cTIoA9AffII8DqfNBSvFkHHbxSgGxaqiXgg2CVHr6gcgVjKgkbaEXG
l4UhfO9mZThEkrGt3qO9L0EqQFoA6VME2VH+pwJI6zMc8z9cWvoHo1QaJXC+gkHlA3ShFnB4tJ+K
/eBWYrtRdzVFI9OcGrzZF2uwdUSIlwHdk7FAJML3kt6foSz/CYOgIwwYKrxkYXsIgpj02Yl4Tn/M
z+ayLwPJRN+uWxGMz3gtSH/ctGJULbKSEOUBdP156/QBEKcnY779eVPfRyvQFM8iBPvpc48wDeC2
BS4ByL+HG6D4wFtct7RVdAIkIwiuBbTCaVchFlTK2UtMXAYY3B0dVojTawss4FieMo47m/jwJcKf
OeDRae64lHp31bbN/NZftLrpdX8Gt1LklEr/u2nVhM7S4+h6ZRldAZWn8xT/U48+7Y2i7QeoDrxD
AElp0JnYvCgHswAKYSclcjPlC5VldqAV8eJwr97PFm58rw7FJISZtycCPNT6v4bzEZeX9tOvgN7u
zKN7yj7jgF/qChSeP+I0yEM1oiH74pPvGYZpgPYevZ2zFV2AuwxEqODS1VKs1u/SX6qpm9s0Al9l
7IAa4/Bq6Jw9+wMzm03Qe4mCj9QlLBhcFsMmjAlJ80O4PK1ZHRcE7s4BJvYslImKLQG4BmbXB4/D
kFjJWgNPgUZNzAME2gsMPA6H2Dfs/xdZ9TCG6Ppe73uvq1gpb0GXB107tNQJme6aPxlcmgIzPGJg
KA0kZhWnt3m7ZWD8hy//I2deHQTObW4gTBShbycKcXDfT4Mjxye1wE8Lsx5e9JV55nHaHPyPvYd/
16CamHcbzDJRQ/UpChkaTAsT604ZaT6a3yl70+QGW/iqAxKO7HKkJfFnI/sKSp3GoViONbEMhUYu
3RvBLbLYJU9VLHDj3krJjvXf/QeET0cDcfnUvX8Yo3jv54ZRhlpPAkW03KMpZFa5Fhftp6PqieBz
B7xMqF1b3yInxk0tI8StzKOK7YQ2iuH2g96UVeyvhVTSASARs/K506/oMsNSIeSeR0U3c4KnDeRV
5BTyw+TACfpFXKHxRVAzwpxFsOlcJSybMAuAupP9kgdPIjefoJ1bA15cjLsVjSfoisGbiBRmKriI
dHvUHYZBuZhtqOOvkkT2MoIS7OCduVRoAsAaZthk4KmhOIDlbFIwvRJMhTMPTheEh4xcTUqSl6a9
byxk1Rp0tHvaE191uKBoZ/OuZQEWQ/pJR9NlR43lLSpQ1i0Az7KLPBYrpkM3Z8CtkctmX4Wcc+kP
EilVrFIxqEy4URuBaXC6BPheavzjDaBT44gJthU2eGt1ODlW+r9F9KSqu1Fjo3oqgmHUhKX/LHDB
8d/i1Ly+xLw5bObhj5HqCjOioW+l7DPxvyuJR/gIUh8ggMrlN6S2ctbrOwOESG6C1njC6OQm5Ly9
32w0U1nfeHsrv3yNk8QsXFrUBnjgIZQp6zf6ULF2DyX+rBBg8QLqYNLy0Bu8Gj7VLlRaR49H3/uy
T9LOtlRbxiuYAbllrwAWd5l20fWPN6diel/i8UoN1qApgrn0flQlXWqN9QnE2T0TnPc+ewpbpOIH
HjvjntQFA1iMzqSNabi2B6Mwap1noydWX0FCQ9TWng/v06M5ebF0F8ZIAVvl95dV8MwKS1Ukj0lS
hqIDL0b0kS9CCA/iFf5djroS5k5F+/11zH0OzV3tKgjcZroxmNhGhH9TGOc5vDfiw97540P+nvi1
JbxJXX/P3MqXma5W7UUHfCZRiq4SATXarMH+LnPLV7qzCl4TNaYFWS6noHsttVlrQRobM1LRiys2
AfAxUQXs3f9Mj8zCJqz6Fw/t+YEbjksgXFODIPeaI9pEi4uKmZLOeFhmlyxEEMmTZbSCbQ09dniQ
NMb5WUhNGqhaSPbXjMErr+4NpdHH3JWI2N5hsuMX/JvxSVkZucRyFuJJH7lQ05BtSFX1nr5yXcwy
Oz78Q2TobkGeg6VlTmI3HQ8Banv5uLwPJSZRbB7ePe0D/uIk1wLxtl34Qwrzxji1C5VrnY8Iuyjp
jvsjBXt5+8SuJ6sk9fVCOZSxcAuJba7oclFtXmAVYTik1W8X48Wk45Gx4NNv6M7zi4X46AdnmGyn
hqHv2hl0B1SEptF6BbcqXJvu5X5m+xr6kGVZL/bLQa6EMywYXz5+csPcFIj6I9GJC46sEqF0DaEI
rv6OGwfD95nlPv8lchGQpeqxyXjOLjbfWchVLT4ZKl096jJn45bV5+l1Inv0O+15be+BjRp37tpZ
XjtiJ0KqAX2p0bjhDnweW6Yn/8mz1gg7IbGyR5xmSkpOKhxe24FSFIg32QrLa6MIEKxoN/w6r7OB
uEBOmnJ7sTRYu+ThzBhcDluh3k/IH3UXzCMlMIoCNQvRnqoa4xworSAOL1DQp140mn6hbkLS/qGd
0OYFz0wldESURt5DY58/eoAUldTFMrMXdlmP60kuvDbLGIZjV7rxeWBd1Qh94J7No1f0KpbJB8h2
Dw2WAY1thJs9a7DUFUm5uoGS7dBPsi+BjMIpbmFi2YiCFhpNHXE1tYNjQdceYUgir6e5vjI1B9yq
A65tIKO18L0Yd8xbf4Z+xaYshThoR/OytqYj7+HO4gARDfwv5KBaBcBvsC9cd9ZiuohF9hr9pLnX
RXU3c9UmfI51ZRL2z/MxYsOebSBJgX2pnViD//tOfLgM+kciaeLV6P7gm31F+lgM/N6mps68wHVF
xmwuTLK6fm+DTD/GIbp12N74WUXfhyv6eeNbcMbYp5vG47xNHG+DXPju+wtiPoSNn8C2FQ4oC2qH
ODwBK9rYD3Otj0gaHiXddiWW/g0PALvgjhOP1qO4fXzQywuS2x90nA8KYumYaIx+xXF6fL5mSvhz
0cp9VY96vVxR5Ks7e/70j9zg5vFBSaoEMjmu7OVT/IZft+vbkv+HqaFvKjB+ufTE84aLwsDP+Wu2
V5kTgAzg1zAIEEOJW5eu7LO/fzDcKxF+BMqLVleTNNF4TabQRXmmP73VWlXV2uYUwGXS23wKxoSG
TUnydNFtbSpUlECh/5Flb6YMiOcbdiwBRiazyPkrC+znvaHoE4QDPZMDKNnHqKm1NfCcfZMHlyIk
g1zChTw6OAKsj6DID0MOvnqHD/cZx1BKJayaNskmVfVjTy/vF+g0uSTXBjJ9UaI/8y1ypal0S33/
ah5qPbcGL7ivzkwznbtodYwJQT64pvZ1oIyYBTtcrc8F+pfLj4PkUqtAglEaSyFzNm/Vyv1c1aO1
tM6V20eO370d1nFj1UtS+W4YHjJ0wJlmLaIRNenn5KMQaQflYFXW+f0yE4GnWjb8HRIyXTW440PG
MSqc/t5AUd/0+HVndx6XChzfU3o3b9k86Nd2kH+RR52Y85/PQV0sb+mZxBQT4T8aRQsT2Gs1jr6F
Enah2xSiIaerk+L/DW2D/1op8k1/OBmvDSwhgm/h9oUmawH7c5XWI8JWNIks2H7m5g52TxqlSC+3
GV+z0UxX1XA9etNhlyq/kXfLB/6HySBbkhlrWhJiphmOSZSzoxm3a1mYYsWMSvHMb9Ld3IrZKHna
Uvn/0hGGcXgXnnoPGpnoBZh5wP8YoufFOq07raNE/7gIe31MIKdrBwu7bOZC3T14j5fDsEWiXSmJ
OlU7GJN9FzzDYxWDw/052Wo8OCzt3D0a0hzxpmRz+cLwO6dtYF9kHPWArMZ+WFO65WyrQr9Xp5yo
qfsh5vjXr3i1hPSAskTSWLWCVzS6X5Jhdep54kuHq8yyMc8NlNK7zeY7v6pNGYqGFnvqilWBMhze
ME16q5ST31ISnpq0hUPkePR1GV3wZZ2AyhoZaaC3/Ne732KAYZK4lZpLn2DtzDlRmFOPiyTiFcBB
IcmLn5KgWPqBMFL4E1pgHzZSkvjSCG1eFzFz6s/YDuVId7lk+Djkd9NxEQJ4LPF8bm0FDWt709w8
Zt5LAXIefy7K/TEEMBR335BBXGhtC2zzquwuKMQYWdZlgDPtLf6IZLzJslf3z9CM1qJm6JI0slTY
HQyRJW0tNamcFFJ89Fgv/GQx1WIEuhhAKskY1jQUeyHS7wdqTzZyutkIE85+4L8lJLBuEfXHkfn+
Cj0CXAAGEDFK+SmKUQyAhpbjcX79hY+iwIVw/s3K96yOf4zMkhobnIqfs5XhrmCryYjoBpyPN95R
vKQXGVltjRQChfRRcyM1ma6vkTTK8Uurh5HOQPWBWIpBNeJYt7Fw3QwpSAnPDT++95fNqxmw5UVz
kuC08vFmTgGCpde3Le7T6/lXmyZWTJBgQ1n+NEFIThk63Km0qPXdmdaUgX89OxcuIMyngJHX14pk
zQaMKZmEZ2oq7VR38wD7jBKmj9JIbT1KCki1ypSfYsSUyZA+Av6sGxVuN7BKZZE8hWqohBfAQkCX
sGXXoAhHRaovQSMiLGqlzdJ2D5gc8/BqxIDezgb5o1Ej3XKVZ9C1L+au4HgJGL95RpCGNKeqrEVQ
SH2RGeZNJBR5MXSrLIPJgcOujnafgPA01f5fyipIPf5SuEqpRc+KUz+JCvylDhnHDIumVqgaSDDB
LEy9xme8x/KjJ52d9ImfMFv9hjzGPCG0qgo6IJd+i8Dayy0A5OcNWiDwX2T5UjQbsFAqgRWnKhXd
JXu2sYAK1cvgZxnrg2xn2mM35HJOFKd2rDSDcEm7FnzQBSKUkgc3Hkdo74GZIGnIsWurAagRU2gW
HtPX7rFqyCgG2wjzG0vqy7jfxYREQeY7OYpk3eN7i5afXGOlt74k4fCXuwHpHHtzojWY8davXHbe
YH/pM2wfx0cylfrX8/X8DoleR2GiH0jVg1NCorat0y851rv4w1Rhdp/G3jCn5i7s8xGm2e9GqY8b
aywJf/9FgJ/s8j0A59x85BRQrwBU0Z7O2x4ESM3podMEl+tlbcgTIN+MM8RLSEw6nPDAhvdB+LEZ
n7PLs2IqaWOzvmemopbE1qYc7DwkxV8p0oy1vhqu0mxUaGxmsHmM9QNoSHwTIrR1zhr9XB9aacnG
p9mPCebLttMLB4dLkYYZqAkZuyCy72WbcVaT3VqRUPEW8fXI49wGj4oqv6lKFoWJA8rxrXQK+096
wnIAXxWdPov59AZrLsI8FWBgsL2yTP7SBAviUsjSJfMs2xyMCEganlYE8zf3mgAtANDaJuFW0HlL
n8y9oy7Y6C2U3ZuJd/R/lFyCxaM7vhj2bGrRpVhCDfiX8s/bkSYFGk1k26eUn4J5x4M4pHFhIyp4
wghcGJEGb/oNbUQU+5+cebzELKF6g8Sk7BMgdxW05l9QnYm9CZba4wiWFo7AHGeiUbsaAsUbPvK+
UzwR3Y0EXBXMhvnIjYbXQPmY1cOzm7Fpb9c/oSX6bjHXLjAIaNgLybhNlNzCAo8ALgkLgMZm21cc
fUVfm7HfvSUbAnb4BMb6Lgb9Kis9Njgy1TJ4mdlYzU5zFU9b2KiFbyrGZw5DtlZjFVjAESpeTtgO
SVdlhdcXLYN2TCSIt1Sb8HVsb46GzRQueKb3mrjAZY9PZIk/t46MLZSEBysCnlhAVC5sxhY98KiK
ofuU8CspwyrDUaHK48U6WLk2qEES7WBD5Yyq3JH95thHQXgHVbXujsaM2eLnY1lRssgVGH8Z0jrW
NCxMU4qQs5XNqY8eRVSyVAXSlWU+bGSBKnru78vy4iXQgDe2U2s5fS4WMG0C4cq0pRsgGC3WQlto
ZkWZ1SoJbR8EdLAxCOHsz9dvhiS2+pOaGp+EfbyJs8AcMCq0d331S5a+nZH8uYf2g1rn46b6DKQ4
Ajyulr/lwwCizumfPsnLgA1HiKAfdiyRemMAJzBzHR5yxcZJ5MYDdI5TynQSeowdsxppgeKh9hFr
qH/tNRGWqi/oKzOJFVikGDZuMQuUvLibTg5zAksH06eOBXziLcMPBGlZf4oHoXUZRXni8rFCnEW4
jeozrzgtFNb477rfxAM9jJ/pbH+c/l4Q45uAl9sNByDMOEJOOTNLNyc2hWwXGYMAotJgr+01E0+m
1VcbaCc0gfNcorURGAah6ZlK7w7/8y0VTZjxbsx6alamF4r84C55Ut4A5uO0bi1PKPN+ViWyfkB6
gBnGbbEIgQuXHJJNSJAwq0SfWCwYK/XHHdte74URRsON6f+faAGxzhT+1Gz4K9QpeGrsuZGvMbMT
0qo1yDQUIfYBaYd3UF8qKh1EL7WwC6+4pf9TrXOF8Edd1IG4fAopFG6iLibIkh1nIxg8Soa0pvxY
vf21ptYJLfXGKWtj7pis6DtcpRSWdVHV2srvgeNzoKt/fe3gSdFlVB9CB+SCYWUUNrNuTw3qBBku
33w1ufXccp+8ROscf4yKfJNrOsrHlm1gKMN66LG8RZj5kOvEijEiZ4+9IBGQjXDM3PNwxA0G49Vz
/+TEmXwB+n9ivGcaAZR4QeZX75XowROWxUQCIENtWJ/wk4TfPvNAtQvP/yTDgRUe/5WyfFQQxVf+
zabL3o8+e7I3oq2lPD2xvQCrTaB/GHhOOKXZQfwWPFw3WDk+13WZk0MApAzLm46vDCEttd8jeUma
Ys7m6sPhYDPVV0gOwxJbRa9RmGZOZgim3/YY6HDzVOq96FQ3DyBd0WTpHAtNs31rwcAK45ZewAvF
G9Ghd/RqzwoWmiHuKf/EAECdEP5/zZtwcI+HeIzPHze0jYO0hNLPn2EPcI3wv8RaKdSiDrmYsjgm
aMli1LUudMTwdaDWcCMF6jHz4acl+ViGE72oU62vfErqajb9y+GMLLCPq4i5zaCE1psI36758YD/
4+drODtUWn1mVvXjb+bR20FO11Dwd8CwtU46uYT4a4LjXVz1z7EIUFeY13kDOAJKNl8alA++O9SY
iGE2MsZZaJ78MfItalJSKjnyeeGIiKPeKoFfO3b8lj1xyp7rXrQHBZQXlBDBOPWUznaCDdd7QoAr
HvtJXc+gpaYIOpi8+qQ3gpQtCU6cebPKehFC9udUpGvrzRAz2yrQPXpQQdfEH3vJ+KwT7oBq7Yfc
wZ2rwy2LH5gn8v6KZNcdW2GHh/Rp90Q15HDW70QCK+MhhdSVs4is34t2Cmf6ZQMDiRi8fxk5o6+/
SAPNTEpm20QauDGdgXXMugUUydPOlrj7Dug9/dZTsMEcF1APgxSLdFnblDzMzAZ5F50RDDlOetex
uxcrqn/EHqlhToQbdMj/CPBnlg7gRFRw6O03+3CbSwkNvkWFuj2bJSk13VXyrmv+8ONYQvce6EMQ
nDtQoQzZVsFPxtWhWZyLLcxdrGxGou62IYB62QXiMSjJmLqSRj7Jc7moO/6yrTyJymITEF4K2tdz
qjmRCKj3j4KA2XFd9En89QyioxphWSM9pMAiY4CIUl53kXxP+Luit00QvDx8lsZ1TWufd6SkwkCr
bV16VI8DuHHILzrjiCXZdCdt3vCuA+HtMSZ5Rz+ptAHZkhpNpDzVGLi3UPAolphkJBTMi9yOX4RZ
mQDLxBo+Rr3s6gxpehWidnQ8R54iTuquYRvL+VON4EVgOlI9crh+Jx+AUEfia/EPo/qHzd6DtO6e
HkA9rjY0pGi7C0GP2UFAxi8V033NIU14KMr7buyAKdkvzBVndzjIoSkKg+B2nPskZF9VwmYzUkO2
vhY5f5/a2qBJOWlLStYu8mhd+K3NSgXBRYK2fXvsaxeAnuL6VepreP5nRWd+ytnKH9hP0Yu27Som
VPy8x8Dwqhl2RSqGtul7EF7RNG/wyJ6xR/X+ipHvtSSbdQJoVNZRPZViPoFuWRZWdFyWZbhh0ZhG
oBp8z2IcNfjYEY6CNQLv5XSbhezHS7ZcRePyk06PfNaaru4RwymeibqXYMGeD8PoQ7/ZPc3YuWiJ
ZH+er7C7UMw6IIuf+fEkVRjiMnOGTfgtfuRmu0j3T1u4zZoRY3HPtzvctXemybJt2ot6AF9S+/S8
LBt+oSYvHlQqR4l1hOnrLCIS0yH+QWK9mzb14cdM427uvocFfnpG1AZjR/lvzudq5tq33HFK3anN
ZWaIDwXl6ZOSYSi+7W7TVBwJfJiYs5msAqqGLC095f9oaWbvsa5eJjunb9iJ33gDABZTSm38V5/8
vJVzOEB3dwux0312LcTIg+WmBha3ETX/YvzYlgts6SsOF3T+1BLtq3Hedk4sR6240p4geIRNd5Oc
t7JqpBbuRusEn12GXGyvdrhGV7/OBpllQavVdOOD5xq3v6kNtNXdZUrgKNPvLfYF5D3ixKrsQo+t
zZ74bk0VjD61q3WBc8HXiYyHOWOwxn5JEE7X6d4Sh0oNlmKA0rv57PBpVXQ7ZB2/LdEcK/0eLNu6
di7v6FEApL6CoFP/4lHSVlY1PagePgc9R6Je7wzZzt6a+QBTrkQWan6gt9WsSJXsE4RsrKmmkY4B
CzA9Tu1rTJRdh/xEPWjtEmqCzyCSwtMY62YAHPB/Zv+OmcR1AzhXElIljDmqv/SYw7kY0kwLeTH7
8sMigCrlNDhiMIyqLtXZk+cIlTb5s0oZMFSuhLAWpvFWk4Ldn3dsVRdBmkCYbpd8/OgJP5pwgprB
GNkRdtCLaa+vjEu1ihkm0wbn6oX61wQBmbHEEMU9fbnQIqpqFTlpkOkbUa5D+ntZ1OGnsGwIlkFp
tYmpDek3pj3n4Bzv/W9TpFT3ILByI0AhgY4js0MWrH7ICPiJ8ZQ+ZChLjSgfJmWwuDNE+TIv0j0p
YldDCAdIiMHSHfEq5NAc17+7I/7AY3AXNHvRnh44ImprsAhpDqUyGnjkqkniezS8+ecUkYL359rt
Va2dXBTF1CyR6Y+8qk0dU/TYdFli4omYbLJMEJ2enHEfTDq8FJkH6UHsLC9P/QVQFynnsqKP2NxB
iwWDHfNFgPK+KK7jBnesEiC/cR6n7416EklMSIShzB76EITRvmuTfj9q6JY0OUp7zQ+tikRnyZkd
Mqs+hPLDqR7GuMms6Lx1hywFD2fQcYkeW19xXxOWaUCdjudaRTTd9ZgTb1bLbt2PAJFMBFnv3Fqg
bwehiQ2GUZTRzZ2xChCN1W6UO61wtey6SdvJHYgqgGriDb0lLhHvT5OR+14y6eJk8jpOEmQYCBkK
SEhFe28ko+zxjfqgAi8NKwi0BYxQhVVo+13dLtt5IuI09NRiy6B+Vmwyq/NRVDeQVNDuomR2v11/
ShbSCAAgWEnTfhxyI3gop3eCiAMUy1fsLePMkO1NAeaxrSv4XmiR+qGxN41YeupAjty53SETjCO4
ZNaacg0YIQ+eImcOnSUhlXgodn4Ubvdt2cDOhuRkUOZmHnSo0b9Lg+Xew49RczKnTi4+3/cgGabi
622HpjPjwbmndNkyKJNb0luLBwMl4moT0e+3NTpzD5JFhgBKFijhWyzG5BUtzonIFPuU9uXGJMp7
QbdTuaRvERj6MOpFcYbAMTIWREIeVJlvg/jbx32hgWD6c5J1WDNEyENzaTYOZ381K1roOjqJNmJu
AeMV0u4KtaRHSDnu9tIDxSxnGTVDIRfF9jar0nqW6zV1PRTIlYOF4fZLiSY+P54GFCHMfY7Uj3li
eowVUoF6pdQsZuXnayfCTfjxGS1axn21AeyqZhtFPMykG97GWTSExtUqyaFicwMThcFeya+yIhVf
w7WyR/ur+b1oV4jpx8q/qJpqI0Jtd3ew2FVi+pdloCRCkR/hr4vPDZmk4SvHLhaYukId10IyU84A
mE0/WJdhS/HeMNb/1F2jL/X/UVsmoqqmcVP83cwwrQ/4XHhYCw4aVbM10M/KPjduQKBRz4QYp9WW
hU4rFIxAiGFvdx2JLb33BUU4p8RNzKcAYF6Rjz2wv/sTCQpq/jy/p79KzMwjAWU7UVFOBNg9qnlu
omEZZCcwiVck+hMjLaCMbo394divnyyvNnytTsm6+fIuskdoLBkp0p3DmT8uoPEcn2NP8CP31xsI
k1S7UnJNj7vMbTFpuvvJJePSIR2Qo3cXA4NjEp3F2g4t6Es+AanfttOZPA8VCuXokLiuTQv/c+BB
FlkZ+7ftnEcTElg0FUQslX37q3sCST5IWnEf6Cfq03kUB2VRbpn62thCSgZoWne6ePiKiuc55ZCo
OtWbahN8NC1kCZoIB8KeldqEBy1lpyrCw/qbuXXgvIjHwxO29rLGtQtD6dNT/5f2i47RR/41qsRT
hGMZgBJ7C66pTKhqbuKS5/3noTYZTAEk04YkqObNfcPogZkM6L55zYdouIIhV9T29MmMGUecqwsi
dFb+Cm2rjuJLBdwg2tCQ2/5a24YUfDEbSi56Dhm1j3i73tvBSNrcMw0bSQINWC4w4HUgjZ51fR9Z
T317dtOQxXK5RRbxRenJizoH8yzNEYbR3VJSY+UIgvczK6L01r+HgHFIr57k620qwyP3SSj82x2z
X6Qd66S7OLC53VwVMb6S2S2VQ+Ui2TGY+HaWr+enAOg0VeZ4p4kfHywxpXftMT7XiToiNFs/u44U
U6RKXjHGHemfzQrJAQxW//u0lnxEetxheH7MZV0hUDXRgP0N5AAFoabaTPQ76ustyrQALjuqTqXs
9TY3OlizBjQT60q4KlKvyPXT59Z9egIBqZHzZpiDc1GZ2JruKCBAaGvWvnHXlpAB08CFtoYqYtyG
qqJZ4aSwYKC/0/ARk2YGesQs23dS9PhqZNVqP7XiIhLcBZ43zIN9nW8XQD8Hd+HxoRp95eFNums4
9jC5ElkbVjHuAUcZt88yDXZFyfjI6G04c+q/arrE7wrtlDkfYUo++Zy7lRaDF/x7KWsMGdQSqzdx
fJI8z+W+5F9UZoo0KCpaSyADmSOvOx8rlZ17t0vACMLwCRHmk7lvZNl/9I45d6WE89vsd/4oozHl
g3zyTl5NIA2OzANn+Cb+gnL16Rq2H9IOs9z8f3rQA5ksimb+iOjwVdcTSpGSCL9xIsHQflwjjBa8
4nJRUA7jyI8sZLZSRg4niEvo8NzZtOQmbKrYGF3qQQplBfVvSOQ0FXvjRtVTAj/kYHbKDGXBxwpT
70e27PZHtVnqw0kqhKQJqHQA82rs7FboRSZHPWFq3OMizZ2DtVMVi6z2TC9ehbl+jVei41Ov385k
zqWnyyZretpJSUAgWwpSIIUj3elMWwspNdbXGihVQ/g4Fdly5JmxvzQDknWw07hmKOVEH7Oj+hKM
l5iZfKL7vOv7qs0WxRuBNhkDHgECBgaCRLxnbHC51Gx0S47crZ0/wClPuMlmhieRtuSkAg55UrmI
82Y4HxgOQfYmbSwwx+SwYlx+QV6NLx++NWDFAmnjD8JUI9KqUhlGukSdkJM9/2kMxs0ql++x+UBT
RfD9FSxmq4byJMsMzuq91R9S0gLqwurR6VVEwaUPgGR6oO+rUCVQ0dy2mgkdgi48FL91fP24AMb2
nfkf/v/o7838wZz9AKUwOPq5c1ud6wdw0qshjC8IObF/h5NOWQl5PwST4GJlk8HAs1DBeUJITAqp
nMVI85FTP3uGBfZCzhM+MPRYgrysmgIyw74K8cQ77vu7euIHF4lW4vL299/beYJkSzYUypydIVUA
tDDbb4RTimYf+w6k69JV/YVVa+w8JLvgMWlgaPjqeIl74Fzx2qv6o3KEkhtsey41pvMaV2uwCkpo
yCxwuuG0gKKyxOc5YpgOqYQ0/xksVAkx4/mGIsrsX9rpuBE0IcLGi67+pyXGdzYKDZrNzk0OcZ9D
y/xSn5gAM/Y/1aw26DRXCSYrvTcNW7swwfjrbxN6VilM5VGi6jwaL3L290jS27ytRD7F9fVzoF7A
3nOLNeUej7hGE5gppLQ31HTbrXJ0WawybA4CCAZfCM0tF5giLfifzUtMbMjyIS8xdV5B8IL8UM9W
Ofxm6zsFNjuiTFizn5q6XRJ5O3ZvNotAuPwKnAjtxGs0a2BJz3UJCOzHS42pV9thIRR4JAZy7YWr
12YaXNg97iOXa+Ug4TnRK/ALbqEUDgbfH4iw2ef0OujKEbHGXgfZtMVwIAnciS0MxNhWOu1co3Gz
JDL0iHXy7n+Pf+DVeBZtZZ1dt1gLEOVb+zZ7HnBGL6e5k2N7urJLDrjg5gi3yVNFCipMDQ3wFLuA
q1EV63dtqgFxQhPCc1MCk/L32K4XKHsh01OzAPOr0Q9HUiOUkUKSY71++dzyID8dvbzgMoeVl5t6
Kr4a28nOl5h7lwN1ppFn0fX1B65yM2wXGFryi800Q0kOPiwB8S2vzLqNQ9L8HKk8chn17DdqOA05
WS7N6MYfoTEuxj+0CCrQOj7m60rTozQgPvjhFGOwZCKBO2+3rrLbVOdZuuG9n1+PyrvWDIz9WMUA
jtVHSOepxvxKtlAwM4UiQGpErrxexzutnGfUKfxep+rwrvF5kZblzfNuWqNfuaavFdDdT30H9P1l
F/j8wIP2KeuypjA6Pjo2/NYPk91DV/1q1lYMXomzJ60yhmwDRZl183WwGpIXoivOHmcyeDSeWuED
rkj8kCsgYv/D+JI0GGwENL7DyLA3RkV4HvFOwrb1pX84fqiyRqC5+iPRQ3Xpq9Pm9FncVU+YwU8Y
Hav4DyG1+Z1NifvJngujgIIu4tQFl1bnmgzKItAK1R71YhzFzyQh8rlXSkyBCWCLLseCFcJ6cVcQ
pWLWRpfaZOD+mi/Ys7aWOcZU9+XMR8xBG4q2KSO/EfMcKqXW9jUFJXraEcg8oa3Nl7tMmWae5IpJ
w8j2t+aF9M0Ell9pHG4JQN8TVwRL8jSusjD4HVCbQR6shXNmS1VFy6D+AU9kV7tC3xbErLzBvWeg
cbM7DKauosq5Q2vrMx80UrPz2KLULx35lbXgzFeHLUypXNC5nuAO4CS05EuPcCOJnNcD9AsL09Jq
Ncw441W5ZnlzLIB8oXkAH327AKXQ2LeTmKPNVd7M8jv85Cd2mJWyuOt8w/AfPO9D1H9NTUJfX5Xa
oQ0G9MPsWUdcw4SKb7XRAe9Sw922l13p/dDew6j9X19mlmNkP5kTllbU5X1J/4lMzSYPx/D32ac7
EwmdoZqiH6FMnkTWcLxfG/rrmfEGOQl12XhPBxQtNdftSxCgTDHoPtxClCc63tnG/LnDOaLqQGZz
ipUTeuN6f0fzEZf9RI4KwJ3WEcONTl1iv2nVtuqKWUWVHUILJOIiV9Cc0YNIypZLBGlx1doHaTmD
InTpoRdd6NUegAddODbNTKelY84i6WuziRe3iwhfSXKLp5GGVbDsyDxm1EsAXBTEExKcBMeQ5J+7
CxmnDNyhVNASXOOlB0IKnxxQ2zG+7fAzBpX1v4Tb4KTyjYAB1CoiIKRsZO9N1pGdifmnNqNnG9tp
hPRAoBbwXoJZ7KwDZYAGoD+/eV+qZ2Uz5x/4eDKxr2mjFbcSSbEjAS9ZIbiRWN359pVuEe4pRU5L
jznGuuEPZujpxNqta6g0/y37Tl/ACMVg7WPKAxkAcce9P/iR1TMk8DM9feZg/4eM6Ieju/P+FObO
KhAB9P26fIrW94q2d/Rywj2qMJdBGkhu4MwWivW29WcN8IVBEchuQIJMlKb+gUR6jlkZ6vd/vFcu
AKbozWNVg+GhVAVMfBnx8HTO029G+QBCcM45wG5r0EDrhZm2KKpjSEok3uQ9nVr2sUQRMw+wkZGG
kkTwo1KXnHsyMSCK7zDhxA4YE6cUuOtoBOquh+V+RbbSnewXbbZliKgfwxLdO3MckPtyRHyTU0fN
uEvVzq8PDFiH5zhLl6lo3p74YzSuMLiTqhXVqP6BjS97dACAtqA+0crZgtMjfiMwjxUatv7uwfV7
scrXzSwDeMx6E0C3pY1m2vZmi349vEzMBqRtiVvoCKy01fcEskskQeVHZNOEdFIW+tHy1siysdVW
hKE1j116kpLoKMCucqH7aUe0Sra/PPrZM3yqpd2LcyjVOeg9Pd85A18XtIcZWPvQXmxQFLocOwDf
ImM9Ec6AiW/j3fNYRzU3Ju5CMubKVDnxPFa8z7clMZclEqaRgKAAnjnFdceGdX3g0v0pDDjDqGRD
9cc5aNYmx8oxLsP7Oe8fc+/jL7g0gNHFL6nlEv8EagcNi22lFPzt5wZmcozWwbVudQS1CHypFTaq
0zKZbHq7qlIXWF07NbLKEOoMgaLq13y4S0aEWL9bJ5yibo3tRjLUAMtJr76M7wsSpXAN3JidfvZw
TBKPCSYB65mKY2Sm67eCb3c4tjG9i1PRRCzzpK9G9vrzpwMvGXDzHEpuJ2YfECFYOBv/DHcJ/V7o
N4zUhXmpa77pX7ao0nnnYUUbm7YLvrt3ZtWKjSVrB5ikziEUU/oHWgyypoEQqC1MXc/e8c7rYD5z
F/xXD6bQgBpbThjodqZotf+7pH7xb2qT9pft/8ZwWarFMfuewPLlONBKqKKbrTEduJqoBPe8tfm3
s6FW6+d49gQ7lZVHQlNbFQGvdko/WrNTxMeC+t7O1D1v34L+S4a6QuViOO+kMpkHuWXDSurvggc5
AWxP/nQJ1gCkE5B4GGI83aJtF/UvhtM1i0uxGzutaPuRrheRp04MbgdHXf5bBsVFWL0BsdJU1RT4
1xFmxqiF5PkmXTmbPK2GU23T7TIaukQc0kWd+9nXETH0LWTzQv5MHN9fQhK2MYQF7n/WsaRDhHdj
jLRHm9dpOYLyEPsAn5vC0+ndNbIGjnS3G6vRZMTsmCLTeCC1R62zpJkHvyowD0LEtK1yC8gwc96j
/8XJtpwLuUNLZK/gZAAezQPtJG5o6czhMWm2wOZBP0pbmpYi7aSouwW8HTzPJvz98p8QlHMQVVPm
a9Sml0d8iOJDBKTHEY4U751gIlArnrtJgkQLOAKew4qLLTgTS6gbiUIlUziH4/W0eN4esseOqKRT
c+oB5vA36jl9nklKy9/9TyF+g9bKVUZd/6lD80rnV7T9K77jzsmhsTndwtI0y3JdVz/vz/glh05r
GEzaJuciJ7zplk7KWOXB6exzUKkctcUQibooZsMTb//F2grD/YodqPKjgpaI9f44TSiR8nUp/F+T
wCoxHeO5qHKUEh7aFEvZxhLHh20Rta2doAIgzPmWoVCVG03eZ2k+eoqW43KsSp0WLTf5nNqq8S74
Bh8W/qJoMV+VOrcttX10reGqWEaOg+TWvGlcrdASyu8nX4pGKffiOFm8HH2iKkAdJ0VC+15ICa2p
3I4ogNAxi06kRD62Bw0ldU2lgMX3oO880f6xqFwdqaObcw9djHKEnBHa3dGaT540Ibk7t48MXI39
mRvoVp5HdSJGhUa3tS8y49jFCy0Hbx6Rnsb2Ty6+x7VWxHGKN2lWymNN/m04HVXlOCKzh7BjqmY/
qEcKS6Irsax9AgAg2z1fDLn+R9tjVhnCQMNLm5qIN/opDWO5i8/7QkBxQbkRTeqrF0UEUS7hwGg/
69z1/ep1G2OR6w7fn/Rm1pr4GFkvTEj7smk7JmYeYU+XFoqr0Hbgo0GGdBkQ1AkSqw3ek6CpiE4N
Y73Zl2ymtspqdO3b4axHDX8PHyERzzFR1LbUwNyIGb0t8Sjbt/soPJB1gKgJfdpBUsVq6qAtrWKx
giMUJoyWbarTRrdT6xeSYqH5WmGKLaWyqgKrOD1F7D0PKrut2kgx+JQXBbyOs3ILY959Ks7Udak0
ZA1dqkMkTM/ndmENuhqaLcjBj0EJPfSFb7TADDBbjK/vVjnNrmOs9PtwQ1yBwH6J9qa+DFPzlleP
Z3hnb2KyVbjRHlAiWuELIy+tLniUFNHa0N6b3ZSbhKTz4SJGKLWyDLrPIIKIJSzhXYMVXZGcr5BQ
I6qGpJ/X+DGBANfBlWYf7ggQGOcT6RnUoR3zuJJaIwaMbCruKjpbEm/tkH4JlGGPxdwHXJQc612C
GMHrFPmMKk9ch3n1mGtKO5SL234ZPazSdAnfXob2E8D3sl/mwqo78w4cQVP4HZH8k5WqRWemdv/B
nDcYge3EJcA2h/Za6/FMfa8v+7bIgFOLE6xy1J+f28TnMmT77OyirMwi0ey822lAJWdHA4aPcX9k
U68q2O+uhUcHSawdo9hC1+7PMojzABROeRIrNpSE8/uR0/F+mmEATWyfvj8+nMW2ILIXcIumgh4O
/RGWUBZspnCmligzseQhcdFJrBBY3Zko4V+55S3augnKkQD6MQzWDdDPE2oOQXxZwc+IfDs6Mi9r
KWXipU8a0th6XOzD2xEsHlZVJjMWHN2aB1x2aZ18GqaJkKe+qhbRcCgcHrF0Tlqb4n2ElXMzMyvy
H0bUQ3Fa/dAPRHL+sTd15io0KkCYp2wiHYSmaxWhIE2Ho007KzjASSZvYad/Qq6RXfx4GBpURm3r
4iQ5SJtjLSKrOt4MNfeP7r+ysVPO8mXVaIYPKg68y/FwK0nkgc534t19kITrmLVm/gkE9p6RsNBN
b0A7Sc9g9xykaLcIvMU2XLnR6FQglaBYApKP/MOpX2h5oC0x5hSmQyj2V0XLWcWFavWQrq2OiZyA
spAnr1nSxIRkztaVJ8iRtE6UIAOOXjQFC+E1L6zommiVTpbugXe8gw+T2thZPXNv6b5Kax5AKiF7
xSLoGr9l5GcYTI9beNnt89P5gOSbOJd6WagH3KaFT85hDGnEEG7uDYZwEEQuIgD245D9pPxu6qSB
sfTDc7FwAR30TUHFb6gxaYqR9eDQKNpUCl8ayQgQAt+xwSgq7JeMQomWXcO6iLUCcG6Wp8YrJR6t
Xo+ijRMuuNS+A8IA1WBaEaGvUC6SPvAl20jGT1hzHZh7OLeJMXuSTzt+8+r50Wod5eOfei3DTXQG
zExz5eVSAH6BD9xczAdvHQ75AKqKG+5xyX3mhoZ8s/YCSv3+YmNV6YRSfgugdCetjg2IVFZNLlje
nxA+5OPgRch3+dcyTp03VCTVg5C3wc7kaEbX//x4fkMU5bR07gskSrL3jEHEB9sqKXyO5tJu3xwm
R8fvVatrkTzcP4B26nwEDzuJVu6xsmrDT5z3RXI7DdZUA1vQtOiME7QnsmNzOVtU/lSEJlVSeOO2
f0F4Zurv4JWufIsaDem0lH4qE1brG9PS6U59Azy2jmlfi+yo0QCtiulmAeCvfhhM7BEaODLEf5nA
/maUNhQ+du10kg8Vz76a7QvaiveE4CDKHLrpAsD59T8DPqBuAiZskElX5PZZSMlA/xgncbq4UpFK
jRBmHGNDHsLtEynxWBDq43gHE+QkfUxJUGdliGUJUhkl45gB2SUkcmLOnTY0ay8SaCNxBmnVBjfK
Xvd806V5a0gQPTWHn+o8T6dAqgk6yeSk9Jf6rby/aMFbHknGdvH0/4KYa7k+WhPIcU0nJRn6RUcP
AX0BNY11HCC8aHAzimpv63gljp0EKYHHcPoJbJ/MoJ+34LhWHMwFG0OOMC1iSHUAL5cuqbzw3DxS
l39xuM4l5S9q/2zP6GflsxEzYlJy2VFb2bWe6d4DyOKC9hRNf53hi6VjEE1LA3q05E+EQADrG6l5
eWfdR7VHe9M5zBlE1QbUw51Dl7H51oH/QuBQCurL0FHU54HsC+hiXVDNZqEs95IWddwsq5OmpFKN
v5rIbLe46dboPhrQXheCj0d/nDgrO5kmI4m909il9ro5qFO8Sxxul/NjOmTzVO0T72XXFLPhrYNb
yczj81hdVTVjvUpMsT4dXs7jUVmUDBvaFglh5QW2wxtwNQfr7F+4rLfVymNo5PgzoIFX2kgif1Zw
/PXw0RclviyBwLYijxx+86tSMd1ohxopBClGvO4jgK0wla2u0S+aFAcu/w3CDMEKuQZxSPCwSaty
NJKfxlM//TxOsnv5N6vBlIS0z94jqcvI5jBNJIaca7Eb+ICAAfcG5DhdIxsY2uRliCNE9Re6gnjV
5pxHgL6yQ2oeZ7zbGRgd738lMnrMJuEbDGZIoyHCrwLS4zXNYwUH8oeqQsykerGAJuA9Pi8rKVll
qsBIljJg6EztvA6UA/FRWfRZqt5Ad2KroS0UjcQTxZet1kSl+SFhR8vVWp0HAigZ8MojzXi+t0SF
iuLF+I1vK1T04afIzHfilVlGjlTbR1H4ywC1yS/F4D41ReG54SuVU2IdnltmLinUtO5HQ0QT0OaV
bepXShOs+GulyeQDKU9zB/Q0sJgB3QmtWIviSoq12O2nJITS3HMF6XWZda3uMX3YVG+rmF5jGKXZ
ZXptzUDvjNdynHub5NmZfFjMGPiXRqShD26xfyv3+Fq0wcm9SEFqZBLcPa+Gvo2RtuO0eh0FBLNH
z0RIcnHrfWZAPUaoPe0hVXpMkzVCB5785Fzn0olP88eVQMYpY+r2Q/rL+lDRmojcqce3Sr1WL059
DyQvGuhJZAbjcZdRkU+B4jqAORQ5R2pIWJs6ICiq9Fb4EFVGhyAdu/5J3EWwgELlTgQ5MjwZxpyc
pbMfjAVk2v4DJVSeUrWtM4rT43FIpGjI836ZOYrBUjUT+tqyanG9M0mO8D8YUPOSt8bAJ9dpasKP
gWPQEClAOiYodeYwRrFB7NXVZGfq/m6en2MKPXSG0ZazLymlwJV7pO5avM69F6QxFifSUYNKvZnt
krs3TuzBI1N29MIafOfKybcKrprgjbokn32e7SOLqG2VedogqkWQKYzf6KI7LiUmVpZv/PkhH7qO
C9VrZE5znOhDkvY0T7Gv+cahXqMqKa/gxnAD8wgxYTSb1nhrkn8WzxUboqWoaVNzkFvYEAvsOZAk
eWd457HrfqHNvxJ1iUV1h8aoX1zIdCiwmSVgN0mIP8BdEHuChnPz7MklSsm9VQNadR5xVpjc3v4B
X3lhM0r2LmOJW8G4TuxlsjChsdRf5j+wI3qucOxuLRHuONkn/Z0psVFVQq1w5Jl7lrfXvVjs52Zd
rbsiWcBy7ywGDOtEozAwEYTg671O/dscmlvHe1cziHTp4IS4/WJgg2husDlxqFQhWl10NMDr96AE
on0G4oE3Kk9boyrOSm0wxaQ4CcRbu4nlnxKTmIjZvbwVtn4qHdDuBwMMAe8IyDVODRvFJCHiSCmt
HaCanUn2CoDIrrqsg5uTOygTWhATJLjXQvSvgAvSK/jlIGjfdr//jAbDg4BwPH640695MqqiMS8t
FPi0uSw0k3Bc+Kuc8YDCFMcnHevP0bifBCwDxHwzPLcQEa0fsx2sjZNIcHKfbSTDsGNMR4cM2Zx8
q6RLQv2TvraZi45GrosXOC1J47YL4j4mgyF2GsPYS49zseWpAS8/KCJooQ76sZT48lmiBD+X8G0x
Wt7dPGltK/Iem6c0u053gauYpFdj+BmIz4NE9fVHg5Thdz7MhMrkNBHbRDPKQnZjeyqxEg1sFkQM
/aBKtxPCgPPOFnlKURtyslF/eFp/GWft1I1zQRvCtpvmWqoRL6h7QM19/vzr6SuJwdwyDBYNKMQW
TDaW1lrhnHG7M8F6TqlXKuR7E75t8uwZ4sVif15/20SP/pGNE7EVqkA3bmdA5ao4kkS5FLUuTbHA
baTl3dO4F8tgq0z8xlimumK/cEO2+j1+ZnqpJYbygpNR1OrGq/utrjV7YdP6hvjgFG6oWi9aeQHb
FL8uo8thTIV32mAESobddhYAOFz5KCgGscw9r6nAw835+msR1uTw/dap14qGvSIgydREzqPQLI6T
TAPIFltwUf6dSaFL9tQj7ZCHiYssNxz7eeWaS3ZJ13nfjFLzdP8ajvEcH4M1H0p1jcNGta7c8NqM
gNl0Mh5IHsN86/Ee7pMYPu9+8T3CiVKYnfuTfWBeFlzfgtx4Er4MIRs+FebTBZnSRaPUyuvdvpTg
8CjfCltQutDOCziFOXME9FxBbLLp+1gWpY8WDcZ0aZZL48WeOMTTBpW6BUpe5ZTNijkAVxdskAAu
mICFrwGeW9cWYOo+5vDoJzyZ2BQAu1oNkAtSD+d9Vf6hKTr2FGA5M5RQTg/dhpLZJ0U8AvR5K2gm
N7NuJYUyD7NUt3nYZ5EsWrHNIol3xXRCm1jwuEilTV6kASnjHxy+ldcwTLqI9AybZRoIEoXoAUS/
36ORc92qlPx5zM5KopIu3JNqhLlRhF88RWP3SGmRrHieSxWwYQLxo4OUiPdys3NNDSTvD9IAwJWW
W7Zfcanup9k1Qq8smfAWJqWjxn6orLKYQSVOTWo+83fFWf3hn6SBVj82qzINeV/S4Tkl8a7dkYlP
BCoREHfetZqIOuI75lpQtjFB6Tcs9yEgCa8+x83RqdIjZn4PCXFwK/yqm05k8GLxQp0itvBBE7Lh
WnkbDbtcCcEn5IGTnVNznBhxTrH6v0VqxrrPhOileoy2rCAuvHemDRk01K/kAtmuxe1Bny+ifNH7
b5zPXEzeuxtUFPkY3hocFlHNRxpCfm2J5XOnRTdW9RkfTGUqgW6Odzt9y6VER4AGkTnP3jmqQ9jo
V+0q7p4t2ucm3GIAI4vzIyYipVC1mOZXcbBMvZfSCXI3fTkweVOsG3s8FU8FZhHeV4sOj5DLzEiL
iuA71McnbRsK28RTLlxitfmnDhjO3LbIZhevR7KFTiEhunTVAKfJPKvD5aoAOV60cRbb2n2M94+R
0d98L2daQ0x0U+N07kUJpoHZvGVXZ73fE4REvdtGBp3qPfzCmMfGbgFga8cRPw0y5qhdDa59goIz
8rA2QqdNoXeM6C3ne0eVQDCNoZiU6H9XCPGB0FnUkFCJY/ziVWRFUx3jdsHVaAeJNE/Ji2BiyigX
HxMnKstws7JxignPT6f96p33vnNpH8o/aIAiwE215bjE/fr4RDzQ3/EDoapUZq+tbm/1OAu8YzkK
2z5W6/U7GfO39jemJWaNJMrNWXYyx370H7t+y2G8goxTENMxrxcpSpmKdYPPHiSU1kd9CvStwPri
wJ6hcjqvucKE88XedoU9fgW25Vnrct4TTz5DmIjqBFFATf6vJAx+V3eKzIYpP0gMUYkRPMY/oX5m
qe0kvuhjAIDEwZoZs/bhspT1subPvpN6Aj4FT81fb9DHGsZCyyyVR+RTPtwjVAnqlvWkwpe/LorH
EN/jKt3PE+1Pg2ws43sVjOoy4GNXjIqnZTHq1D2/REPMaYZsCg1pcTzoSZIsQXx9P2Wj8iCaygPI
jv/9HWx+zBVwUSxvkkYsG/FXa20LRylUMTt0s4y3RVRPcDnZ4JmjaLq/ruoA+fktGKbUaU6ewr1Z
hYduUW0iy39F6FvAm+epGzVAc8KgbqqSrffDILhfy/CYy/JSFCXxSSp+L751HeJBVCRCifo7sNc5
ou2havBip25z/T0AeIJiVkDUYCdlzFiBOW6Pck3Kvzl1uIAs7vqT3GIbKW7emymgZZSt4xPgi5ve
6zPqkZfn//b2Q/Jxx6cVkxKu0BBwd66ixsGCpa1yQsejBDSH1EIrEOSbWZNTrTDOZu8mbgNW5lr6
JLmh00UzETL68K32NpZCin+3zqwbPLVfARHOhQskv8VNFawxKPYC3d/tgP/flzBrKFQO3oXYdoD8
BWSBTNqg5SWrGp+JG1b+o96aY2TLGYcaYoxRorNRdFKT5+rYOtxJl40dob6WV2ErH92ePUuQupXs
3g5xyh+Mfe43K/DbtBwunbLGfhQ4/0gldTXQZrn+F1QcSKg2ch0JztyP04Hqwt0vdKOUBIzLyPgn
7+f+Q6Kap3p9Ym9P/qXq2XKW1oaCd9E8oSWWTYfUCo7DDSLIHAD2Tr2/NzrvsTlqERMq/g0roZDH
CiHIiSf3l/zJCVsisCdTOd68qOfy/xgrPBHn0z06iuLB/X1syoYQSTenNVw/i/+zyWVL9G5Pm14Q
yRidWNWYLdWdDtdk7a9uOZ9oTrGBL/5bk8eIRHkHr991WpxvlJBkNvaVd2S2EBJ2ZWx7NcXBVRvs
dVdghD9inQP0Hvg4nleJGQ1iU2cdw33A7z0YXU75zbeM5CPpe41SLiVbTqPGGFYH1DFVR54AyDgk
3DGTyYEdS52QhtERMX0ROrm5/KWWdn27VVJq2fGBtPsB1HnHDfHIn0vnw/Pax9DprXgBV++9Ncxk
fAwrHo+XFsWjcViE9i1ySx1wUq/S4VUeeSFpAHStMFizd1fkieWrg2jB7Mk6ZmtRdbnhk/yShNqq
BvUdRa72VgwvekHgnK3ihvLNwy6ZGY6Zt4OHyotEeU/QCAO6oz+suT/k5Q5M58W9gTWBKbPaRQiL
UQgcRR08/P71P9FP3Xj7LsPKlt/30w+/gqjz0ukpauXc+Pj7Y9ysk9FUNE33AJhjLTemx/1vf6Jy
cosR3uo48rggnIyHnkHM6FAwkF20HIDdldHGrq5myAO+zA4OmtMuXUvUIHYFVTFyJjDFAwWjAebB
yaIUMGEpR/xxHv2bDByjar+id2CfxfCU5GuQus/LRSiIexH9Fn0dqC8BL+003pjQwxSWpkBE22mp
IvsvkjqhgaBuWgrQnku1eg/7PCvzFmG2QmE4up7Njb3snrfrp2eTnP3te8tg8tnEVSvAKU05Ca/+
30UDsF4QYAnwJZAhUlQjYIasUxH5G/D++6qFIaF6JpYxhHgCAV8GyZ1L2bW3V55DUYOxKcjJDYVV
9hVqGQpb6D82tJLF10ltGZ3stYo5xpZtNwUtHfeQn4wUX1dPyKABCY8d5B/R+FIikHuI7pTAEKlL
xN5PYsl0mtVHx7+B0H42tXODLOnCrCfasZq91uM3U3ljxruBKYjYScSbkFXDlWeLEgQbIy4cJ6Ac
CXeNdqb036Pw5pxbY4dtH/2Nd13xXO0gBSwhG37dNFYaWSjCCkt8tP5ZtjNFeUEkYnwRqP/ohgZq
AJ+iKmgrNrd/SYjnTNuWcGz5puDu9Z5uStZSCtyrNTobq4YdReNwtDif8kYJEyStcdh2ePTS/xch
YD+/aJ2mzc/mchnD9NY8PqtHTQG405M/Yg/3WLfhNr3asd5kvD9m+7nciax/YOmV2ckJdYBEXqld
gSFAfZSyxtCI0UVqiuzgMqaNsX8bcQsspyO56C7FQEWzexa75IWRpIurY5Mk22KSAVtH0/Y7Z93j
erbSeVFfnoYO1djh//n7gN62r6dKPYTvIiW0CEx0KBLf3md1wFR8GC+7ok9zGGBAgvAL2mJqIpqC
n3Eed9r26UEduQ8Kqcka+Z3OZENZqRfM2ceI1sk+SVTWv63rVD3RwfohtJwBWCDUiNG7a45A/QsY
BWSQkSh9B/sEKmzkplWtKUyyPliT/mSmFD1OKtpTNoiHAiqP7I7rmyB5V4PWSBWYrNE5KWT/pK79
KC4CVjjnePV5BhkyEn4xhI1y0bHNotN60ZpyHaOyn9G71WqaF12Fbbtc8ca1P8JxFyX2oyI660k7
Ek0XtTyi9y4fb/m1t27I26gZzFiDmNuvO4+mT5nNPyeBnRJ9tZ6Gmuhq0PpT3lZ1IOT9kTfDwtjK
XsgutvCgORIwTx5d9V4md33g9I8apq0cAxJLhaM/a5jc44VzinlzjizTye9Edruh0vkXT/A51nOk
KRFlNadyjpMRKyaivj5yeLArYtwbFZ2JGpjUgCYYVjRbrdAoE2uZLiTlhN0pQ/XQAPElLpWDohPB
2Sd81RE4N+b8iDj3XRwRQNWuhVbk9YgGADP5K0JHgrxAIbDOrxQsHPo3cBPaexXh1OS6l0LUnpmb
V0SBtoit4TVp5DdAYwQk6xNntX9hSj0u3R3KMDkoB+x17osHCzLzsFcvIwmSYiRANeODMvms2nQU
7OxRajECClzUaUUZobzOqSzLf0pXoRhQ9JN7qBgouVTJFRfGGe2XnzjuDmHjJdtiKkLSnItqflNI
ic9QbSLUp5qfeUI1Bcbe02NXL5jB6iOFf+XK35PspjmDNBF6cdLDA1WamLV5pWHjqL8iNfLXkSSO
QL4CMr3sqoyjbcNGPJmEWdpZlLzgUozWUWh7FVmXyk7egY0rT0MGGTObYeK+tFMVP7zRZGGlD4A6
Bd473I3+CKepqpNKrKDqAlcSjIzOcDI5B3O98zfghVLr4be0EixnkmLj58lgeVFldaqmotf3ayfC
WSgyEQBKg09EoEA4IRTNos2jHWH+/+wRFkQOgaMgGPS/s4WdZCEyKYIzDQlnJf1UfrxtYMf+ebca
UDu7o/El3KtE1rhN8vmf6WgGMVmWPQTD4C/4+4DNSixBNo0TwzLhVKh80grm67yuMAc1MlvIOrjk
dQSCfxTE34/RGeEmMpBbLP4O13g4TUFJS/hY1ITSNfIA/ufD8bXDghYHD0rM/Uw2fhogXZrwi0iq
fPUO6/lboYAl8wj1C6sGtn5aDW0Qf3o7+cANw9HTCjIX6SwhBmB/iDoXjdf8/ZYEw2hWA4PxHqpT
LFDTnlbQzCUbgnr4LBSY/Jm3/I/JiV3rmT6EeR4YNziyRZ2yue/pD8MhOXEYk1bwoyykl7JxFXpS
xRhsDmVNbUVL7thZFI1ly3Wp5a5zdky6ckn2YEu2xbj/RYtXVi4Fl2XZGQyt3MZJToScgB/j25Me
4IhUrXDcMqmfs+88+aFHnh6XChI0WZVxK+6k/R1VeqpGurIbQWpyuXAJW1Nz+l+MToqFZPWowEan
sjbXn7P1E4e8FSio+A3xj0kSbMwXA8aZ7ZXndFHUKkBHp94MN1HUR25HZVNeFdyBoXT3A1NYc/Mq
0tQncwRVf7nXtDe1gAZuDUTWIHor64aRvxfkpNqou1lrAu/l/2DbCxj+0WOnUQbXr/VUQRTGIfIs
CvR1kGmKJX5YoG3Xz4zWZAg5PeIk+Ac0ZueZzwo8Jjn+2qKWvlXvjNBJV23iqPpeNqLo6qrdx1T7
5tghkFDn2JHRKShHY/QTYNELzxqEq6UIs/0r1BYapv3zl+gEamHmVbxmWxvq40xgjHitVuay7krw
iQ0aSM4a1rrc2IxXDUqP4QJz5MuHNiijjweciqSEccXwqrpCkIK7ulabVghBAlayYCy7zhQmLe7G
3mSQ9rPbpaA2M4TLkJ4XDD3d75Hl5eU8ZSAh1RDKyrJyt1zFeChvJyCn++HaABeWwajq01bKj8Zv
Ij3pvsGTZ9GlZym42SvNKPuaXwqnLgWzdfj+blSj6iWpdneuyBH+3fQ1RrcNcIzXdBH8NWYHhm2y
grwv7n98ZaXIqGiD83wQkS0mUn9Lsj/W4LMmul5+N3Yq3fmMpN9rYPB0C1wjRqDWc/h60a/f9lt0
zv+Vhm+HeEBcf/x6Vkj2Co7N1OCqCmbG5nrKhAek1kaF9+jSEvoI3Qh9XkFGvah7G6SaVNxk5dFp
xL+AhMbZDYcHNPdrlZohB+Hr4Ib3+IGGn5+4/ve1pciPhi8B2FMggQMlOsPId0++K3pC09BVkAm7
Z/mNY714FKrJZFUSjYxXNs3iWyNr8Fv0Ff24CEErJnEsJTMm8Sy+hU4cZX1AxCXVI2/y9dOARKor
cdGZx5ccKTwYhV8irRt9fE+gfaJRMVvZqRl7Fqf0G6VF4pCGTG0RtgNZeuAGlwd6y5UISeXQreq6
xB+ZgG+l9apK2exT8VDRqigP5pstd8tRMmClkzo7IV2rd1c9mBLqRJMhSzampcxwIPpu8WigKnr6
gHPV+QFebuIZe0QOQw3ZFh6kV8pNmqRo7UuG97gDgW1Q7Ai03qvcMXh/Y3jTXTFFmFxWEV73dtKj
DqmoOREgFUyd0kXeLkzCARiIumxPKokawaIurR1pIeKogPylQLvjnAyMDKjzxHzTpL3Ct0pBfUvt
m5404RW2tYG273JIc8eXQWiE2ofQ/l8o/ylYT0JLz+Isqh3tqjltZRRKCQwD/lGRcwvLVchRYoeW
1580zvmXRNLioRZ2BNzECXE3n2thp4dA4XyUQ/5/uQ0oqzY9gFTA7qtdaQW9CDNv6ycfc2PxJf4P
9IpG2lTTIB7G8/fKnJku7LdI8IyaApFMkjWRR5Fdq5mJo2VV16m8TgCHTiUKPwUklcwlCLF2OmTJ
rhBfqGlQJjco7s89QNZuftvtJf0P3mtCurtK9CrctUiJ9GmxASOU99NKbeX6D99nXIpMI9gE7xwZ
QVfmHmb2zsbD9cYe6PLJr5BTDMby0eW/K/qN6A5k6mtKKs8dXrF7CmJrVZNrLBeAKfpjqcU9FnrI
nloaTwBd3rcVRs9fXYxtXOna4AX+ADbrjjyf7Tvic3Jb3pRH2J0SzYL/ml3wXasZPDLwf3AN2ShA
gi8BckldvZc8k/3jGr9+fu5/QPPaJerGv5Mp7Xj8p+eHhvG+o9GvjgmU5IM7wCP218hQx+s1Gaun
s1kz8Twj/kTSD/bPsVMmXn49v/LaUf+kvddcecHLD1qX1mW26M7xXvP/CeNklF52liRSmZE+O/1R
EvRyHDCRsCxEnIQPnpgzt53WEZ7OeAS8kLkDehTKUO/WItJVN5PrsH0HvEX8pQa1xNDvr74xb1Io
8jb75Y5CFPexVip31MYp4vVkXTCilU3KvDJcTbhh75/0sgsDTobJ1I2PYi7ury3FLr5Qto4P3KUK
uGwlATWK1HuDlI0cimuuhI2qMnp8trs6Yt3VYYHeQZDV3pLNrCXbDUJbOdc8rm9xa3FFAOoQb4Qq
cNfV11+d0jIxUA1WDe31o4MnREaGFVpfSmrvvmA2IygP33RvCW72oMIkMaQrW1g7IgRWyfdz5iq1
p6HeNgynKmWMzItSN+BIllidfaOEK+p1svMjcm0I6qyuV5mqVCkT1akkr1eiSFBRWFG9jfbN1fzL
gXnnSwY6Pk8HISZTxIh8dnVrqqz/ytiwZlmTYAn+y4VPqyMNViNG7GpwiDKdwJOaRZ7ZzqkztmRe
+gtsCwsAm2RInQWIrukPlWC5xHes5OTRhmjyOIzFlkVK0nHJKDf2SI/Ui8yb2Y7OHPlmwje/k11Q
OWba2mKp7tukQP6eAS0PVyu3kgKclD0Erk4M9uYkuFPAE302uZgD2zM/WKtavYzde9L0RJJUtjJ4
Lr22njBxYt4mUnCzRq3QakUk1zFcSrWeODIqlk44YkKCzLM+ZiqWPyHrWGGSuHBg/u0efmt8M45E
6L2qhGXkt6a3t0Rslq/EHpy4J61Y7sv1wNb8NXiQIJXvXZtG3iAUlgJaeTvUaddL1xk8s7vXa2L5
mShXBrNNecDrkcRbMJFpNkbJUjhkZpn70ARmS5wFLhojHDDRHsiAmS18Sl39c7qILPWL52rvKHMG
4PiRAakQJIQ51/1ghlHv325H59LeR2/7ExgS8FEffK/euxpXYthTx/N/phtdJZ4lAemr/EDhB+Vy
ICfGmI9sbJCK4EPST9PCIPbXDO+QHs2pVPmadURygHAOOSzTxTjdbCY+3aFwKAdY2py8qTJcaUKd
it0uyURu/NI47IeuLhuaq0IFDhXnJy4veBi4qzIco8VdIjPwk6XxDoeVmFfYG1+XVeKdZCrCnGJN
S/6uYBu1eJHE69tkZEnjjdjMiUXAmhyRpPt+8S8mEqL7xMTKE7BY+uxcoAg21L/mZn6nn3DPHyJ8
HExCsz+ksQN9BIM8FnbVrawFtXtZwruUOKWykWeXC0NGGVnDBEotCgpCjLXjFlkt36po9ER6Kjux
hsAje4cV6gC6p1vf7Jj4qU8iz8iBFx/HOvBgwXypGFNuHrV8HrcG0h1dsRp18GhIVtdD55Khs/aX
NenXJIxbOMa8eWx6IxWTNPTk8KA4MnpJhuv0qaEJ+Uh9VPz5fm4Kcdb28EkkAn21Gk15ByW/NnfE
bgZjohDFtKnK+JyGbljUmIAEE29LnHfre8PcmtNGQFrKtQZDOAy7YM9SCowmDfjLe2r4g0v0K6MA
8H1WwHfYuO4yY++alnwaczF5wiwmE9ZleaVmFZM/GZcyT+AMkaEbpusQgbkLOXH/d4riGPtqpB+c
rRX4zmpT9GHlWpxAsRGa5IKFz/cyCT3kpoev/KWOwVDv4RXDEGOrR1brqAJjHNg/qsalfdoewIyj
rRYscVvZiFLdg776T4+qqX1G/qPqjcg6te816GTXmbXT5WzToj2GiwwrSzXKRi6mQ8HBWzSzmvwJ
+cya5qTcAfbZT/CoM2tlgofpQPkhTs6rbxjnNvvoviS92f+iGK9uBLaboOKg+HVhB/A4jPCvxAG9
za0UE/IizJlhK8zuGBjItRTkZtim56JN4pk8YkeE70GV8R6Vy/uxazagTN6XutpNfsJq9IMhRX+u
5MzsaitT3wdThK6j9ZTaVUkPFRMQ4YhjxFKHSOOB3iD3yyS8Rg9rbHRZd6p+tcHLAmq0g+8OutFV
kzwt153/A7AMi6kk5taRvwj4IFsdGQFZYIrOiMtKKTXlAXUNQBb+8c9xL/IvznBuwSMjZnCH+v1Q
hea4yYSWFGBMax6vwK0nhQT1WsjQwcltHlB0jjUfkEwCjepvs3AQKmfFWDrzQByM4zt1QSiD+bIj
SuvRO4uTbWrgS/wSvC/Pi5NgAO+1tPMlBFs78M2MQ+jv6Q3qdA7tkuSQLnrdcLL6C9N5CXD2qRwQ
0neAL4VpnnEEgHhnvj0kDC6Jnnww/4c2asdD/KuA+LGfAZz3IwvHO71KsTJF7gCkQL4XfbMXL2ht
4Yl3VyrF+IEv9BuDElOZNEWyKPJ/tI2j49ldj3T0Z8OBBuHqu9RFc1rLlQZdDvykgo7fk64aBd7Q
Z0cKnvDZrfeXt90aVg6eA+MFiQXUw1ZuZkSFYbdRrzLxY0qh/B/Tzrt7tB1Z1gomJ1/RmrLPLJm4
NbHvGydhiByBOSgDGNY5/DoWyk9RxzIPOipM7KQuIritZEF6sd1uYKW2+ckZ0zO4Vq5n0RCcA1Zt
sq9PXub+Cj1nXAWY0SL05yqv5PT3+xdhcLqsMG7fdqROl5ngBcLqNvm40mTjPDN3eloqdkFBADUk
fI9dkVckfacslpjP8n80qb5QPpZkraKPCFsfmmAEKOR+quoOcEoDHVg58Jxw7x+9+zYHGlK4RGvS
ejWk4FbVO+Tm+jozswXidf6aK/ZIVHxfc1HuqawLIwlHEBXv9wpYktv125cxt6IeDKPDl02K4dPp
8ZGm2B7/le7HeXqnda9kPf6f8kJtfwAk8GfVU8xhT1rkBUzy8hfIKlkIJbusF/aK94uCz4RBGCvx
qHWDeMOgCTzcU2UhAmBzaGUHzf0jIQeJQ0GbpNhuyMfynYQeI8ffV68e6wTMB1FsYiB9fJyvtG5b
cq8jbTsk2GilSpbpcbkSoCxbqFUkkdupyuv0QNHUY1USJlnPz/1nmgD5OpInETFhTlhXZc1wImEg
p8yAIUYOh0yUxoMxus8KolH6TaE9fVkUlcvZasFUWja9Z/4DkL6y76g36vk0XYv0YLFnVB1/hjuO
KHqTm3oNMxXeqJTdxw+ByB95k43r9XVu1TS+97HW0+dPCQ/Kr3TMeaU/YBZ5iiCklcPHbDf3+80g
G8s+two6zwv1KbvHKKdtAjeeykLMzDXzGWt2HxhQDqm4hedGRMr2UqyfGaspcOTwapndaWIK6dMi
QNdC6eyv7esVtUqOuQRHTZoFZhcTIH0YkYi4SvRvVXh3WTUuJUFdp0xnrA3w4yg+7NYoPSjOuOow
KWDU1nqiSGrW6eQzHOzQbU+61k68OtbhGs7WoVkcWmFSle0aMyIgmibvx81xKhCJta1Z6cZKikZD
BIVbHPRdkt0Fur/B0f/pm9+cxVVACwFMzgwugFrRlkVj6R5uTJirKf3U86qUkbSj+n1SoaWxQauE
EDah5WzHcW1pPqas3dqoE53n4ef7YDfJpndyqI8BDA6qFJbwtlpsrwgF3UvLLOOKGihAkunkWw0u
s3Vg2W8NBLYAEGi/zm5XSr9jP6+jK0auq7tpu5Q3mFrKoj93+j8N0BuAPgif6cHkPcvYEh6B8l5I
BpaTPV8n+xJbQa9PsE3WL0W/NOWW8WpWtdqfVTdONR+oy9BGqbaxh9Fe9UlFXcsGB5+xmGeUKjM/
+FNNTuC4k0aFGTv0KC8ogIq8dwEykvb43fE1epai/ISkPuoP01cGB5pUWJkNtWoBA+cmOIFpNzMM
lZrqe7MU+fbubHy8IqqiNRihwsDhQj58/MGqejHdEpTLGAQkfQwpaG6g1JgYW+nlQRqMDIN7JTLi
IDeAujRft9FEGmui6Fx2Oo77frR9pPneLHHnVTgqBR2c3jPpGHs2MfB9cRFOfDPG3J+6ecugZB+6
L6xaeIrsCMDg9gmcCXr40v8enNmPHqbUVI7CgSJgE+MmF36siTcYDIr4xa+UYcS/CLL4GI26EP+1
mz1IH8+v723UMk6LprBa6vgWokZ5RQb+YOHMVpMP60fB3Lrwcr2Hpwrz98jPBfkz8HKXOLj8KSQq
LgG+Y8wAPV9BSvMGrd3r6tpuB+dS2rlANIrrrXXJOme4/odHeNKoaj/ctO5yE+JMOBxrZRHg+FCV
F7gjwEX93Ir4rjlvNfdreSrP0jQ8r8LMt9TPIkf4rpC0AUQI2Uq1miKbCeL8mv6Kpsmg+FpCKMaQ
1ROioUHvXW3vliWD7CZch3IOQzIQ53JBTFCHujBVNtPyWEwpJ9g4icnSWAg46x6lbmoZJMROsFd3
vKo176BnjXcqZMo4ndrl2KGOxsbIv6Z6FhkNbx2QqFfLOu2DfSKuP9VX8dSxskhUUN/b4G4Noc5b
RCwHLeF2SazDVV1hDELBZRfHa+jmfHSgBXvIE9xJ2UpYwn7RhhOPnba3RhIJ8aAPx5/Lkdp0htZu
NUn8gba/gL2V3x3GqffySd8inplE01yxOS5FE3fSM+Sehc+XqkOY7N+eeNTCCvtG5TdvUweQqSw2
e40949uqzwxPU/5QSOED14+wIaVmUSF5VjVD3QoLPUcuLpA4w0ccka3xWa3tY6dtg4p+BXjbqKMj
2ItzI1ijUbftLRgUdnQehWwYtNucjAGXcWibN+e0DcFAlJ6PdTyOCJgwySzdIz/Hlm0IHiTAoL99
M9c4LWyKBv6SyPkR9Ky6TU278spVE/wDrEfvnNTH4gqdSxyb7jU/N5awDT+TH5acvTvtTxsTbCno
MiaO53sTQVuu288qB1o+1+U5bv59dOOvw+EZ2Sc8FZg6szYLo6pTsFHDynz45J9Gy+LyHZhTl3/B
htIHIqB56VuAr+/v5Hb6iUwPf/g/3YamyD5GHPQYDSJTK1tdiH+cFu9sos8ZmzgU6MWPYUHReQM2
GPbbI20odN81w/2o6r4oBLr6q2iWpG13FojpWCpM+omf06G0cT1fXPtwayZjl3DQk64FoPWMq136
mWCfvgmcfgMfVsOneqHxrs5MIT/JvPf3byWZdV+97JMRHv8R20h0K071BWXDUPjlf02XLsIMq9qh
4X81tEAxZgXxC4fsN5fviYzCS5AhoglsXc8ViVUfOJ80kmAXfat56r1o33HyyQ2bxkf+NHtNBJ7n
/pgmmq8mRv1Jzp5J7l6ooicfUiXbmLMzylJANmO2l3icJU7RkNa4Wj3dfkps5vn2bQQjp0mUqaY2
5UznHJDPNLcZvmGPnwSSzCAOJlRLpHIhqFlc0t8GfR2pSQZP4sRKI3MZ92i4+2wUXnLSrgbOwyQL
x6UdwUtANSKUIBWZvx6iR1NBwj0xtwunksN1edaehF+sRTtmTGPfHkNPEe5n3iGo6SbZDVR+st3t
NQYriY6237c6GQl8UKUjgh7D8B3YE0cFaA5EdKcXB1WqQnJklOqToa/JJ70gxqnS9elIXpUd4Vmk
uN/6kNFAPmY9Qbb7K7RCZTkYepuQRGQH4WK2g3vr28HtWBBlkW9bQj3l9IOce0IOcnb1jwVsIDrV
GFP84I65w7rNwKPLVhRCCkHxcd4xm0qWi6TY9mGbx1HC1K1m33AkKHvgzaIcYVk1CUox5oSJU0XM
AsJ9UfxcmOFfh/bZAP9y+j0tHHo9mWOJOy4Eisk6hmMpUlJTVSYOKlDJt7bVF2+LrATHnOayuINY
QVN6xu/Rc+xD/8gfePHJArspG+eHT+sduM4UsZdOmI+PyAjMb+gvgPnO4Uu6aDlDbfzReVaROVF1
Nd1BaxMP7NiUenSdtArIGgerdISOS/yg0xuAKI0AkBVKuOEn5NMvWtC7bLUVWBTLKo8RVXVqsHAr
f9uitHt1KPmgR0x9rvugp87w927fmVDejD89ryy3GII8NGtaikaNe9oRwkNQsiejD4RVDVB43oN5
b3esmvgpd4mNzXvn4BgHcCYP/8OYlQG2JR2IMZLB51SF2SKfgUuaa07XsemOTBWZQGeuEcKitad+
8K0q0iyflOzyKdQmyXG7MDamsZ+UHZDBg0264uk8ovQH3u6ZVQPhQOS1GRMS/X6u9Hxb6KR1ysJc
5wGFduuBo2/ompY1UrQSmM5uE28DPYkUTs0yoqO9UwRY70ZAvfAd3Ogzz1FweAT9D2gqPsPL20HQ
WHBZjYxO4fLnHasSdwOmOY2y97XzmlUB75OFYAh/vqyVAzKeCTmbh0CVmO3sVWUmUy0ERk1brmDr
BATOl29fvaT2YaseEeLg6fvBQ4CbhtbTroYgVWeW2WyiI8VQVl94v7m3iBEmHeRDcBdmCkbOUMB2
AqitqiVeHPoobenpwfUiPerP1gMjXRq8uKr2oFWiGYeUEJVY/pKxWR2G7ovFbLuqgGjl5uj7Ya3G
t5asu8UOOL4xzZ+OVdv8yN1UZiIP5X/BWu+AKQzzzZWEqszPe2eJFXlwI+OujCejbFh3uNsjH/8I
UstJQXy2tEYvvMn/3B9ArBSNUWTvzBdI0bTkF1KCvDpXFaIPgvJkP6RMiQRDMPxACq+1YLjEpK5X
4H+1hbOEEkfhHWHe939pdq2JT1uPf+bH9CNjczgyLCiPl48Iu5v6CcD0pE2g635qENYDCzeXTZYj
fVo4/tr+7+kmGSaQmhazatCcZIvUg/aq0yPL1J/Z2/V7ogpWpqSJ79tsYtHrgTH5GKAz9UqGKEKD
xAuU/3zjxYwR+6mps2KeHMVyP7NH+tAGkYn9iMuSdsU7GLIc2Xx+ybWFxUxp2dYNy6CFLIkNiC5z
rnvU5HH1QpirxLndbBYeAiia3nREjTEiP5hUnnbb15LbTz+16pnHMc3I4MTIeRQGgn+40qfAJ8Za
UdWEimnbtWBKJYU7U12pwxBQ2xxGwkORAV5JtvwJMl7rS7EkByNx5LjGjtU5oCTeRnvesLrp5REA
3yxD36vk9KDTkIUPsSn90YYJec2tz+Xtjp7+LND3ojnKQbJPncUGUbuIy1ifuINSJS/kNN1+eWsY
tZ13Jb2HWdwutwdgT5fA2FylSadHDE2jUF84QgQOThRBRLuLgplhz17rHptbLGsybGBXFYK9vPdg
le8twcfXobxLZdnIA6ynEvisv3LxlsIshjJ2/3mgb6B7XY+0RVR89zGnfEWq2Ss7ir90ISlSuOK1
XWa4E+UOr75Bfcgjlt7syi6oqLfqz7APP6+8cDMEg4rfzoyGvjl9+ltKEHrYLUEhaBwxeg6pYoFH
pj16RhjEzLRVV3l0+fHm1o+344kFFIc6HrPWWjCQ3CbeOKbzfqGi3YxoLdqPCorYzqnarkmFQDc6
ouSX9cu+mDYZ4IIqgih6qhGW53rTbmIrkTVSF2xvsiGDF3/I9dT/tj9cJCFsWuH13pvw3mOHevTr
iuAC9nRvgc0PQYVkSdef1bu+VsTK5oZnV73shy1MgH5kxKY5UhO5fUJLN5YjQP2qiLpEnZHWWODf
EBdMRJuy8Wz8Zj99mrVq4YNbfxgrPXxpLLwvMJuTgvIjDMYlg/+JTW3ysH+FT7G3NhQpOjGZViOk
YP3MtSg526mxVc2ppSB/4KYfiomtuYxMVmLATSNH+tzuD59QntouZr9pnlMFUmbyc8pzhsHQuFlf
uWgusg6BxXWc579J0GP0cp2O5L+pmg323GYCBF+5JNeZp7jwGYsjlAB6OJmGtyOHe+EmDnYgs610
Rv5g1dkkfYOmpfnmmI7MltNTv/938O2iPGtmTGVBuFCcACbl2cymA0Yngy3/3hf1WqrYsffbmrUy
uF2tFlXwzJl+0Tws5tW/mUyGLL3BEF/BT8MFuY78mbAewk52+wOIrk06t2ZWmnUHEG8a16AjaHM7
t4EEWvSmTLKn6E2hBImrx0l/TXy/YNxVAWHLRRVx99Nr2U5U0duXfBhXZliWpQwPityvFxhN2RDc
dS0T8JbKptp49EAEEwA+fIuvtQ/GRQ/rNksd3Bf6BHdt1KUPoNk7H+fwWnOG1GBbLwUgXNCgmMY+
Myc0Pn7QVaOCx5BNoemuicnbtzlBqsL8sdbXBLrvlPXlf9lZK81tvfEw7Pp4lUlPaZf+jH8F+LTQ
8CvBizFKZR+egpnvYwyQOiiewD1VeksrEvTVsXgfrKxSX6DspfGWXgU93feND4labq6ubMPpIsZB
SLSLligJZzaLMIbQI6vYqpkY5NUTe9NHt7mffw35F0f3otNEZWziyBWmaz028Oe02F8vxZLOfV/y
/ZGpApurLXHesIm4EO/fw0NhAZ85hz6deIU89VBqi5k+RdeKGlV8ZbKNlUxBsoanylXTYVHwGbH6
B/Enqq7OZXV0uekmrLesAQu3HOr1eA+432bKdPqI9UiAfZVC37f+BHMftvZ5SKCoN09cndXgG3ai
Bh0fUvY7RuEY6WVluRAVBimVWATjs/A/cu0xNRmuYaCkN7+8f2deFX4VvSAeTIpgg///TUTDTPgt
cKZEaAmKie/tBQTaf9zglSrViLagRIuVOPzYcj7Uns6D+bagh7nhmJF/8CdQ2aY7LnTJC5x0gBCF
axsrqMGZXpl8eJimHV/Yt7vUTDkzKcnGR2G/vwPbeqYTW8syADLEy+PbHkCxc8ZublAFz37a6DJ1
JkNu9Ae0F+a2B6Fh5UqUeOckliASLRL3ujwhidNnD/AfW9v40F6HemXvx7PkOyT/akUmMQxW/pAe
fP8Phgx497M9nDsLKvwEiHbH1zV2/OAAWvLZheLP/Qt/nUGBBku/56CvptQFVJtXlue652bksWT5
5ESWUTVeYO3zha7KunxmL9Cya8V3CqtGU45YL5A/b+1iGjGnskgnug6l3F/ZZZVjeeLlbR14XLS4
UIatJ6accecB3r6FnkSXyb3NomEPxg/wE0rWhnjefGZmb/AEL7A2ZRMVG+5ItTS4G6o0j0BD5rbl
sE0d0jUIWlyNADwufAR9fqkX0RSnKLHkB/wSjJ3PQnB82tya4D2iZJr+zoTv9vJeV6ptYeeiMwPs
zkWVQ2McBNr9auF7TRf/MykS+VZGhOzImyPZfVDQ//tD98u2Fd2NATLBKNr2nFkU/mHmE4sQy52I
XIq5o5OQx7XLvmoAmhA5w/A9SgzxkFKUtd7AhKhkKtdV3fb+54ZGAtkDCSXbGVJ5hALOQudY9WBc
0tqPcZjFWNpwj+9/B975maCs1WRIX+4h6eE3oLWBqU1TkC8geYmuvdRnQahqZ9XXk/6zbz6HO8G3
d23vTJncFma9Ooc2thguMnLU6FavkgbvEePQZ5tHdP/KyOR+eFQYe1sY6L0NNT2NovqdIKL7HlLQ
aiHWlb7tnHNptwoHhlkuf9UIX6B8QzbBJA1G0zU5G4CIKT5EIBYRpGhWEIaAwHWHSV3ms71booA5
tbxjPnitQn4K4oqlf0UKvmlAsLXfr/8SIQm56h/39c7hn4+OXsKt2HDCOR0Qo6ePzAksq2NlD4KK
B7XSynaOkbfV3GYjHFptewMSWHRsikitZ10qlarMVLTC4wOdE+FydUTZzO+sjDxA4yHAVOnPyB+s
KB+T9n2hfzv1AYdkNfCIDjBzEBEgCRQriBVS7HFx7/Kxxiam90pYiqBe2rYJp5hyi1uvnbcCgsi8
x3qiI2bIYhM7hUzBBz86MxjQTMHw+M8werZfDG/D+wM4gOKCFmpIvdDRRqxKaDLq/pHAy+GFtMQt
vW3YulLIQVnIWgby+BaXOYaQ6/OWUAhgQ8bgMIzvKK5coMDES4zLO9bQ4HQdXGxMQotdERI/ZWIA
ZnPUV6/kTrY+FlfwExQGtXupNErMTFEAGB7GZvAAezrzD1wXPi4dFULNTBEOf3UvVVbdaYWeg6aM
TvZ/53avsmrC0gEzlBf/3hRNalPtxY/fgbUwIsRUdPzH/a4r4pl+ixgmXMV9bEXYDflHG0T7PaTJ
wnDAwlc5AwMEzR9Lqo3oyTvNPKlplqye8Y2SZdmH7xgmma6cgotC9c8/p6jsnL+ahnV2AL3mksBY
sCOOeinWWHzF1Qt4u4g6RPHA2feTc64LVqRQOqFImozimwA2dU7U675P/Aded3MZC8znxgXcqgF+
VQW6TX42Z2MZmGB2lOH2qq/01KFoBOkIIoJuprxc96OcKXH/ko8wZuoXTz5Dh1XEY/LMmbsQw2P4
Z0xNe+9acy2fVW3y/V8pmSgjB6E5NHnB0cZYjvm1AIlK95nhq0Va6OUf6aD90LZjPxH2gUTang/d
8A5XiHA9S/Sbz47nHserxRM0KXZrjOrwJQ0krIKOWBPD3ObFIdLseG1mkv0zDqPpIM0sPmyRI02m
sChz0w0ZeH60wqQz2kpPqC+RFfp8vrsUB3fKnYRUP/hhnK+sSryMhK20ucKXHJ2mij5S86N24bm3
GzLIA9TimrlAfciac2jsP7n8ankd+hE/jIQROf17sX68pl3qS65ySA7J8CNQu/9UHW48NfjvkJmK
eUdHIEVusC0akB8Ca8IiFeHxQfioDFsQ5swZbU36MWRpQYZDL5UPIluQI/zlbTm1rLbB0izab707
UxOouCxSOSOar2O2OGJT2mzcKQwvjhGJUtQZlHlm1SuWHZ0MipTO+N9GsaoB7nq9wJ7BlkAuZDQx
GVKN+1MYzbLNhFumemQk6zDaAWVoiQVVGlWVnHvB/sfQP+MOT2Viz8Ys7a+IuxWEMnAhJ9gyMVVk
TGsWZuxinc886qPJduwChgfjBBvCTyjqxHJRMyuF2u0mcIpsLmce3Y4oj7u+1WXpa1iFW1jYZ0mq
Uie0iSPYoJNZZumQdZpUgMms5Er/AKhePOtRVfIREogs2djhgYQ9xssxDjl0yLFjQ9HAWtNJi9o6
z5v1GLJ19EfpqSoKIN7/ehAg/ZbLjfm6VilNU6hWKNqjGjfLRguEt1q75V5w9sxryT8/BpLDlnFA
HFbn0IMpIsmls09NSOWP/RDv4m0frcg3EgAOaNMaNI4YYqOocOg96s4QaN+qx4yXFUF7gR3BEugl
yFep7b1WbWI7BHBhajaNfCC2a1lqZ2qpx7bKfr4MZ83vZJk7f5pq+bsTH7WWLI1W6jTPVLT3WEQK
afpaZ0RmV041+0FOeoIKATRPiIVBtgjGpu1VajbXvDnWzEQZiAzePh5xikjjtfRQurN+1gOvSea/
pCdTrcinzbcnEBoD0ZPre0TPqtj8g+Y9UgvG9dYJp71PdNg4YqcQzgvDoECIZtVGhxiUI+EHdzWl
Aie9nBlPUR1skUKu4iPJEtO4bAJaxIrppNXOFo5yaCOuldirDCsvOHHi4U4tFKZemeF1ycVX20kh
NCnnGjWxjPANyEsL4nA/QJX4FuLsrNiCcdLfvRiDYl0iLl9jMd+uwmirq3+4UVyvaOMAG40qgxZF
N9N6sCp2bo9Njb48C0papOuV93pnufVVNv4mrhOv44P8xGEynJtQCuFY9hFYz2sW3Z+1Y/DD+L0L
Ao6G/iZLSAwkoqrygZza9A2d8Kll2YXCGwa/ybEWsDJAV3dNuksghDN/+PbKCkWN2m/GoV4XPG4h
jShxO99woNZ/0xgHEikj4MCXe/mQq2uSRW0G6w6ptaQBzc74GhSy3jJjsBLNp9ZhOa85RnRrbWU1
LG6CiynPoObNnmBBTtPuIOuVnlH5qHR339uknUthTDrIbkBz+Njzg/EuBH/kcidHa2adCPFBzOFS
1rJXQpHY65YhF/jXZ+lC8Owl6q459mzauxmC4DFUI+k5clnWTl8uMEsQam8aOTelvA3UPJ7OKDVC
m2yUmTsTiPLf+aj4JpRaHOrHI+Ch7waTGgsR3A/nqzmvATDR3vwV/3ZD7YydJVEjRxAKWI8PDpBn
9LOKablZT+TAiIDVcU/pOmJ/9uTbD609nAdkfS5eOrdqZl4exyxqCpd5aFdEfTdpFtZQYi4UBRIp
4TImF4l8iFxYKlzth1LUCJGeIMMoS8dOf7ThDVuTdGiACYoMVOE7QrK1XxIEljncDY1o8Ad5L5z0
CtwpcFmH6CMymmB8vmbi8uGVWUCQDiW/rldppI7y6cJlKS2xqUMlE0WCc/j0iX/2Klzr+tUlNHZY
iunoWKcYtH1R8Xa0OUj5EFOQL+vmclq6BOUc0DdBu96Dd1vQjERxZD/7+ZHoGqYQkvS61UrHgr2P
8h1zm4ztfgnQ1rVgeqyW2P0JHUyejfInmA6qXOu/lmO2FlkGYsfqlnZoVyPW7LbARjfJE6chwu8I
RbfcobASQu4+ccHlSoJJ9w0eQHl4Kr11FPEdgBf2IoR4w/tF7+iPb3a360jQ1oOWFzgfOZ47dbfd
+8u02+RDIUSprxp9sUnHHgpY2oP4VL9MoNQZirvaxC47m9gakrNDPTv2r1YABQwRU9u+0OIbk+8y
QVNSRpcwuymL2vn3owGb5O6j20URGdYhAVzBf4C1Rlni0jfBuwZcLrZDxNzPPtAxramiZQqJLDXu
YaxDMueNl6pGNa7S9hGRoylBSedS5zLCnyvUa5/M8uapNa8ra8k0V+Gor232Xp6bAYBIdsjHu4Od
lq1pbKA/Qbh6l9FrTR6GSzPh6GJe9kcC2bDDfSXQOZZd4cDRqBfMNlq7sYsavMisHB0unyO63V8B
Ou25lf3LKvWEPH9RQjM4khNqMwE+pPcBgvhVzXibB6ihjUQtrRqWApW0L5eLh2E9EAY5lBFhH9T8
X6JbqAgeHAkpZs0tSqkHe9F/0JL/AyLuOKC8cWI7szThSG2aPDvTnIWcCr/+zE2eryo8tLlnXJTA
dzL+QzjO1k3hvI+RqyZzzt1nTSRDrzo7iP2K6a7aE6OpXd0lYtPRqNKJUrVFQjN2TxDW0zaSUnje
btzyC9x4ve9f4Jd8qID1Kk+LhUunT+3/XYrp+uw/0FFj9Sws+LNclunCWilvkPMe/BolSyiMAcHD
hiYe9LK0Hqwly+FCmbCJVy44e5afhujruT9i6azjZBnUkC8Pz0R3OqgV/eY3dD3Z7i3hhcfk6X3P
mbmsQnQ/+xG6u9YP7B4oHqTYOtA6jpBzaP8BzC480PvMckv0SE2+qfCQzfjo4TmjaoeqA74MZnmO
UYLOTvZ4ULZYUsy3uko/SaqFbCZEmd3XeB6sy2D6ALO84Ai0KyFNyvNO11EAU7u9Xne7FOoqOh1t
V140qvr/zFr2usqwwQlcrNqurt6qzyyr7a5Dq2evSQnRtPcZ+3WV+PDnqTA7mUYAJXfsA1Wsj2BT
iUo6O6ptKVq4g2LWnybg4Ul6s9cBUDqD3QpJyg2qIZojQiGOI75c30Tl9bwiNiosbLYqw4pb3OLp
i2tHl4mpE23iGl2irFjifJKnZXR8xH3Fs2/XvHyOJD494nS9xvT/bsVZpS17HH5P0gOTV905pL37
zUBvgg9Xh2K3Gkn6mJpPyOY0UeWoV7oKp/XxRGitAKH1KmliPytQGnitgCE+0l4E6mJZNK6Bf4lV
blujTwkV6cZMkU1ktY5IXj6+yUiJwR0rmD3lyDUzwV9XSttm3eGkxGUNWFJs5QmgmdR8HxRsnu5W
niltHuUlEof2NYQU3roAsdvsriJPGtcVbtkrsvJbI35dR38NeFa4f+P2Aw6FEMzwsiTAzNmQni5N
B395xWal7P6JSM4qrlYTmW3sZddcvXCs1FlBDE6giHbEsIfMthMUr+avvgZ0Q2hJNftIsOaM0koo
EivKM1hRg3Qfg+and/joZw8vEUEDZaeSE+/sOZzmB7hwTWYVvY7trNdc8ZJXJQ/gvE7NvrXkFhOb
kTFjjFWB2ZOTnUsg7npHzKCAhqxyc6VgLWCAg2bAl98uULWkOYxBrEqwf33bWxjCDgyRJZO3Rvqv
bzkcPj9fsQPZ2xnTTy0SEYsjRCtBHtup0lmJ01y2kBmHuWZcR09D+To3JPPddXBxkRlkW8jXC7qq
7jqdUA3pSzxiOR06KpT6QqGSX16yJtpjdzCCfEXNunPtNOZzLfgbxdqGjzqKx8iB/Qp+Ue8ORcoj
vVteHKxUremoiQ/1VJ5K0vv2GnF/5UQH4cP+z9OclGANcupZrgJNpSdrrs76keMMoJFx0Yvh9HKm
Nxpl/zn7qOKk9jY7SlEMzjr8cWEPToR1QfL6iy4+XCp/jg0x4L1wk/59gNx4H/Ouls2rcSyT3Ed1
7dXxc1Ewc1xnCFg3wRscH1A7NkyBwGL3QzPXF492w3daTFuSmSmdKBoMly8SNqZbZ0XOH3zVhebt
0H2dojOrYHabO86yToGXken3fJnEpCKNlEMCt6bEX0/xqewVlq1I8AmEaqOCDyZuuNgxekQMGTvR
rb5vPYrs3lLDtl1RH3QxepTgX3e9Zp0uh1AvdefJkSKh+Kiku+gxwwHdvJhKqJHFhr9JhkU+MbQj
YJ2rMvdnSg2N7vjjn8rnrj0ZYs7taCFTejkhcdwh1YVcf4nQRu2fZY63GXWxq2GvMCQCCEP2PuEP
6VVskN0ak7sLI2lyPbzQTyJYX11MTnPByQIwWFEqTrG+6TQmJczqVTeCVfl4Jvhoq6wQkKR+qUHY
ap/J7MEzQiB5G8AlG8t8Xsdiv1uC9w53TbeDIb/n2HcstFtSXELfIq60BBeTbxKQu0XAQRSIGWgL
jXth31/Hja3lGV+G70+OVwY0LdLAN96Dtq7onj7+0dqaXKkCBIjAwjJpiTGed4sbxvHTXjq/g3OW
aUiw+8/RU1TLSYYcrEgF/zZ6piUVpMcelozbRsD4w5VaaBAnlk2fq+mH9GmU794ez1hNPNdUo+pL
oY0s/RZnAs+pxHTIYh4nI810jTDrwO04SWWGTdnASIicFuVmPg10nMcNbHk8EL0QnFd5/iDPzJ4Z
N0RiBYBB+jWEDTy0ks8dtpD2mYNecr0ZMeX3MVkSFaY0Jrz4KZGL+BW0yMdsC3DoH3zhNcAXzrKx
Ifz3S6IjSMbxYD4TS0o4Woup4Ijb8LgRyht9usyTrCUBz6m6X2JR0ksp7iIKcRT2xMIVyGazOGcB
Y9cr8AKrzRcfn+OrG8gcVX1Rw5zClCd4Jc/cgFbNZeHeeIkNO7immFPl7AwUu/7qpYdcK1Qn7fE+
bKCtiM4yrdkxW/OvKrl9EIsh5w6uNL7M0+tFIjdtE3SdRKzKk8e8SeNYIu4TH6QD3a8gw4A+uhtB
UJJgyLX1K5wn878yXSCWhdifRuA3TIDewj51J3MC+/fVuZXUWr2Kv3aRUEdJnRXcqE9oRd4GQNlK
gCrqEkEjXjYKqIRAt+4c1lZgwYtcMlaBJwqnsXkPNdHvi3zVLdqOqf+NPbpsaxGB61hNd6RJxjBf
iQorcKHgt9MgY0vrV/L42urbvRjNSA/3j8gB/oeK82lP7yB+QLIWnIdH7qGMYWT1tbV0SN+3TiYP
DW8Tj3WWYx5xIwxkVSy+4IPtGtjbNqdPTWa7T//vEBmVz/GH8gxj9cp4/okZaxzfWb+xXhd11lhf
jqiYcWjk/wB0aiKq4uivMtf+tmOhJ54pa4LkrIEPDST9RI5gp0XhVIQND42iLj/CUfdJkVKBQE9k
OT1Kf5s4Ly2d1s3CkuDVkJPrZ2AeNqNtdhD0Z3678ad8Cqc88szgFOS+lwvrxGyyMQNPibGz+qP0
DOc6/nfnucVP+BwBmgzEkobdY7KIg/AgvSI3KRd5QvblkLeSDGRf2XZ7qFT96evDknhcYqc33gPk
MRvoUFaaRhYjqkpF0Ah0VDvDvS5MNk6G+3H0L2LQ4uRdDJ+oy/VYunRVcfLp4wkBlCFMceiBRxTy
ldo8nEIfbqZrsztAS/kuIcIt0k3Uyuwf1KmVYzslY4/zLh0+0ui9c93EeyixcbGNuw3tgrIJTc2F
mo1T5xmu2DDpriGPw+RlN/SfnyUtEPvFadJhRoP2AywuQeBAsASTA/Cfy0D8uCM5RyQpeGDp+ixD
wXyo1YtAT+VQF0PoszfL792SwQUcegyvcGoqLc4ZhbWVyYH6kWooW2AuXMF2JqCYJ+y+cILy6+5p
5yOpHh17oYWbVJcF2NCMktRIZ74HwbfWzL5+TxWe/THPCter2fzRGGEihHEg76A3E1tgVt44wpMn
ujfUQy1467Gob0YjNZ2CbSwu6ql2d5LBihBi6l02FB6jmTcTwBwhPTn3d6oKWzzROgv56inmyAvU
QYwS1Nv4In8jKoJksvGV3osN0EXQBgchki/kuD/3gWaFWcFS3iW2DuV6RneW/wbWCGEaoz9jXpDH
mdIakYrnnlQQ//GJ8ZEICrT55GPIEY4sbZpkDYT9YQG1KrgEa4iozp42VN/89aMD3zIvgUkVCghC
VBKTdvaykopc7uVuP7RkAtSspiOlsD7dNID+uavg58Ssk00WBXW5ilZlIYuVjgZA26rdKQOsjiHx
ux9pFdm76tKjuG23WnRatgwUAwlMtQ5tVeQSh7ESWzysNpmye9VRKuGbFRkrl3MGRMAXv2khASpC
h5ja4oKlZADXW249VkfoAuvX3XMFC4i2/6UvWOLt+Kou9aQ7/FjL2iYQNThOYp+XFQ4Lx44YXggR
wYuu7WZ+jCihebDK+oMoJ56qnmnIfwyBfGUuk1NL8N3W56quT6B7a5CLLS3/lNFYbeBeCVqKV07H
Aw85Gg08Ck7MTef0aOXGEum2Pw1UFgt7h83lgfXml9/oAgQ765/gsd7ilcqXM71juvFsfanC4mwI
Ux7xTR+k8cMOYBWMwx/b2Qc7KFWM0av39uLaiWUj3IxZ+UoAWj309ImqMdpjKNWKGBXsGFOaUSLz
+j2C7E8Es93aygFz8XZNnMlcHClHoRvUuVsDxuc5POxxT1Y/wO/NnT3vgL/ZbVRikuW+U6SJ+Uai
3Yzn+jh5FkDLzkE13J15t2nNGMWYYGXQPu8PjN79kR6eXpwQfealOBSysicVOTA1D9v7wwYMtN/H
itCfAl9Lkj3TkCZn5U8cndqlYmQkpy3bSwMZWJFgIDYy2QvEYbj/cKR9eRqM4ovLiY6qz1EvrHM+
AqSiKxeF6yWH65jZ0LsY3u+p+a6D6Ns++nsuNWIuqhss5UvjpVrPTURWWU7Pfe8AP8ZwD20+8NXI
TGtie/utdq1iaIhy34NyXsleLxjIl5YLizsYxJMfQQO7GiVpZcDPNmv8SZG+perDqEGFZNqT3ql5
YmDY1brXv76UOuf+Q893H3FFkWl3iYC8pp5VTCyIaB3mBHXLZynI4kblyOHNWfnJvUCjWrTiGsEX
U7ciR8TREAx+7yvm26Z56PchMynqEODcsy18hh1WnLFFsRqFuiT28Kwfs8whTAXS0+TadPvUFfdM
h3uG5ioahJegjNPxfES/HGayqqrXiDMM95FQUPRrk71q92/Yr47XwPrVZyMsfK+F12MeoRE6JnAI
hvZP66vgEJm1zZHdgEvq4cDoemSDw5OqLUJBmij2evhJmIczxVjwSshhME62Scn+pfe+G8kkLE2V
qTwEsgDUxd49jk68SFWQ579coLf1mrAQUXYWcuAEtWggeZIZM/BPu3cpZzckFHdO5TZyGo9/zXXI
cHRIKD1TsVfqcFBzgS1UDA47mfIPXt+ErF7Ci58hnRcyhiScc2QZ5W9IInfdMXWsQ82tEWm1w6no
Us2bt9tNvqSkrabJzs/6EpnCLB6MCd7ukFfvDMtQLnk6UNe0MBFD2g8uLfIM1VoA72Z95wEtFE3M
i3dW/jzuqzxns5+oGjxsBwxa3siam3s3Yfs1CtA/XkcuHDiahxqkjF2jlGoQ05zR3NtLlvWmqWrP
XqLtmSQ1FBJlgy58oRGbLvcC+SmYz+xHvXBwgwa8bE4rGDvyvL91huhZKqP6wSLX7fFrlN4Ku04V
BVqMSt/lMZP/J2tq4FfFdwuSTrHAQHOK3IZh1Q3mG4Mijs+dcgja7gRvwyiIqwrApY3l+JTz92vl
I4hbE5v8+aVfTNvYqtZ5IcOGv9tnoIvdilEYE6aWGOE5uN4dtn+8qQ8D6o8LwjeX1Gphl0sAJV21
Z7h8Ah6qz37ZZYmhQR/LMqNmoeWv92nn+UZ0LEnUPHO0KW/ae9QtxwGXELIqvh9EBlYTl6bS8KbN
MRkynyUX2YvrdJdvYN81T7maQZnt7rwXX0r6P6GyqJH4eb4LHiblCWjBopFh+yLcfAA4ZsCbnNW7
dGAqYfOFAD5fKlW/fflwtu72F6u6irHuZ7wAhYxtyaAFF+vL1G354k0kfoyezoSsLXwwJFXeIm+l
w7vDHLNNCRdw5huVXWTwmsVyiyb+Gr1xcDpEyGfbP7/GsP3PiF0eJOh+haDBX3evCj1Toef4Bdyj
b1MsM77Rx+vNmj0o35JqZCiGWAEu9yZBMiBXfAGVgi0vp9J64q0YucVWGBTf0eaMIOlHIJ5SORJ/
8ERGnJ9TSiXfleIPvrJb0eyseayxA93sfxIqR7Egm7k+1IwmYr4c1e6yRcMLekorcaShxrrp/6UN
HFSOQIaNCoeElF5m1zmHl0XLWM76C8M2K1Q109G0R5oYa3btovSJqg9+dOyKOcL28JFiaexsRVeL
8GCNs8aYunw6lrgfSkv0PDbcO3xKdTFKYj0Le8Wg9Y80Zfd3EKVvHmkFtkV+1ycgEZqvIHUweJ35
KHNJDz4RTbgEO/i3Bt4y+5m6FB2zsNwFjAW0W49/AwSW18/9fuIiVnXwwdnGDpe5djV4LrUqYueq
xF14LefIVeBKSzcb1zOKrdur4YYvuvplyVMSCTLb7ffkYc60ntaFAKFCcUdvuFCj1ZYaEKRJI5NJ
vPYX8yHuwsy0LLg7OcleRXfstaPinBcV8y8H4vRGltMnIBvD3fvdw0uahErZaj3wO4NVaKwiVH8Q
bzv99kc/vauJF8hKzid+r48upwOG2JvGnAOp4S1YPmfwB/55mtQWj4lZjnQsr52bj6OKQk7SuXQU
UBxCc1md/wiUeSxbyt+tJbwJ/Xt78w8Mj859Ksl1IJtv1eQEJggmbrhRxN9qurz2x4sqbZUP/SdP
6HiT1OoyuAlkYlTOt9P4wibrZNo1YJsAEyyu/F2E9jZsYrVJPEIs2OoqfrOUCSfAowf8BMFf6bx/
3tnXJON6hFVwMnIHCknH2eIydY1Ip/mHVy3zUlkgOv8e36bWei7h5tbKkQYUS6TYlv/NbwQLV1U3
g/UMK5XxB2OjBW3ePy2f6CUQpuJADZwWL8gKdtkhUJ3x3zcjX74iJf82o1lmu9Yih6MSHf4Tt1uW
sAaKaSVAHfYpElQwF52R/k87SKS3+ufyjjc4gcNnwpl3as5jeUU4CQVlDOOWyay/6DSEDDLr3YMF
VposapHLg2bhXE9mzdj10xRsyhmaV73Y07uTYfVzD/57edychZe5n5KdKaW8HdelRf9xtytXzURY
mWUtsm8MIWz0IMef/uQHLfqI0yXUzASY6fQAiFi9RvhhQT1fVRwGvW8DdyjtiTD3bxpwLdChgtoM
w5d1U1YCN7LLfmJUl7xFketajFC+ZZwQHmxA9TS92XFi7lyRVB1o0pPQdQ1bGL2GsJJSHMbcnjaP
FBPnh1bFKG6jNd9coYIpVx2SaFxZuvXFJLNMz3nRWUn3hSgoDogflhk318iNJJa35bDl0KTKStWX
79lAvaCF/CrmCnh3f0M1ExlNDRTT01zeZELn5D00rMraRu9haN2OAuG/KSZmhm+4scM+8a0mCmLc
ZF6QWy4atHYlw6wNiVnvRZFzXErwcjblcKLpHU3BB7pgXnQRTfHawh12TuyEBU/W7mEgKTQJhnbM
wxSR4KGpGAtm5vZQOVKtZsoRNV7/ekWROdFTRL8vU5ESE/tP0OHVlN4ApG4XciMqkBh6JK/cSvY0
GNbDlWmQ72A6QPcXZAmx+O8C0RgIsxelYlbE7lS4v4Wreovtscy/2uA9Y7BhSIQAigpLfKBZ3j4k
ldvVqzZl0G6N6HRri3vqhvd1/bX1+mBXWFGNaDPtGxLkaaTPRqsybHiL2EaGOhlx6TDEkCXo4H8Q
8H/ILSMCwjReD2f4+5HPBWJ7IRbVcwwIVpqJdiGZeGPTBFyYtSqpeIG4ZE4YO7iUYBO7uXDYKGNZ
MYwMQOpoONBVoIrRUHb2zj8aKDMGy1qCen4hPQC0MOdu9OZMCu11ne+4sAomvToXBJipzb56UZtI
edDlJHYtPaPLdv+xc2lRrIAwpvSEJMNGcdcYoOfCk8SV9ePwb2ImtpIcRsmDOLOZmFfDsUsocTac
OVDBm3yhxKpToJaWFu0Q6VSZ6N4PHLxODhzRQjIVcdLJGTtJJYha0E3ABGCYhJTHwEC4LRZyFJyk
1/cg1/LiV7vEWeMZo2cn7cfPIFNg20fq9LM3/u83wvWaz4UbnW53zhbxVm1jpUDxomf7KFI1hCUW
u9u55X7Z3F2paFyRnYkPPDXlYybj2Wn6r7t5AS/X78+xsFHvv2Mhsg1DfnGqPNHVPoj2wRMX9VhX
TMoy0aYFyJm/CROkUGxyNrHdTVqGaZZwXA7BMSHIdg+KybG1BreFQLot3u0240afWVMA3nDCTbXT
yst8Abg+u6d2COFYMlC4Zy3hpV7u8vSXNys99UnpLmb9e8O+bh73haAWZ+aeqGv9hGXz24yEoKvm
Vwv6hQ/a88eEkRvkwVeVX/KCSIdQmMnZ72+24FTgZu5sdxqE7b2DywPhq4myqZGoqv7e+DNCk76J
WcMpjOmR2Cn00Iqq1WH8xD9LO+QHQ3EfnREjP5Ca2wjQksVRt/vcq7Nn2p+ynRA/wAxQ24FXdxQ1
jD4WGL+W336pmIn+5iF8H8oSABPxt8ENOA/Cl07KxFPcibwKT4D6LtZmTZC2NYgQInVQyzxqPSgK
hee6/yCyv7Pxftpb34V/+zsgZ1Xo7fWCAZsRHq7kLzbBus53wIRwCI/pc4ZdoH+OBhPh/OdmXcvZ
3sHroIFLi+XHWdfqwzxEanxvN56XNUxZaEUBj/F+aXHke7cTAqLaA86VqlAFDYmM5d7AoAmNd3Cv
ZXDcRGfSiNuNvZF3JGQ+OHaBC6z+l0PacukfbukBmqwaan5io7SH1+p9GLbaByCj51XWS7MjdhZu
XAEa6y/cf1bZNmhWATNb6OlwU3f6v7KN9OKKp/fee1c1jPic04NnHDrTADVcfGFHHs1d5aWFjF1M
0+NjKdfByiOFFYvr6LyThkxP0rVSc1OcaU2ER6t/hYssfv7H8DTm6D5VAwhbJ58bnhl33iEEKDXD
USRQUEKUm8JToY7t7edPNKcbO3/cHMZCc+3QH7qYILfQjZXLCEivc3bNkrf7k1lU4mOaHIkQU7K7
9nxeXqDP2BZYCwGu5wor4E1LgA64kFiTrnKQ1YueSv0iCAzjOiyyLrjLEFOI1nQkyARV0zR95yk7
HVNMo++uSMboaYh1MKLqskoyeLn3ypplXbzYX6GUoxP4wlHj3YPDUxVnmSPM3s2Njwn1C1XlNGR9
x+Khewzh/M+32AgZeUYS4jjhlSVjwNNYOzz/rOo4zNLcH0dMh3xEr8cDgN9nN5EY10BuhemVAyjp
qdSnNi6OAw7m27B/Q93wumfD9J7/FPYnAG2y+Aft5Cn8Tr/PFPm1hZutMn8KLcvMKQ2brZyCT4aK
m81uQF78KmGHdVpFHnvl6m1DzK/qqzS9PiRAWwAT/yeuZWMf5G93gs7TIjCmAXh7gXGNUKaD9Q+i
fZOVAQAVTgUEFZc0CK0Ke+opr5j9Pc4bUpp9X19YPVHwqFmIAVNKHE2XR1gzDTMol+v3G8hVAucP
MCX2pMnGD2gMaxavFVIpImQwhpwxOu30kc93DAOgJR2jbbf1d5A36ksyzlT3LzqvAd8vnXRAS4o9
V2Mm5ozZwPJHx13Zr60bjqFhY5TcTVN3LXIj5ys1bKu12Ag64rx+Cq5ML6kpOVvBcCvtiWQGPWup
pshzch7p6j8oRh+A+mdybwzX4xbwcknbNGfcPGSbjcsEUDS82or9sE8oM4EDZqwHT1oCurwLdGGg
0f/sIyU87HSXT+CFjxUfuixDr2hZHHjfmPGJoy7QZykFYWVkriyJaO0pZxs43O4AFSYu0Wy+iHkC
oEWn8T2F1F4rNLZyyfjhd7x7I5mPK+ORhPqtkbMqOZygYvDganfJFM/fLwcaHB8CpAXGN6uUYvVL
AwCSRx8zBRzRyMf/ZqZexMtep4QCdSAhptnPKh7AaDddxxK1FgbbXo4okxXhAr4SYm0LsGTEO15W
sl6VQZwqlYBx7DHAzEv6SZa3sBXEU3+4Itl7gQ0VnYxExyB0yQQl0n4lRFUQwSUgdignS2o9c/+j
vkKdoGdyjHY+NWgXhbOr1kzFMmdA8xK2OU13ZA4199nvXzzO5wEq59RuhqlF/5pANWYT0mOu0ul8
rz58NFjaje7Xss/sw7KSyC6hPzZ73jYsBK/QgaAg1eldW53uU5G9CmMnUx8wpSQ0+8ZI01nLfaAp
sp6VfYKO3uXSEQBahxiuly+fuVYVtMl1pn5j9s48dc4s0pBaa+pcZQVVtpEZKmVDVGEsTKkwAbrN
qsIPRYWnIm589d9wH0KQ2IqnWFGLZBwGe7YiKwcR4JtwfxrizwOOPB2ka1YwFG1CIddb8rwrpM8T
6DHMW5BiXF+s2tRXguben/oUd9dECirl4VNERNXfgOQOVmAbme1A8Ut929eAb02YWAOScJ22UPcQ
iPKd2XXzHlKSq7eS3DrwZ34C7PNAYDCUVL1xb/Qvwp85QUvEGwY3Fjsqsu7SziTUC90dhQ4pdbcH
y7yY3BT5rAZA+DFOqsDmw/1fTSho5cNBXObF1z0Rx+8bF1X3V90klsQWjnCXc5+xTVNSBzXOWXiR
8jEsz0lO4z3n30U7K2kEag1kJbLxHtb9wQ2f9AU83xdXjLZiSqSNpMiUgY09PZQOE0DLb/08Jsfk
SDyox/rntXa1xbfwDCgdaWyJk/Vs3P3j/BuWrKApB5T7E8YGKsiTwpo5WyytsSzOX1YkupLil2Sj
MqD7/Kcufjs9DLZ2AT3BzjR/1XdMhzww9O6Jmvcv/+2ajRFYibodyAfg4Ce1shDHW59ctCO7qYWc
ebeJzQV9cl0u+NUt9KcSivd3tzPJM75xwDxXjSv6gT9E+5+Ej2jl3afxlJkK8dDpHwLX1mkN18AC
0HgKkYjQVmAwVeROv3c/jNF8udp8KQICnQFC4QQF9PUw4HG3MHtxQEJ91RAYXknlS3FKvoUqJoMh
0oALqx4Kt4BvzeAMmPlUlMd2A7k63EC80o9gH6apng5oR8Bs9AgFHAFzdT2/iLzmqjpFMujd4gWD
Oq9a9VhZmKle5Jsy5Rcs9gE1qv7BMpnvAnpBKzZIK32qLHHsNGaw87GB65hHEMBAKxyrkB/mVVMm
eqEFy8fcH/HDx7UxAE0EONM5hiKe3MpHIPJWOSeLIWFnecjPXrQBVwSkbg1horDzJ7Ieff2UlWUR
m6F0zwcr86zTRrxTkqCk7lijuMUUF64voxqUkYSqPw+WFOKVPI9gvXEdwLhAqflhsZD2rqKqK3lo
tAesqd5NqsDBl5rmKW23/wMyyMJR/+tDO/SWWOnKD2K6ql2HuHB4lvKgmGbqbRs6lrpZdJ0O8Jd2
BN9S2HGz4sFKdkMMd19vQFgsDhufZnVGFeL/sYUnyFfm7g8Nh+HWszXO0ELbsj8gwUeMwnlwRUv4
K311UUEE8gaTXuBCgNv2fdDPT6UfFa2MgTz62WNv6JDu+AlFeWPNOIqPqp6TP7PoKbHB+Hyb8gsi
TmPEPoWuZp+ebqiCDDLEChMtoZbMwmcqMyP8M8M759x4YuMfNqE8zl5iuXy/8N8OYC6rqKBK4F75
+3Tepkuq/fZDaAtcvED/HH/bjhHbyCT9NB2GEMdgffaHBwGS3cXcNpRodCF+rXk3HXNk/v3sfmEE
Ax+PnaRwE8K1yUTMBlpp1BIkqPZnmZQ2wzP3L6pSmc19BjfWAfDt3SL004ofwR9XzMWEdGYIVRh7
Jf+U/dZw1Wz4s/i0t9ZQ6hCAERTxeHE4CMhY66QCjWbfQyn4bVzVyvwcgPakyajNM0GnKROps5Gn
HAGWFouytYxOVQ4c3PIxy/6kVLUg6k1vJRw9TNpO/qJoVavL7yOuNEm7ImoDyALIrd/KbRZ6b3Gq
rBV1W8gx/n3+vQRHWv7GtPZ8VHvaYjJwn53Q31n10bX1wAnzEyoy9YDGW5WLca6IIqMWrA357XII
i7a+hqht8TBQFHo/+qiBJ+ED101So4kSqdyllVVh/2Hut3gdHIurtXmWiZnXZnl0hErzKrtNOeLS
FKVh+u0ZvNcZ66L6NP2IPbeVg9X9fGAHAkl/JLQgJCDQ8vKxO7unCsMzBVn5NWGt7t1EcbY4u2Nm
/nyClIMCKsymdowktLHUeDMi+beUVoi7WcXul3HNUqlbUlgQtMKXS2CQ6VWSe3G72xP4cr+dU9BF
bHPWyMMdi5Dq+Qz1P5xXV4ycdNhKclPVnZu7TMMGsamATC3rkq+7syHi8MsV3iLEFHbL4zrTP5hg
TD2zcvrR8T1HX4at9se9GXpFqtPokXqhiwsop7KyJftWCxAR5fntUuOHQxyqA3zT0JSWt2Gv5OvW
wU4otYk2RbOesXOk+LEBaiCpi53wH6wkeyLlzORG5HaFX9SeAE3tKP1a4e+pcelRiUaTj3hvI1Ij
cNHDTZ6t9ZsBSvqLJdVd899JOrq41N0QljrNePiVzWjQkCiOJC4jvKfbalq8h1zXmClKq6wfb+ow
c5G1K0dhkE8HX+gNcFqCzNl7jWy4BdNhjZO0fSq4l2w5xjt8ObcTRYANR84f6HK90t9evzmaXR43
8TIhyIjrkiBv26CkVGCchSGM0VcSlYBP0mHHz1GaMqutgmur04KqClOIutAbpIUqhq3zVoE8WCnY
WZJvFQ7M8CjAYuMk5d53ts2ZfAyotPt4lRYxmp/gJegQvljnPHzJbqP6FjiumctNiSvplxnv+LuX
22d0xPZ36feX/InamxwqD+Irx4TwnUwxl0KClexCBIrFrR0t8Fsru7JPMqsSqk4Rk+cRhmw5YtKl
I2CaJf+PJKHYAdoaabdPrygui3005j3MIv8U2fUK4tr4uyhdBjEX4tdNmt8OmV0yhLwG6hKqfaAJ
3uDuHDc5SP4FN82wZfDxGGA7MQvkFDmfhlYs0boysBruANaByGoG5gTM1QqNOHcWKciBsWVdQK6T
IV4d5SLLpgLMY72mUUA7/B2MTkgPujq0uYfyW+63pbe8uL2BusKAX8H09xLu74RUh3UiXNXP/lUw
hfJYg21hyc2UZ7kLbZlHrqHkmULg8JFjHJuYy08ZY+yop1x5ZdEiCP6dAXa7zjvdsb4XIlLzSkZB
Bfu43ezGjcjpNwrYdovscg9uboewtsHMJCF7dkHO1te3dNUalUF0rJBkhb7hzkLvoJWMZk4Wd/s+
QteKoK8gpPu8/FltB4e0Beo4l14VnY0/5abLYPkIBXcv+h6HTQHUaOZZExFfdgbt2H/G1Kln+Tnx
5J8dqf8vID6qkeqkJ7Wb/ixxeCy7JGodfdoy2ToFBw/D/d7gYYgJU6ZiE4DfDDQKcNjWl6UcUJ2s
Cs2sSGw59Ws/atrQ91JdG5uOStFHd3VlTiIS3HmqdnCMZu+Dbr1XTDmua9pFlYIDyMu9ofvshjNK
Xk7u77IHq+HqApBDXNZePpw3OYgv/c6297IJo09H6D28VrGKUIqsNq1AsPJ5e+95lD3Te3H1lnOo
zdzXWF0wjelKYkObReHkLMMm8zrY5/+0evrDtW9UAdyEKwa+ihJIjK12pFb9kCaM6web0UgdOSiW
Qlx4N1ajURDbpJdg4s1n9emYRj2lVTGm4QQ2VlTuxsoz9J7GA+mdnrzfHDGPwEFSHQaSenHKefX9
K1vIp05buOXiFfK1iYAZpdqSNXMSYyxBY2Xd3ANGfoHwCSqhtyp01x7oxwYN7uMyLc1mCAcsNS/0
BlqVtT9GkGUBOMyMwRhVMhrv/WQaldLDeCWUBU2WlbWeURVXDCMhayGnBqp5BjDxhQQs1UAMOTC9
CfZApwpEPjO3494ehNb7gD+3LFsE0aPJ9HmtN85cP+6zuv1IT1osi1KAW4HZIwTYYEr5sItXZODn
aBeJ8D5UG9zX9+cfn6x5n1dU6Gpr29IZ4QxgbuN5jDPsreXJ4JbXM75rACKYTzwOJM7G2z+KMsG0
ON7lf6v7ujgeUhQjVv8e51ORlbqtWKgbC4FJKVHUY26nEYWm7t1S85gCYM/njxtyQ3PD5D8GqGze
F43HpOeWJ0DKgTWw8yurCs78GztOp+pW8dgEQAKES0nJGglXPtD4tDEqctr/xttNczBkNHCEB4bU
Ty/XR9U6cw0KoJRSmxiLJxBfz+ShIqfhWlRxkd+R1bTTEkDUEc+iqt3u/1CxZDCseH1X/H+hFJoL
FOZreUXb8NipI4QA++KnD3slgnU9avo6ODv1UmMkIVW/xGOLzVQisIJHSBZcSGrxNTnpZLra176d
KMEdrbgxm1TUTtS3l2vbJhuR7BLf2jMKBmvLmjyYfY24G6ccXRi49Ys3u2ZKE6C1/IZ2zD3C+5Fi
cYcQe/zid8H/SaIRJNAc7YZLzupJwYz+FNIITdqqPkTwNXlz0GB9iDiQvSYyg7HwXrb9jhkGOui9
N+7oSlEuLTzkPR9iG2jdQKTdB3QtcR+35rSafM8h9ObKDt1wadJBJSl1lcpHHDTONALxJnNImIBZ
v3WOvkzklhf2TwfAIruF3X5M/3RGXHBHBwIgFgzqIls4r7WRwkR7R+Ggj6mIIpDsX7U+wFHl5UZV
h/xLr4E+uJ8J4tATb5hsuJDS/3s6qFT1ZHTn/7emSMNO8Dn6umSDET9pzIhoIAlf4XDxSkn15t0v
CA4TzcfaTfeLakKiw1z3wjkzgSCA6QwT0eB25zMipiwPq3OhWySiqZvR0mPuW/FhwlsI/M3EfOru
Vcp7+4SrwM14xN+k8x6OQliiQp7uNaHKiEROJluKWsMnedZAx/5VDt1QKYJpOjlBWwnc+f9kk+w5
Vnyx4RRBCKuNtET4gSJ5zTNUILPCcnifE2hIkLyC7rH4lmtC/3GGRebEpgiZ3zvxHGMFSGAOUqb6
8d7swfOQvl0yfFbvf5V4Id1sx5knxmpOQeuItja0xlUvHtvbuoMBm7M1pZhLI8Pn5NxNEaqU/KhK
PUmxi8O8WQvd+4BFRjT32tqfcW8V3YeN5tmcdZ63UeTb6lSvyR66+GiS9Mbw4Y7Jd00MeobVe9xn
IokUkGJ1wREAbsP/nmsGHLJp7i1E77/qNsnekNJ6dRDwlJkWXqHwXJIlmnh8zUU70q3Z+4dN3ou4
OhoUEMkikMZSUQ3TTKXOFuCNAeqvXGeR09/01taQdYuPLyHFy35sGLSR3USFb6J4HwoTa1CFqDBA
FHNkIEDKUFgvzSLP7MKgPfGP3zwizAtaHKa22phZm8NGjXSKwBCb4fbavWSnObjDUWgYCFUP1grA
tJXatjylw83AlPdSuZpWJBD4U4cSZawcre2XNTsqnlpr8ViFUQza+CjPaHmz38Dh6GV7KQ9RhVdt
8NuMeSXAdLS+CuuCkdEiYZV9pIk28H1CpJzlJVJxHyTGTPcA0UCv4dStv5W8hWFJKTRrrjTbQe1Z
3dTEf/xfAw7CQAnpAr0P9yeCchScp/r5TWZgoYejw+wo7mXgehuEmays66ltsB0Rzq0CSY4UsX1j
muxSHujc/jfarLNX8AbfhafIxBJ78C/d5mwLnr/7LBgWxXMJdTa5QShq9y7pelOpFgbgsIbEFyyR
LEUhPXWcPHbPsRh6Gn9ei7vKsXAZjv+oKrJC1AJrDA0yC5/NC1c//Zs3u+/wSD1f+kUrUvEji267
jrr7IRJ3dPconqNIy9PDPmBIRKwlmc1XeBIskFY/QirKB18+E2AkzAnS4sEsYd6NjRizWljREXig
ucHt/HRIHNWWB+ljKK099f7/2UbPM4idiDVHB3ujsSYlLVFl6d4Tu87ZS1dpcJO82sMkcdRK/M5T
w9MZuyJolnzVGOrQjcI5HoXA0hS75058rz+vaWffuYfzAuw08mf8U2+TCyBPBrPHhqwPppjKnpSz
XtqiqMKXQ3ldQpEMS+9TG7dsN130JpbF4opiIFhvUQM4YFM5Cug2bljkeHpg3cde5OJVoOYGP47b
qPC7OiNGkSfns/JtPyHhxZ/MPjz8481DaaoRcQ7fRvFEFz/RIFGzjk/TSZtGBwvII9/my+/USNx+
BLOgnSEMDbAOcZHsHgyhR2QuFI9STMD6pSSw5pS6D4ZOO10TSJoyXZdJQZUa33Ss75/9DDwiaspX
FoV5ruOtt9QbUjbAI67x3+LhjKOVUXQf4uG0672NV/qXytzYrpzlgDSa5U4jZ3i2gPVp3XZcq39X
0Aq46Ty3RkafHyqCykSGS7F/o36c8+VR3UQxvz47DQKk40jKXGumDYfGGa7iK/TaIzirn4rXvEdl
henWFuLl2PcQ8ued2dUUfwrDxdnF4gDbNLkd8yGe0Tz3f1p/i/fEr4Q491S4kdK8ZLkXpxfFAFWt
tgC4H+uRfgn2582qxxzxGQHx/L4pfFSnm+MEr0+g4PMdzXhgo2Fb/kU6QLy/0UcmXwVfjH45iKjZ
EWz1eOuwAkQI1KeFiuK7awUHFFVe49Ht7w5jxk4EnHmGh6ZUQuIq9jI9GvFYvv/wKjxBbisISPSn
IIw40UrRnz9yYC/2ggqqHFGNkYVW3nBb9v1I2Zgj1R2igBhKLDFJeJAdniSBML/X5jowxPcl6nQO
ca1y89gkjR0Ja+LPQm/vw9h4pq/xxcLv2cr9b7WhXTJYiPl1GrwHPZ9s2cnUJ7HauNtPaWI+AYxE
IGbrNQm5tCn+wi7HOxGYPm+zGSeTS6pr1hZqz2vrt4mIhnujjG4S3bKklU1OPLUURsQZTCNYaU5K
ttGduoqQohcRj5z8rVq/VSKmfTj823oj7kWGzY18nKNQjt1VINhQnDIz8Rzs4fiQNKcmGcHdbi02
7ITbVvRrUSNLkL17xyUWbEKVncN3M54N5ZIzEXU5j7Ds6GwOSngVD2UGH0aar2zjuzNav+wlZEHQ
hc8MEHnfd2xGIR5r0YyhhOuQFCGALnr2I2LMvodNHdsPWLvJidyleNkeGsY2TCEO5QWnRtTGTxrr
PNoyJcUB9d9bD/QI5d6/VoQ6R6icZ6vEUpw2sHLiWK6Mb2rRw8yF32Q89uFV/rgytpKUDM1groRL
hnwXS02RK9mJjodVs1GpkA3roHpXTzAmpaZYM5hPH+1lAozsipa8OvpJ6AF1vBTnZQkrJCva4zzQ
ncAQsfUAXrDqqqYnRum0kEMTLWmbq54PQGU3AlqyV4XhEcOVsbJbd9fJd3JH1m2w0QvYfOfGS96w
62vgEVAIp4imVwgDnSgOjc3chD3zV2qHUjaKoEgd5W/JlPBoYL1PdSJXVcDK8SoBHL4ES8VTJt12
UWzSVVA2JzLiR0sIN1yXuzYMaHK543k4dngp4yT9AZ2AKbVK81Q2N/Gv3gqPDrczPcyjT5MTA0Qf
koiUQmLcz1abvOU91kbUJTs71FyqLAef5hYb9lyQ1irfuTH9si19h/1HSCUyV489it+ZCDXJuoUB
5CGdmtt/6mFg7Ws/eDFu9iQkEtKFz7wov8d3s2TsmH++9c18n+SpECGM7PFMpC4yCGK1n5P9Ki3Z
YuoOq4Vh6qlCvtBo3825zu0mP4rXiMDB72+RZJi5bUnYYcwZ7lC/+aSWzyMwl1Pl5l2zLAIDIiLC
I5JBnemCK+QHZI4LwAdNL+AA3V3aMk7wXZop8m9sRi0X9Vs+hgLshMHSy4NNo+hGkqwSYxmComdP
nGliMg7q+yGGMr2JBv9iZnHxYsDJt24qlsN4/YVftggMNkNcybPq7uPaCQD9fX5mLtJwZltXLsLY
yLsqfAQ0n2S8XHbctHXPrZVeJtx+ugnAk+vyBr3YB5dlyV02Mi4Rh0I3fW/A4ZsNF7ZLGQ4VsTTD
C463ucNhK2XD2csScefZVmVP7O6Dx2+qgSW5mCWMO1/1ASwZy8HMXN0m3/a5uvt75QIam6Q/2kAX
N0JVWPjh7hmDAA4VpJufGgu7fkFN/pt87gv0ilfYU2kuvfd05RYn77ZzV63qMP8NV5zwMymREdCo
Q5NSmJjpd08PkLPjEAKoY9m25gWdr8Jxn5Zr9jB5ml8HfK5qaMcki3yN1E4CFcwkC2HxvlDiVWLt
HyYIkiuw9TWXjQfKnPlSWS5WKlIqGcfTyjA4gIYxMhC3X6UuhLY2m7UHjkf+3hrbEep1MRoqresf
F5kD0optfZKZwFZs5t6geoAfMIZ1lsriv4Pc7Pi/hC4qFId24lW0dib9ou+MXHZ6ruyEOrt/bKx4
E+2NITyj7z/zjqSusZfCOeecMX4crhmqM5drz/O0SEIpTN4QgaVEhmVNs8KDQsZzAO600/fh7NU1
netVRJld9Im9B1eVzeDs0Fe6Xx1qbFKaunbvVevcDrV67t3vx5hP8RurtR492l5pE+RP/y59PIW2
VNmbe9JcEae+sO+0i9DJyjRrdAGVffBOlov9k30StCWEP7ItRQdLoD7RbRLct5gIy4/dtri85Uh9
++NA+YaGbveZ3tDqUkrFDhp7fSswYzwvORfiP9T7Qxj+0ome6MgnXe+HVeLrsEzMyr920Mtfh6ZP
VbCR2Jrj4KdTIEwtFXbiUtzxFGwSuz30EPZ4yQpfTjudycrih48Mo1sLS54fY8ozfMJ5qWMCd86b
PptDBKFxcNMbS8AY8YvYha9SPYUzh3LWz0Lwpn188Sce3/J7Ckyf3P3z8IIDJDkYYTSHnp/Aeiez
NaXcG/S19fzn1FK0o46LR3iNJcqn1/hKWO7CFyeYUui73EnDon8ZDIGi/VG7ZG8ukAUbo2FzmEmr
/b2B+HV9AW6MLC00Bacocb03ISG+9rMP+ahrW9YKRDyDQ3upmJmLgX7KoyEjXfUbiwLY4xCElnHW
tqCdkmiEQoZeEZ5cVeTjKlkPtsjtkKi99nSrsBktofp3zB2i5qNV5R4yefMfa87p+Hug2hshGuxb
k/G1ntLwe8BUdq0uTBuH9i9sqWV4HrbPHkMqsp759cAmOEZUTvSuV878t4wWPkDJtRlIgjNP3DhD
KXLoFLqU9qgWJH9Ykh/dMVhvc3iDEas1ntpmMuUOe0s1QBfajs9LUtLigZ06nrDnRB+SNsLQE17T
MRnDI2Aja2MYssMqG764CCF35ybQlAOvwIUvC0YO8Z+Kg6GoapknocaIjVdhsVGeM6l16bYh3T2+
c/W7Xm2DsJpAkltoRm0UnT73tn2L+5mIGOYbutIYwwv009QMJWq8McpJ3cZsF8BWFUkXbqFyNLbB
EVTBg+kNtGv1CXt6GsItMRcRWXjwxaQ6612gIq3xQobABJQY2ca38CF0bkl6nCMRcHh0rfjqB7MI
kPiMunSE0/ifo9gDi6c3UuKpFb34bXGM3Trx52/ZxpTCYPnQQkQz0Nt/g4UmMaJN+dsrWih9H7qO
IVECkcZbXV02lbkAH04dc2Bo+48usdGQPR0IoPe4A+MQTpr6J9Scjeg/xO/VIQ/qZFW+KShnFRSv
z1IKSTJc/OwdZzShwGJ1sIoHhqoxWRyfNpgfciWW8GVBJ2CDa7rO1dgsLnHFPdCSOQDjaNJoGnmE
xL2ZqHmkIPZTf9JYzx1OAqopMXbMP1onzefOS2iGNUXAMnPw/jH6ImWUaeewdtWMmSwIniPJKm7w
K0SWPDOriGiiQ2rGSxD5uj2iAKjRoHYG0CvI7Xkpx9Kje7xppotPiGwVOZhO0Kf6e0K+9/16j5K2
P0d+/qw/srxZfUipfcODLiFREA81W0cGNHcDo9LGysB2Vt8EhOmLg24izUumPeCybDaahxqP4F7t
1Ap8Dg/eggiMg27GWIJ98nX1TWiRaALLs3Bg5b9UbHEzCN7Ntlfr1biKL2valN0PfKNv5LCuNv6+
mLrCXct5PmnnP21KkZval6/x7M+MV7xjDEwU09S/xCcrZcNVpwcK0+EuGKhhMgz3sc7E/Vl6f7Sp
G/nFPai9RLsH9xUG3Rf3FumSKL32Xu1jiJH6y3jpf4KUkxwiPFGmll3rWZdAIeV0RK/vsb7RD4pX
7FU+HsqIhNHk5yfKpfD2DVIW+HyjSSnIqo+UOXcbEkvL34nqPO7Ux9xPY6fQ7E/wEMJF1Fm/lN9s
6lF6bTLDMPqpnGWlKEugtfcEnF0g0Ivzig90rcGbkmzDurXLAft6MyfoGpQZmu92k53ThCrQ+q1P
utjHGb5hQb2+sBHduDkdhGq4aZkjUj8kDudFkWheuto6Nlei7E8ySLuTn+9cJ2UvAku/pAmidI9q
tzOXQNTnmTbgcTJXVgQNbfYbLrWhFn5tCgpP8HIv3I9HY2dM9tS3ket0lupNnCZbD5QJuNGBBYrs
8ozjVo8e7ERhDjHF/juC4xXCy+ZllCfi7DpfNGk7uE2ow82v52MQDnS/G4iOoHH0WhaIbZhAC8kJ
gNs+/ZjaS6gWJgAHH7cgenpkGWmPDmpz0iGV19b5gsZ915NU4oJslWPcLrOFVPr1iMmW/IxRlINZ
LYfn/by42OV+yvveKsmiE+QEflqq7H3M25xj5rPOTEgSElsUZsS128S8W7pWAl6J6468Km0vgUpB
VyDaCI2rCaOIqIXW9CMv3NleerSlVetJxfzgvL5rg7Z1iAcNu13mFS+2m93f8WukKUF+GqhuY6ZU
AoQV4pPrgCOtyZuHFRMwvjEscnjTQzkI61YjIr+/DvUvAdEYsqi40CKCn3+bVXYD9x7v/vJ1jS13
wtCVQDbse0WIqtCxvRWf8sNmIouKA3YNr817CfboZdfywRfaJ1ViqEsxsytU4d7yuHE1WfHJ+m7w
rrwv4TibBWpFuRBQmnkJSiAsNTHWRsyeiCw0FNEtDSnNQ3VA5uoS7XNz1y7KyIsyn2XOcWcQSEXq
4sx10Tox2/kHC3UenD9J5QYeA0RwicADu2bcrPWgyJzYezoF8IS2TS/r6tY7Q9r0pMSWxe/f9A60
pm66pn/ofOaBTfGfWWMgKuZ2yEG+3hRHDbQjIthUnQx878Kzit6x+OJCj5QGZGq6nfH1wyq69TJl
epJ0qhL3NiRlXwuPDcMjCjquVfXkC7EczGzVoGBENO6uWfRbiWbSF7EeX0EREk70ktWUDDWDvZ9X
6kx5hNyr8PSAoRPnsKqJxCdDEbNGyo+NA1LV0BlnlxfxEFBRg2oydV9D9XyNec7LbWWU1LTthapJ
I/Tq8DwC88Ajhd+gJIbBkrr6LXhQRY/bM8Uhd/nqBWVVNOi1mZQmICtBpik0MKbb9SAWfkJkp+wx
6HYbi9Y3JQjKT2Uu553wbyQodCAE9RPu4w/zgiN6PTtolkflH09mpCXfl4EbzbieZ/OzbE4kxto9
3JGq4x4bZYnOP4NoiQQIF2eEdFdOAGs2vqIif1gjvLDMdirrAQrxyzmmn5mUiQC7EG9mR5Qmx9I9
qI5cYn/O3/eT7+vrSKVmxHFwEU76FryA4snbba7uxsNFR+GyHa32zIow0D/QLeOdUF43gZhnXFj7
j+iHhCx8CVNyhb+4S8qYOGJ0gpd1UoGPLt/o/i1daawTao+PRADRA5JCQCSgwsHIly544/7COyzR
UU77zpDJx3PmU1jLzlv1fhskSfO5F7Ff2/0SRFpQEO9jhCwBcmsvbP8ZQlYYBjAbVfc/TpeL+FZb
grH0tMKAdjoWCtPvmcbWWDPG6tEi+xbmZd0ASsBg8bOWe4alWYQ3YtYiefP0S26pKJFUCu18nGkx
3+3dBq6CvgN9nsoY9whBEle7UZ7zqLCZ97/caIq0rsMQHevnVhcqDJP2Yxt4IGtM68CZqWrFVuux
QeP8SA5wBX2w2/LYwJkscYE+m9pjuRNmZUZyhy3Gdiywv+AO8AL0eR3K6KXkVAFIKG0qjxcoPETo
qj2TRrZbpz2duzBcrBNXNDPp6lz2+H50zAZDsfsfgrxSZRHi93pC73topAKp2RSgIH7WZDB3V4+M
QcW+qJM1IwFLuQ4CBM0ELn5mOrstjazwR7ZuKM0g61p4GtuYIJ8dGFT9LYYeIxGJ6hcVvPlscTla
Al6uTaEMzuD5m6+HNIT8iIsiDhPWFRXUEm+ZdfBq5bL7+3nlPfNxoo4Wza7DkB8knXV8tJc+o87D
4b003OhFD9o1OnE1ha2gxFQ+St6HWtVdX1sl3DUqSDY3OEZ5nYU0pGmMGnKQxOcOAHK1a8REE7MQ
NnvNdD/u0q6EKi0Rm2ifnlXDQ9pT7+kssXLfAgbB0RPCQUrNFXLlpSfGZU2YbEMFW2eiY1eB0EOm
JinKncXIaLe6ng/Va6KF23PQMO8o3vQJvs83YWGSDRK1ABWqn6aOv7JQkc1PE0WZf7ANXkNl7ohO
vOcsNCHtMMzt1nZsQj5LdRWoAPDCaVWfraahusyyUZ3mPBQehIo8u5gwUPJwRn1zq1lnabZYWIdl
k+0LiI2BT0prIbwryZrgOf7zy2kBJh6pACo5oLkZ1YlSB4tCf4qUVAzvWNIwZpcWZH6XflvIY7q0
FCQxHsXQRJj8IY2s90PvD1WIsiWnNlKR4wgFWmmFzu/UJz4bT+1VJvDgSui8cSu9Y1RsvFRxAEMV
dvlFTeexOc9Z24XwkYtAKZbTl/9vp/ShFk87Fgxmah/YxBxOiBe5bd45s5dcDlEwtZaVBND/cxwv
9xgDVhV5BL2w9rBJktZLt1Kdywbdjxd0Sy+JBJYo4QMc+yPmpvGBU1S9cI0h4e+Df8XgTX9NXav9
B/LAyT1Mb1X56s/imMIVrt8+SNzdfdoByrsku85aD5dR6ZBdjK6bgme91FPXPv7whOAC92Ctj6YW
v2KqW5WtMdGgb/a4wbiQviyZSVDpOLkyQSwFzvz/DpRfoi6DQNgpKRoTPMOPYkoUww6CE08xRsXE
FfN+pdmqaia0k3+41gUJI2UP/6bPgh0XGuV2bcjEIRqWdFUzHb7s1F0NcyfLCBv9duND4vPUfL2P
lcqIHd8mtFOv4q2ShNdzVpXnT28s3znyn7mJV0B4aq4jRTMJAQYkkBdSKaKTRLSbabxM8ExMjP3q
CyfhZmfnLxDNKqoT0IMpB3xGvlLYuMz7cZ3KsvasQ6wOKNPNjnUQDfwYOv6PfR1Y705LiblB/Gmb
bvrgqtco0exw+Lf+NJkJOEi+uYS7AI2O2Daus6O6ZDIOQcQ8Th34/5CCFpWSpqMp0qCG7n9uGpk7
WdXraD1UCsnmn56ydnAo//Luqf2hWZOXI6lRFaiLrXow2anpSsVg5cRxk9HiEk9mkdKDUORRFiSO
o3vfvDKz7uf+4eIDzpD+fI6qGAwcEdQS8dC06bF4kGiEl9AEfgJomng4Y0Rz32L+RY+xQEBggOGd
a/OvTJLaEC5bGnoJxlH3fdseMYiJRq8q/0ZmJJooFIEdhJcV4kGl3kCcBv/DQlB+9YgALdfhOu4n
5iP9W29Nwi07kTb06xOD8XRw8v0XeO7IlGHS1kQ1MwuvY1Yrrekzpd9789O0ng160hPRZLv0RJY6
ngrSCslBGyYzLm8x8AVUOGBBoOm+dWLs0ma+vzUOW9yWgpWsfCIcZHbNRr7iEL/7bx+EM2/SeDPf
iUprLxO1Max6IglqbjPKUl898zsVG6mXmiO25CMLUlEYlCfDs0Kggo+Drrub5FBt1Cp3UrBPo1GM
TvR64dU6FxGAgogaX8YiD+Yi6w6KLIHylPdIv2O/6r/OqAON0Xyxi77zWgIYzFjXfQeoI3LQot1Z
CauDlx6/HgSG+eTraYoHg7X7fWDyQIiXdRMc/qwhiplB4vb9HYBqyfMiApfJQtstO7/kVsyH8RHA
dz7F6C7pa6tI9z1L0QJNlIh9lUkxtnvasqjw56okxnPPeEbssR2TzCsFegWIYTeMjaSK1Q6EA0nz
LYVl0wZjHpnqmhSlBUt4OmGQXYBh0qOMup7Ge53QzO1aWjyJf+7x4vebjNXGDBCWq+wPDrc45hDr
9yBD2ch+Nuk+VYG6MEuIfPWRShuuMwWIF93L0opEtlqDQl/4BhsQGYYhTvd4U5e4YoA9sYzQWlgl
/3plhcetiv5q4C34AKEl+MjN3KFK8AQjWdprfL1khMAwwvykORxrHm10ro4HTI7zMKVDHkz3y3fF
gyVFRuFuX4MWyifgzIGvMrtU/dnApThOl/uNZi1s/kJXV8LbB17k1kf16t7CUvw8Ujy4OADVhAcA
zouCuzUPj3RHDTUTUU0Cc9CoX1q3kXm6vdQapBREq+GjtsMHfM0jVZ8WzmN94aIhr6EryNGMlEW0
0nbM28bU2MpuwjCmmGKp8zrzUCh9IufCjfcQMfP/rnGaTAUTktLY4CInT2F7pDZgfag/MPpB6e1Y
qJeZnxBqq/B8CI4B0rpJR+mvbZ8rKmRUO4jFWqPZbkSlTz3kz7m3LclH51PtGis8A98jUxRGooqn
NZJGC+417Vf2P5Qacwo8v7XuKzdT5scX8TimiA11tY87eJvYon1cHsSMRncWcuttULkraDh9b9MH
PMDzCHqGuM4e+7SPVBk9PS2HbFpf5X2/eQvKz8vPoXOV9W9Uc7DL04Et7TaKt17Hsy2oTyQCdMfR
izeqng4CxrxXD00yQ73a37NIyd8mguQGMw5L6u49lD1YZat0kqhmEeKtknFpuEZcK6U459wXy11J
xCoAsOszo3/s7lbA+94lmXKCqYWm1dMmdUg3//JJUMLXzetoWM/KVsvkgpComcw12uA+Gdcw6yp/
B5lC8QqVDhyMus/GuScinD24eFGantOXQe5cXSUN8rHqVnr7oW6BYnSfY87l/bx/ZT3fYu/7ocLj
VdEYhrO+doBLJQr+Eq7h+a3I0Jcb5jQEhSDBhnZc/lAyOih2N7Uen3GTOF8FmeVCv5yF3gFNOc00
3lg9hdpSooVbMUz7fYalCHtDkvMS7SWTe2KAIJZRQPq035VP92lFQC9VNWn5Vx7uIgU5ojNQZAti
3W5Qqb2TPzQeIgYEDNOu09Hn4o9IJmlaWea4OXdetN0dkirT0xpLkCrqj69wXqzj2gwWhwXLHj61
/zfJ9jjBEMXjyS/mBdyycSwMnyGYHBxsREtap+TqJhtKCgdcrXdIrb28ARaOCGkDngvDlGraCuKO
UHr3ODmjkIehveVQibG3NPJpC8L7JJlDRhTec2RAa706VpSZTKjNQGnCT1ckeHQwbeK3Mgwcr3Dj
LpeZ+cVZgI0eCILPYwBRNb6ki3UkZrHEGn33SPS56LHoQQkUzS1rxS1HwFdcagREqULIR8zWSXhA
VSDzsSufTkPBNhGbGlitscgP+8NNhJWvIbPzJQt+2ctFNMHFlk7BEtqPiSzxETflGHJm5R+XFlhl
XNPootbBumdqs1pHMbjo30Ciueyx+2EpsKfBSypn/2HMLvFuBT6B95hn/wdhbNoVQp3j96JwO6HR
zViWcu71j2KkqN+V8Wkd8AMfNCxCNgWjydrjSWmm1lJnodTI003LDb468Dbl4lZukOxN4uRxXSHU
NtySNR+IpLwADzA1c5c7BwTZBQZ1r+1VgDcbout2Z+LL9ZT2s2DzJylvTx9oJY7Q6BpwShhqjYOZ
MLOWbvxEvt7+WB+w4ofpMLscTZISwu/mukqsnUUyXEn5fOsjL3FevXx538HfrwJM7wQkzLPtWtve
Va9U2N0U+6x9hIa1oA5xpeeuKYBu4GEnYl7xBBX4W/kr0C/qGIs8VRYdkUjWaoYgELuuAfRzlB8S
EhUMplUhskD2qKVM99FFt8jFqTJdRuNArzrdJEuUx/e+peBfLvMA4y+oHXIpniW6RTH+Wo5FJ+Ny
dAA+3PGTom3SQlwrrHB7xixliuKaS5A8Kyp80AHdJmbSjphK3VftIH9qBfKWqXKKoWpOfTgJrP4i
d/l/CBHde+xVgInuz74leJF37YWc4WIv04HcYlNK9DaEiKn9gc+Cmc6P8JdGfycpId+3L+p5gA2/
YWcTSOiERc4vrAkpoFULNWDAsyCRLiiEKMJdKnsNzC1wAi/JlbnFe854thtAychM6kGjWvbBAYtl
9jn0todmc5g6rUw1dhPlGAlVIGVstxOeOQOZwgeGZiPL4U0ho2EyTUyVcDoFfPOqrh5zMViukSXo
1ApDl12SmkpR09Vgsor6sF2Zy7hXz2Cb07hhHaJUjPgAuIsYe8msDITUqw61/n5MOrH5KXNDS01+
TVGD0CQlG9x5q6zoFkXB91KhHjISsV3AmsShB41qqQeO9iqjlaVx9gRfRjPXeIulGFfRm37FDNXI
Rh6NAkbSqU83vAIy0kgat8o4hZ/Tv2w8NtXL6sH1ldlQQQ61gwkq9lrStD5Xbj6OKosk8De6KJ1P
4BZhQojwV/gyhRBz37VuFdzIhVi5IS5JD9RFNqZSM3L8MltRzElrv2fxu5AylMiLZJK47AtAGYHf
JHf1MnWVme/6/xSwzldW8Gl7eI7jut8Vwv9SSCDt8srbmsUbXRbc9Z9ijYHStA+UG1keQeyQsYZM
LQckDvC1O7MS2no0/ZnLVgmIOmSJBqyHyY9xQksT60RbQssmOC2MMXumoj0VJaxRY63xccnmuAnD
oU2J5iMHCPWNbfhKBbfCQwXTrdOU0bq/b22ijFMNiBPNcL7hzaDa3gRlF2izZfd/T4oexYMdY0YL
EO3PMsa67xqQaU92QQ/JSFB8Y3E2ke8cPjTG6T91h5MPE7YtRyvgcE1iiYmonQy6iZ209gPAjWLd
+7OpRAf22bD3lKfOM9n3qaKeNRBlCt7wUHvsOd96Xl5owgA55U0FYHDRSqi+NT8BM7eRDNNNve38
51ymZkAq4+ZtRMCUGULkugmRKG5iaZ8rMRE5yxXr2JisP2pbcgroeSxLZhsUaBs8geYmHfeftgU4
V0R5KDcEzZtRJGhghe1rP2LJaUGFd2vEUjCOlHiHiSZDkctydOU4ixUVomST39/54X8FT4o3yqft
eGG7rjKqkMP4cc5q04JIyZW+wEmrWxWqf+2Uqy1KA/LyzehMaRVVCruJNU5o5AeO+9acW2G4v4//
f2Rr7zWwEFnR/FX9/Dktel8TZS5KQNczx+i70jWXHCS9WvtHz7ZbBqXXI0Td8ahr/Dg9t7mBTHZK
Q5pRhKTABv6RANtgn5B6y3hsmV4kWMOWyF64j2w2+7tIxb3eRf6XHK6d9iCtDIaqP64rBIVSS425
7/3O/HwRHqeaeRaq9qqCjY/lGE6fuV/tBUw42YcTi6pKrxlSI3ii7auPfB8RXK7cgVvUsCHWapy0
JUUM+BpYqdW/B8PnoT0hyibJ0FxFmPKODxMQEzU8BhbAQXYNfrBw+6W4Oh0SwXh/ktBVLYSF2Fv7
wU1KMtfdAXvp6rN5Gp21qolmN86c6nskQsWM+OOAU+uGMxCIlw/PGM2Zocm5V1usdNAcn5qxvVqa
A2qeafnqwDiaae71WKYntp1G5YpgN+QgIyQItUZrxqRWMJkYy7d0M0tTnhJYbRFi6vo9MWA0d7uT
M8mVs74/kjC2MyQUjDBxLRS52AmUwTv4O9OEX0ZTK+8lXgszQgiyhiiWyXmjzT7dSCQLwJLpaFH0
spVHOIkw5yFk3p+cf2cYAaHZEzYZ/gT4ddZEDbjNfKRXeDEty5H6CMASaPyc9EI7FU0CFCSZDkFj
0/+OUgVje82w+6dxoj+I7bcGSprLTCO3F2dxZrg7PaowkrrgudBFWDgvwd6DsgZAcgPDpNjlJIzo
xWBrFEMGcjSej2qRoE+OtF9ofR5eDKr2H0LcCYmEgN3okjWyMbvpfIcsntdieV/WT+4AwVJgN91C
5Cji0XEd07TtMpRYKyDGaqiUVMh/TWmveJZW0w/xU54gm+b2tXw9XBpk0uDHZgYfEjesLwCD5LS7
OMpwMfVXJU4ai5zkIYWQKZ9D87X9nqp4vWfDRrTC6/holrQB9FOIMfvV1ffdykEAIsWZp1o2QThm
qsYA5mrOUgpSzqGGPlgUj4HKvpxbIz7XBPsamq1nDAtdgaCqlXXt3Bz8ZJPeK9+7K7CFFWm/10IY
v7CGgx5INpIwOY9ArGRWui3lRn8lABineVJdJ00Q2+j61bMsjUozs4parj5hMUyyaYU5Tbgj+4P9
HN38km73f4jq0SVYW0WDxb7rT7OIwHWDzyZDtmuC2dj8WdxYATEk3Hz54hcrtemNcsZckfF9dfpB
+jAqepCZBWDnvlYj1/TkEUibk9ySS4+ITdAQ0LoucDEY6AW+TTYw+8kfc5rODGHX/xC+h0/o0KX0
tbHr/G3IFQa+/WK1X6nwS15XMWK4asvS/1P38HMdEUyeWzdQSd3hm3+Ih8RBmF8zoFFAds2Lhkuo
EvKudzDuj5GsenAClfd9QRjjdSC3xYg6agI4KJQ3lg8/SnVkMzJcaxNXrVVl57nfps8/nZ6D5WWl
NdBycw5dGxVnMmAvFOKFcyTjp4S/Y7ZopWrFa/BFcLcYprSNcq6G9LqaidGZDcKSVnG5k61ofKU6
IyO7qUISZ3TYlNuBc3UBP0t+hXP8SyzXuBcuI6IFlMLqNcVrvGwUTrlNpVq6LLiNNsuleZb9Mk7c
2gMSZU4vegXcjAOEelR8AwQDdUvFwJ5dLCkl9+MuO/xaUXEaLt7eBJLN0bf10IKv/PoOW4m7S1vv
cxNBHwR/pyIPgnBRGHbSqhwi6uykn4TCLx0toeJ2YpEzzQDA1blimdyIg4BJ6hY4fgwxZ5mJb8yQ
9rIsb16cOMKnQo0leHnrM9isHS8fJKoPyftELNYKDZLzIhqKnCWeqDydbDxeawb9/3BDeUbWaHU1
qmAVJe33iBafsM1SsYGOxXVZMrPwlqkhnO/Yq+x6MxPbo7xzp7eWCt7ETF6lr3Lv1Wuq1HV60pPs
2Cs8TRyGhEES6NkD3ukowh2920As8ccTUQ6eWzbVGqaAI3cDzK6gh66xasIDNGQOPisb5eN2aMwu
DJ9b55Y4w2KVN7uxI5Rn1LkBOYKtG2yIMpIXdCwqzXaFjKMch3/9tNEPAghiTeEdjPHHjimbsEgN
/9k9ERbwHIlQ3ZivwsQb5fOnNWH9vkD84vlkPQqkz8Z72S7Oy39eZNN+rdPELsi7f8pOI7eoWj/z
sA2W2EjLMzFnEpmbbVOjFt6W6jYN63RTwdACBspH/dcd54D06VRfTngCCDIeiDUL0sFZOB8suH6F
95+ivAUqi4P8bgO54UuI32m9m90bt5Aw4SmjPFhh0+Tqlns/o0wGejmW3c6celQ/HyjeONlyudyk
YHTVFj8KjsbaYufogkHlcKj2EJng6O2RTQXlH3EQ1cfCqji8wiEieeCj9IYE+yL1zbAMQ9LDSWr6
ZXsf9EX0PsBMQU+SbJlP9CwoMP1uv2t+7fA4Ma4wQOhtw6T+6Nknod5TzaAYQXLctgNgjRj3csYc
ycDLk0aU6VOdj8vFFj2U4VVlTFUIytMjsDKND+a4X2ZnAtFlAMRkyX8KUEqfVUXpsidj5HqmW3eh
lMXZTAY3cD6XjgqYba8uY7My13RwXOdyxUZOZPZoHUoE6VklpmP9mJd1ZdtV7wapZzYR0g2VAggR
uEYDR2X/lHRrOg84DVDR0IGdsyaLnmN7PDDl0/Ua/zfIS4Hc1NHwNBL4Hv+5rI3dcCGPiifYmkE1
UgXI+eCgxy5xQgbxno3YfYS4mdJnmyUQKPrrLPkERL4uAaR5DgoPSOI/uCtn48WORfycyRKCb6Ve
syYG0rh2gvh21bzAo4vohuX+Qnyc9OhAZw2HpxC5i/6+7DIrCdzJgadOqev2CC2YKtLLELdzMkFd
NfgtefLxrnoK+pk4WJB1NFC/M85DgFvZGWTFtERoc23ME/hcDQyDlDcDpXVhEFOLM9U0V9CYFQNi
FIPJ2OTxvhigMvMQjOQK9BjxNErv61ORyx1uBBvlXOef13V3Lf5+Pj5SilIprkOIAsq2Y3wwUhP7
BW2+vkKxWsjYkX7pMaN9FEjBYOCY7DgavIsCqfYsSdtvU1t+U5oMI28XgDUESsaIsKi4hwouu2uM
dD2i3vBMOw8Y8xAr56shTMI74M2NaKBbHH0K4AE3Uz9NOnNvyFikqmgWMcbU9RoBXDshIhh8GBeM
0yGSXiFV4ytJlO5afV3v6xxKvGJ+GuBojtPoFmkSeLSO5dfUtD1AgDNSlkiO0LmIZcVLzvFB60JU
Bq9WZv5GS91weButPRYchJ5IqYhN4CZwvnTILkDXtFNR76852igh/MaotFmWrZTiI1fur4ntaDw1
+LifzUu/VUpkwgHpjtGLUliLY032AL61V8KkuuKOwP9BqA5cfTvl0mUzKIMbR3uWP9nmtKu0zecD
Er8y04jBCsAppUfFwrai0X1BiDSxv+YatwiKOBpW3swMP4IXQoK9jAohm/H5byFDscE8UkhDKlUA
u0rOyIlVNqgAGtM0O45JWsSOPnrRFStHCmuTdj1V3yo4r0qrHM0+xAgAN7FNsAdAPyIdHwtDRsXK
ks2T/XR3XN96/RIv2dHeqbwxxL2wjuSI5U7JoRxO5EpqdHY5DGm5g5vcyfbpQObglpLxe+6AnNvw
s7Q4NmLnarf84RoNtNpy8dBFLJCa3F/pRgNZycrjKvkKeg+4sPUiGwQgP4CjhK9ZaN9cQuRVCcU/
k/c5d36r32N65aTBmoPZ2S60rSSvPcB5hOJov88JlRcG8n0siCsO4wcB1JbRuKkeMy7BR/pPgyEs
rhzIME1gLRT9GRxspa1UCVKrBMFIRfuBZg/Z+5dkfPFBbX1kwiFjVPqqDsInCf0BDUptoqek+UDQ
llyqtuxjb1m6AWbx0pl4fnQF793lmMEhPwyKRKYFqTe5IDtlmuGEySbEE4CIaHF1ElnPNszMWJc7
fA4Lge037rMzjGqX6kNA/TBp+GR9Z53n4vUQYXInte/HZdKRfrkE2Ht2gdsutiuOBCAaVDh8Lovk
7yKyd4yZe6u3mTe9AM1wQVHzEKvHTroPuyWnTGSFYYvHbvn7EvRZRbogqNeY7qxqRoN8vYbzjFa1
lII+o6Mft1IAEoccfRgM2MPI+mNquDVdk7/spV1O8RkIbVZHB15dHlYGhY3Rw0g54Q2a6nbFbH7o
4VEa5Meat2doo2htFukoVeF0AkS5SrFUDtmUJnDXOQzu1hwWvkdk3QyWPdBsB/+46CQsrUrOZuby
VzI7Gu7X/VVOwNhwZDZeiCG+3QF1R7qA22qnft6JkgAx+4OPLFrdLDyeMKjRrGYdSuXX6smimuwh
zrNFu7zXPOc1qGN560O/7LBt2mZrEWnxdgwfrJf0zwbStvc5JXrk9dLXA48DmXSYmIIrFWtKjxBi
JWcPP4wzrZye0zCbtWIrE58078YKRm56ZvP4ygRncdFEFIdQt0meR8ftE3Szk1JXJouMeEHmkgN/
7J2Q1p6eYSn5AtjNJANioo+Gxm4tHMYUzlK4NNHtmUhB4YLqV/vt6F/0JuzAfSJH7Qhxt8dSdjdV
deeOwiM4zP2cLuNQW0RqrLD+ARx6ANNd1Lq1qaQaqUNjW2GGCQoZJX+d14jUlXiHzC4Ix1d1jfPH
Od5PlPD2qsWqTZaTWrfYtC2/yEKkIqgOSCMBMm/6aRlyNPXiLeBZDUAQWUaNGwdys/yn0sN5deTv
lwJr/3pgAFVvNLB8rSk8WAzl5zK9k02YYCJqN1OynqfDuDdOppVbs9iApThD4/TdsH/iAcTskuEC
53mFs0PTtmshTQHOIf6IWZ2gowSnnwZQh5q+RcxpAFENbty4Oh0L5JTYcMaT3oqNUblPeysCD3B8
3k3aMI9MTUSKs3OmsnjlT6qdQZ/aI5yH56MClQ8VLYjAauRQJpgcCcEIPQKA2mdhHL4e4oJuz1fK
S0T93Kz5dN7VokOgqO5AZ2aI2hQR8MvN/Xnn6lTN+aaZL6T/wi5uLJCdvx6hG1l43hG2IBD6H56E
7S6z86Gj3LoInmX9Lc4AIjOmK1lHd2kNBG/LwJ0mUPWK42pR3rZPx63YKKVs2brdfc4+FXtdZblc
zWIzXXBpGG3afXl8VjtZtEM9q/avJtidfu0O/7umf0kkMjssgmw2pUlPMl1sv4eSAbTf5Agod57R
vyAfhTfOFruIz0DneZ5NmmIquOjvE9tVugRtbu8rhK7ZLKtJJQPOYvayqWBUtMRi5GsxjhZ6CxeO
IfnhBUFbYAQee+vmpAZIW2Wsnhi1EoJlxPh1ZXBawaFey1N+mm9XqCPo4w78cbxe3MrOUdhZT3nZ
c2XLUvpKC8fQP+a1H2xZY5PQhIA8jPAv0a7yHOSvVWDmwbrs/2ILeyQmiNAC0xEm3B9Nr2UoGeGp
H50ubmNSLJ85zmM0I2ue9Krmtp9rzWtAapeqseOFWEmMUcfRlxboxnDJVD4KQYMLljSh3VFfYHdC
4Yz7lIiUQ6NLGfhKT0NqnFSznE1isJWMqSHlOEu1dzb51yXEHEf59wtb4UfcHaBwk4sEbN4wnltV
ukdZOftgZ5GwfNhyif5gQgS+sfMnpSoXQVtVsikOHFLwnTTWapxixLxdR42p2zueITx3FotY3quM
XE9lRJMNhbpM2+dKc9YMNypE05ufTHr94wgtm8KycDbxo1iNQpP8tNxUcLuWZBWh4oZSNX6EVU5T
wgeRgx2VOGgjl6vFkcTygsILUd+xgv21YnvND4Ht8dPwkcWuSSt5dLo5XvUvHIxVi0jIeOyhnkyT
EypwlXJrDCBv/mdYvM6V0QyVCzCu6uNtVp3Z3Wt4vL/6KcP7WhqE6O4Ar2evR5nHZLtOayLx2Fcc
ZNxWFyOQZ3ptaqokyHoGk2p7ybCwsoKR6y90roWZ/pxlIfErMc1117LjVb6y8VqOY2hJf7M4qbr7
o4/DGivcjUQsVMmcx4QnppZE+GYvmplxRSUacW5InOKnmrEkv/B7ly65kYJ0PfUz88GXKLfmKRY6
HBWNZpiprxgYbzWJADygKsFqtdscXUtavMum5Fmc8MxN8B6YXAre9wPs886exFi9k17I6lvTiOh5
fb1kP0f/XIZ+CdiGaq/fnMBKSUUjA1vh60c/2gW3J3uaNUw3kSRK849W6Bic67wg1mkyqu4mcJiw
LtMW3shzucrsLMMPMIgdOR31KaqIenIJLe7jax6IHwG2zPaLTNJKpHamaX3h3QyQqqglj/VXWS6H
pw0+IkSrkSxp92uAmS8sP/2J7uVY/1HZnbWc2v4LdhrwPf5Ny0SUBPSnJ78oZ6j556x0SvS1CTZA
qlXgIZb/98XoUW0Y+d444lr7O01cO/eQ4PlPyg2GXJ77FQ96u5CvfxxMVz59GzoKuqRkvHeD6X77
m1frdaT8MZs5n68yBpA3E6aiFwt/BGHigsqEn0gSe6xrL5OI63Vbs4/K5N8oxgB6jR47Vkedkkka
WZ3N1mnyen39ibNvS6ZNLQmHFDkYFWb42bvKcivbA03gjqPJx1ns5v59w4eS4suE4H7I4qJF2GUy
u8bS0GMytJgI1q/ZjUCe0OI6Kyf/1es3ujOqqYDg6YmiqN3vlwdQn//tDxLhTPNOdjPwz1AJ8YEF
Gd/OaMqM7cNoqUl8c2/GV35wPpof7bcX+jkDRKU0sL52TGzAAZpI3metk27+NaFbVYZcxD/3RGST
4f5l0780dN4WwgoT989FiQGIVfASNMe5RkY0SfFIeFbRItknBvyShCAtlrg7dZlvF4AdIYrAV8Id
Ra731Db0ULACo+weEYNapgZDOQXQoed6Y4R0oGmm7Flolt9UAk4+SAMHIGUn/cwjS/xcMM9gjVLq
yOs6DwCJdr9EpFOgKf9hCcXC6ywJQCSy62esKZfNZFLxsOm7Y/x4KV9gEzn/u+BPkuvKxW4ISYQY
vDwjwzm6jeLv8FaeqhAiOsRJ1OPYZQ2vPZErSYi13KVV1IpnmmPiZ604JLZsMhxpw6qV77X455Ch
K1SfXOpDqe96YJOykAlbtqyWvbUg+aX2BlQK2hwvdoF3cPvq7Hf4LKzafaQsuZGK0wae81syoNTK
htlYyJpWBXf39QWI3WviZ4IVm2QIGU3xXi3G1htSFeBudCpappmO6rccmmyxML5JyIJ1fOhz0gWe
QsD9pcSi4kjRVe8/9f7B3NlNxDmJNvGF3gYZsT95auyKzYaC4m9V+ITHHTx+b0D2W91Lt/pSWy5Y
dBkwYpGPxgkZOhlqTpKZYDwCbK9mjqaGYRnEo+D9RyVat41ScbhvBPsnTrnwebEmiNlyWz/HmB5K
8E93RiClPlCl71dXJ+FplLRfKKg5H2TIi97lwvlMvZrs4WQS7k+7tpzf5OvvyCa+KXtq+IC6lCdm
rpPlwxIgFk8LKfBJ7pYYyHY+7VoDINwtUwiIJYI12ozmrqx8BJP/diuXN9WpsuRxuRpIfRhUXJqx
fuSSQ3Emgy5JPJ8daHdqJzECH05UNiXvrILkAHk2HiIJgNQ1gZ7jE0xDu5dTHmMx3wXm+Qnauecv
xh2jlA5jzqMoJt2A8t1ADOA4NS9MUI/GFxlxBLWivE1HPWkMKKvpVIWAmh2ZFZfdvLualyBpU0p1
kuoMFq0LUSQ8I+nOZwCeM4L1V8hHoK4zJThWQyP1Vpjt7QljqVhyVSfx/wSfOpRbUMMvwJM3NCov
l8Y4ClqWoYB+QMU/4XDO3qXGk/Q+NenJvP7hcA82gpV2BLUr3fLJXMuxTSER0E1oKIzfyrwQ6u84
Pjf0nKnAr5Kw3soGrt8OKoGsW9FmqtDTU9LdIFFDzv+vJKgAK+V4WE6W8hD9KXrLJaVrVFfICa2B
Ww2PlNACnhodHFzgtZekcw6h9V/hy/gX21bjbORKt0KCCz1O+x3RD1xcZODwd0kqS3yhNHIT95qO
P2U4lYFxEN7KsrNnk/PqYs7XkhNznYSCnGUdk1sHD+9ATP1e0IPDeqhJrlNwfc5g9nIDq7oZhU1z
OO3sLYQ/fq7IEwyfV3kouy2lMPPk70Oj5B+9BOoWHIWC5ePQLQh1VTp4eKc0EfSWbpMA2RIWV9uE
PiAwdgCYoH1hVRTnBk8Bu28/zODhVNT6tcZYG5DOzecjR24UnEordGq+tcAvOnpMdSrCRVTzRGoP
uuAHsANunw6JcB6ePawe4uSjTi/8x9sgYOJV3FFxgC1cN5ySjXtYLfkMdPIbMIEIdNNw+dhaUEtE
LFmDdfS/TMscH2fwSmgwc20aKiJricQ0uc5FKgLxKpEE7CGi/aoTyn4vniCYD7hjTlaNM6Ulm6dE
JW38Zhl3RvvWKkESlNYL/OkCwNYk5FomFKb5tnD9E/22iiCaDmNZjUBX1fOFnhXZjcCYRACTPJxe
gRPtW13loy+DIjYPaD5CCA/tDRSRbpixOxpVPK6/CRNdRTXz4/ui2hUc7MRRmU7Nx4ZE0tzjyCQD
1Vja0dvf7cdQu9PI4yLphgcOKKp0xTnsQE2B6iZNKp5FP0FXfDkxhs/D8ms7ixF5IfMtEgCG6sVP
HVc5q46ll78dASxe/O9dGuVQblXgAtMrxuF4OAqSe6jDIANLaG2aFZcTPBxvByQ/y16PDXAFsHgx
J18ztG+nUD38E87r4QZIcMGql4OmKj7munylXFTunwM45kA/lojooLU+afvhkkejugm9FT4yc6PP
TSncZOWB/zjYmJj/Ss/PzRb7BTjAY75tz6bsK6Dq0mjqWpdoaTy9VGcaz9Cg2EJNEJSFttV0RAD1
b2uXLoCBgPk2EjJ1BgDkp24xWxOqBf3NvodH+baJcXNyt5QeENM+WTe52t/eobInGiz/VBABwFqv
wsPO9A8J4Dfp7LlrLocP6ejlgcmRIlwNsFBSkM5UtRiGpr4pjvM9fdjqsIXLIJi0ghAiqRUr9Ruz
crtlNqbVEL6Lug5JyF+cwT/zoOFyOLHBaNet9RMvlKpRs+KEmcFjNyX7JZJ1XmETjmi+5P9QKuk3
Y+hg1cn20OooREu9D5oEI2cFu9lUEXkHAGHMA3o890Zz6U96Yez9ffDAXN3B75b+1Wol/uLTs/vN
C0ELfy9g9rh3QkPaub5WgaX7sWVttDTNTI8FKkXyvBj/N4y99zdR1cNHZl8/hK6wNy/7OgDZdB64
Jcdn4D1U8mJcXddsMZaUe2LGBZ8PD1HqyYGJg/R0+BT6XlDLpF1N1VlOp++csqP8TJo9K8eflwYR
KyPAQYmIA0XJaK2/hPa+45e4sA5MuYMoQfODTU7haxR7944m9jQTNcFgcvzqgRN8brTOtGk8ElXc
JUZtq365NFER/HHraq19hsOTGJJQ3zj6BnHhvPQCVWYYOXnqvQEba6r9c3I/YjGJNBNtry/gCMRe
EzURT12LpHnhY5Z9O7ahKmetchR+Su5fL5rC2FjedLe63kuLjHk4X3w5AplMqtjgSgcv/WTMGL0g
/yQaMc8ZbdIJYQ8qhhKFaUo6DYeTYeyhnesGT/qN0eEOuSBFH21k4SYzmr9mxwrP5fzbVLjBKedn
DOxNIDP0LdYi0gWKb41ftPDwrsTG66hpI/n+57C4GGKV7Psx1okNN3mKgGyWxbN3jeKiYU/mctIl
PABuwLG20ZZbj58mXGENaN8TxNDdq+UX91x3bMSWcG79NNUOKm2qHrBA2KGAjEs7gUpR6pBtv3Il
si2jUuW3bDTIY0hGZGdQjkzuZers6OoNMNpFcAO6Kxy0u7m+z5wlZq80rJlyNOoQpS8mM6bRvuQQ
5SMqiCDO5AObrkjlDD/gr66ccm4LnMuj8hK19eT+YtfQDoVY5Fp/JQ1scRW1A9ko5MYaEHgCbQBp
t4bi3fm1jOSGpcMy+ac1EWBLvTwq4TYmSRtWnL/8fHUhE2aQ+K+tNW9rlfKeM861KEd2dG9l9M2x
UaYF8W079ZqfSeg6WDu556R1BaZvdxAc1bEMMlhOvVSj8HcpKxtky9/p8VgL5Xbvuw+MMPEh+sfx
kSnYzWuVhBxI8OJmYDtmTpjPcPb8C1JpmSDYIpWGD5tgOXVFNVClX3CHm3dIgdhx5MbFXSNqVsgR
o63UtRfhycmwCOp5svl5cZ8wGgvJFk2sI1/R0Hbeal/kmtQzNTl/KOzyqAFo0fXLebIJzkZooJrF
EP4LNs7TpztIOJURoMH6xfRM++CsPCj7UyzCIxDqr7p9iXMeeLDJeaXAjaUN4vuQo0euwC/b3zlm
viwVakWVuNj4fiL0QTviyLXxiCCJEsW4e25MdxQUlzNTb9epxQ/KYWz0XcHGWKRBGBafjD5tC7bE
FzuxMm5WWD7UTAcqHFOw0JPAsMkVPJ0x1kWhXmwQ18xRDrR/szX4xt4u0De3JKB8dHblabddpULw
/p9vXKkecCBHxbaraEuv/acaCw9UJGyNtT2ELOpiyrwey9IqZQcNV0IADLtoGvixd2SFsTL52vyM
9H35nCnZj7KlQwzw6Tidij3XxvcqjwoXQtc1S72z1qxv8L70PNX6b2UocxU/tJ8ZwbEl5ZOgEEFa
/HDtkBNLlbKZHf52PBy4P2xUjxm5q+RoNGUlfqaX59wRWpqAWRPS8+ujabAXDlsA3wcRR7AyC5uM
gMPEaeYZblVFHklWYz2ZG10mAFcNST7c/NrEFyMi1FwB1C9E7TjXnCudEjKrfet+cN1YYxSxMG6y
av0Sx3B5Qi82KpIV/H6yvb3p116fKdEqss3nD/Npyw7GcMMA4N6EIFAwT1mFCDCbcZsDQrG2HXk+
W4sulyHNeHsGbK19uS0yPHDzpqqltjcAJ/ErSZGxT3hrDtiIZcn4tKVUpO7j31DKVaw+t0H/sH4f
larxz+bEjSny0OewHH5YfzKSsYKLiGek0MotnpORSTVzfM4i4qzPmW9XnIyZ94JFeYTyCZHajNY4
WZOOOUO8TMDTHxjkfgi7aFbmg6RMqp5rrct3eo5gbEvJPWF4iv8F6UlM/zT1zB3bTavYgv+Xs0F5
xYOfnO3E6DYAFC5OtjG7dm6hZfwFWhaCE4QYNw0pAueYNkqYYiBCH7wPTvFL7q2mPoPXq910cuPR
5QGS5SM9ekN3auk4pMGnYwrVKlF/IX3Fgx18SucJR1lBr9cU3l3aKHA6Or9RtWKzbJXLyYFY165Q
Esh7+w6uRbfLHj1jonfBgL14b1YoYsDsv3O5K30S6qPVJqTaxhKJU9q0PEhWRxJy/eFN+GD1RO9N
46FIVC3KrpWVMg0gnbqFvNbEWcQS21IxzmuWmcKcfoSiN8oFSrJ8fcJzVJN4F8u8fMDaymHksRud
vRCmQEwXWC4kUixvlylVEyBJFs0jyAgnJOki69xgNR7EbzT4LXehIyJi62EJCwq4NercHyuq+YQF
VXycoEWzWhHma5EgZC+olarUvpSQ1OTiRwHU7o/gKX1/eeqnJ3eXoGO6iUkrM7YUz7ZpIbTYp3mg
DSE9cTnM7B5+WVTVp0Nyo54JjV1BpxY4ZZP6IRQ7UlvluJdYCRRniyNNTl9PfR8rQw2XA1O7tLKO
1u+uZK9FH6rMLsy3967ESkPAwh4byQwMwUnodF8uNcA4NOXXxWzHZifs3OMMchAOc2iJ8M9nfAjM
fa742oIlHIwS/tX2oDFcysTbsWBz5e114memtqra6HHdCCgO8HuM+nOYTG6jv/2WqZqB8AYXiBg7
uqmLs/BGKt/8KWor6e7Yx5V0fn7k8VolYwwfeiFWV5Nk0/oi3Go5iQ2K+P9RoPw60lIBDAiYFkRh
08+PGRCwDeQauzJrPeJcbWL5LeahccP28OxcN1w0MVyWdbO8f8MV6GKBP7YvhfTvDcwRSrjaegFV
AWjcVZxLHY4cS13Gt64p40cSt1POMDaHzUj6QbdD2SnSVGREgpVx5gQApW2H9w9EAi0NOoHomAoC
sLKFymIC/umVNqcJq08B18sZ8bZrGAc6cXWZ+8UahIABp9egZ0e/0XlIo+SCy3nrfukjPlb/kRUL
LL+TYeCPG0Z1NRujsFJxXKrNRfTX2xDzTGA9OEhgbdgA2CypXNYaYseMrWNyYvtGsWwyl7sPIPM9
V02uWBiaStU8/IPCJIgtdiwpEaOER3eOIurwVJzTEpPnTJMcNBe9rZ1zIUSF3mXEc//dtUS7zy5N
UW/EmJ+OMS28LXh8IcVwRLovZ8cYj13iU7VBskwGce8odhiwBUBb0TNCtmKJrRihHN6h8vuypNGs
aJrUxsq6LBy9DPDVqIj5rm0P9Fn/BWZ8QnhUzhBO6h6bMaZkcWZwnT12ifiZ4SRMe2OkPdubz3cd
dzufUKTWerk0sT/wjPduVjmrPPUz/rtBV+0zdj7P4ebHPalExOoc6snGI+WitnWQZ+EdmkOhH6J3
6rFrg1AfZ4xefaf+Zwnunaub6XGoNKIkQjuo9mxqc0dPpeTDdGsI/QvnDojrm42B9WBI83nu3d0F
GEQQuSuF0CG5l1iqms9QGcJsoYS3pJikBNmlBC9uoo422mVhpDsnHeZlqoJ//ITMOjnIpzB7H2zB
9MVE7sUZeYtqrlDGff+zhLn8XPeRXvjZRGYvWPJhiIVxz8KbMYBuhypF8qvCzFA9d1yyTL34nsH9
7S4xTrgareoR5i353MDRxz/2IS3TfyT4Y/xCaGiKlr7mMPmbYEkfvNk2XJzwK8Y/FCHYrsWBh4q/
GsVr3LqQ4b3Yo/POY4ldJAAP6aL9VLQtGTCML0qI09RcEW6ph9+7W3hb96XRJJSMrPfh9inENKXt
Ld57mpygkTz2YZHKgCv2QWGk5C6ARhvcgdZZ33HlDq9f+SlcneCGBCRAUsFAMGucjH31+3XPVUl9
NSWfYM7KjETnuG73pS+DzurgSrWrN0PMdMolARBg0eZNjo7bxaQk+W7FFO8wkD+DBpSOYi3a337G
EK2yIZ9AWHAYXxI45RY/YcPdDe/CcXyDHcRxYPSmuzKGBH7PiCWwKoobwcO8mFG4zBzPYqV/ouxf
/4/EtKEefUw7rY4y9RX6weK7Hsc3PtA1+1TvCYhtKugHJLn9KXH9cKVU1xjv9De0lWJQbk+kmX3U
7L8n1a975lhA6g+KAwFlpByk0fMeWh/KPYqkTcnfbPFtOzA3iDrUmdQ3YK7aUkNTJlkxst4qeuUK
Xx4ktQroWypBSIecW4VxwzvgMSFh1jrb1RLn9mrTOtZS+KyxpPY4DOJ49MGcS4R8T9f+gTWLHDgN
JxFJZU5fAH7GRbrAp63F4j35Mm+bFi7Vt691LsXM9P4I2/sLdwo1W3EsMoeKZgxYtJjldaq2H3PD
VKzh08LKaa7rEAULD9G3JO0VOnitlpAELMsM4/Al8rWNl4q9T4jkjJkUw56E4BNTLUXF34zRACmh
3zpm6qRLkwsBMrGogw8JNlNMGUd9kmfw4QkM+FQqzbFqVjHM4NviHHr6mFqkUdcJyfA8IX/dXxM5
xECZK1thgkq+xzV5X+XP7FhSgd9U6sXqm+p3EbSyVOkFO0Z3zbkMH/NsipFBz9RbyRxSFIz0IxB9
dAfxVNYnrtjwDoWw0S2/H3BVC8G7Bj3J2F8mNm6PpPd2Z3LgysAVkt8tHMYMKhkw+nut7vwQ3hJJ
edBhEA8SKhTUIhfyaXG874l5w+SeFhijwH4BkiWoC5YAUcgH+ZLXuZIhe731+u/wLCFLfm5rWdhw
v+xRIirrNUH2zABml5sVtpaQURxNblU2y13IuOXqkukJn+bBTf5OxIH+Pn8AZk28how6no8hVDLq
/rGwRLMlA4kPgHfm+iityrPv8hCT2pwKS21MFf/aPui5UqBFduP+dS3en0aacqytSH8czoB+IUUt
52D9EY+Xc5y9TmVbyW8cXl48JYU39ifW355WaqjeL0V6jClFoEtSyAS8J21JRH1kdKF3MLlpNN1Y
dKsubIJfX8YOgPqaVYJPeoJt+vBr0NMUnKM2oqMLROz4vk9sq09Nh2gu5pJgw5TI/mde2qhmVl0U
sEBMSwHqZa21K0wsMfXWb3xPl+nmaCkgv7brCoy9yco/C8Q0AMQGiY3KNJZkgjwa/8ygadM2n1+z
0pvEFMqUVi8hkUAmBKRFEsA2Fax1mJAT4jfW6YDJrC9haXcoa1ad7c/57qztBlkcy/6UcgOdUxVr
ELpnqnTEAzAoiZRecxqY0Cl9P6NPZt2tXagKoHm3d3Dk2PjiK8NSWr+qC+9p0D0xctORkmTuTe0Z
R/HYyiM3u+bSoCVoVz33g2/EhCy7H1mYKGL4A13ZnQX8Pm1KQqwFK+89RGopxr9gfSLtiT0qGRRc
trxvg/7I3j5KeQij53/wOia14kNW5aEozewugdudvRzj9E2tezVMdeDCekcyW9g+sYJVHWinpCk/
TGmyUHXDJo7PaYzdy/fpbHne0aSJJu+8Nbvml/zmz0c3rjbdHaPV44MliHpYqiqqEdQOGkTE1bUQ
a/pb47q4FDw+YHl61CL1Lqjl/9VPeL5s/37K+zlWjtDbyIDZnGkJaDhAQxYWBdcVxUyf9Xzd0EQ4
OnkPJj+Casgs+S3GwHL79bqjW3jhY80NVMP3aWPPUkqXBz1tnnjuvqT40CMLy1W9DAst0L1jX4Kp
JrKwKshca2I3WazF5wY+YLn7iWYODOvnk1qiONlD5ivNc8T1X9rBrskeSmRADdmy9WSOiXdkaGAA
P9z/V0BSzRFu0eEeWTmY/bFfd+pgxbiB/jWghGu7aDLXN6L4uxfO8ch9Ic/RueYJN/2QK5cC3jas
Ab3RcFglCh0qzuJ6V71SPySEwLx1DBhgbOBD9y3Mz0LfeXL9jthr/d0IfT3STknWPyQmHLodm6Bh
yJIbPOQmabetliK9toC/XKgM4wLnJii7IFq61X6C93b04CWVnsCdapZSelS4zPLTIRMaq3A+CeMg
nAMzbLd23SfmZRfa99UhRzQ2uDmsyGadOByFmD+fyGFYiQPQ2nxrPjyogCdJlEk7zabH+9fMsLs9
rVALy6rITXlFTd+craN0eBtuDEOCbxzhKlMDnO26/0CXBF9U/t9ke6Wgfo2kVD5PhDDYL0tKsPa/
x75bQX0BSni9R8fUPT3uOkKwa0NYsuUI3cLwj3gremAwubN4s1NiLOdyagLub1EOOjw6tkCj7SUZ
mwfPvEHoCEH48pDL9bucllaK0lLvFHsZ/XkdK+FJJlSxhxXjg2LrKwDC9gqnitywS/Jg0GozF5kQ
e8YVh4xqxOzyf99JS8xxYtQXWfVcyjvrgGbmyGkDsL1cbxU18y520dHr2UfOHaM0bC9DNi0vhNNP
Or9W1WLnf/phaMjsO3D+/KYdjcwffJ3IRMwdQwDpVQ1XBVOv5S5DhL9PGIgSaA/ySWgUPu+9dcpD
jf2CgzXy8AZvzdkHRxko4Y25Q9cmsbNcWqMTgr4nETlWNfEti0GQB6NitZiD42rupst1pXklYE8Y
VL8fLimWcIFlDTZ/vWdy4+ByJal+5qc7I2QyGUetw8Urp4aHQtqIW/SD1DBGeBSdBGFpdTKyTKm2
9faPXIjnyPB5FRGUtj448CmqaW5DdlvUuU2EJ9FnO1t24x3JFHU5KYzHHcHwPj/JOq5ednJ/9HW3
vVB/HeU9+y2acY1oBgxEVUbKFss2SyGNhVeArleJ6RC4F7iALpps/gMiviWI+nWxM6gedV38OMRu
fyfyfeDWvySxS4Oc6NgCP400ztO9eQ19N3IXWjsKvUX/ddwCX7uNeURPnKuixME8A0/bX8wA+FvV
pwSjTLxDXpSra04ehzFh8EqZY7yEM+1X/nQsue++lyeZL9AX1LKzlnjW3DSTELkzNy12wtihyHLP
76cjhOBIGZfP0zkWSPuY1nqm0gMbL+9b1Ib4aT14ByKIz7VWvV58xy5u81dMSXAkf74bx4mNzWNZ
iHJyx6eLQvdCcsjlif7w6Zc61F5CpcDOBR8AEJSZLxx7h7EfJgGkv7hrABlXTov+XTQXNp5pU9C8
i9ontTQlumovxgZ5MIaok7urAeRrso4+HUtaacPCYzodzs+GPiGmhJ5s+AYqYSgFPB4effTqDlJR
uJXfMRyHdIZ3me3UamjH0x1o52IeE/it7bFGMv5NQK4TTHn0m7I12sjo4u82P6ZHnjLidCesh2AO
FdivxlDiag38c3Yk9LVbg78hUVBRs560T2JAYXJJqbCXN0DTp0gklWC9bebgsfUmKdL07KVkMl7u
9ck0onl0gjMStH7evMXXVk54T8LfksYUfIj8QrVqZkJLD092mzljRHVrvK3LpXy3bNsQ1o4Eywxe
sWZD5Xncf1cLQH2LtpwLGD2e8p+3s44DydXDyqTY4olMBGYtxHd8yWv35hgOC1dETJ+5zkRdHF6n
ESVv1H5nd3q/R5keTUnU5Qzq7FEmx9tvQLk7D7Dun7V2SIXkNz8vxkgFZQCbz+TNLNqAMEQgH2AE
aJLM2bPpswt8nOjs9p4ffW64B1obDfctgJ5DNHrVPKAE/JOThUO5154WNlOBrEaPtZuWk0NX8dz1
uS30uqueGzlZqB698149F0l9qDkfTZoLJ/LcMusk1wC9rrZNHOeH/HbOC1rV9Nl/wkrU583Bt63o
7AIbPOPlM3C8U6QN20HbBJDlyWckRgT33ZBdAiJVT0NHe9rUMrDm7na07PgnPWDdRfgIZNAYr9E/
eQfXeXxSIxSeum3514BZHaooaXBD5/Lwf/l8E0JaGpHi149A3hgZ16+aw8s2tT6FvNCWrVp9hbS+
uyyTfhL9m5G5ZJDss4dH6pviU6fjdXMI5Pn0hgsF35Qzs24wMbcEYT+9TMkVS27EMW2WDxfF7xkC
ge2xyUrWEoWh7AI3J1+orbZzh9nRkuOd6QL1XiDbityhBB2Y7oCWU3flhENMxisrlVGqlGAd8Koi
+k35BIKWJzkfPJCctlu47GzGiky9FO4JBw5+9yzPEZ9Rb3kSRgzZwqfZr109NHgpmvqJPI0yOVaU
Bi+w0ae6Q0SN7fhl1GXgyPvYQR5c4v3dN4FOZaMydSmUuEKGT5pbAzihY8/2nea1JIbg7PTUw0mR
HBvSdST5t5wt+hdVWXoXFtpylqAl2hdIH1J+vpFG5c4i8FJUp5mTrwaTGd0z9+WHbZzYJZ8rF6qV
Q0Q337AqB4cTsbXv98c6Rc97jMDp6DNz7gucoR2VhuNds47HMxcCmjU/TBa32cg49c8tdwqcaZWD
k3AIGsI20CN+2PrLQR6Q8qNmqETZCoUch2hNNrKZOsGDLFLx7MV0d02OKjJ4MqXCs0cOp+/zVEFs
cH6ZEnCCPkjVd0hHrd9pEJXjGs5Ti0j1PwYmr0Cw60k5ggsleVtCIBjummA/ImEwa/5JmLsK8m/r
7HU29VyGLhVtrC/vJl2U7gFWCkJni52xAAJWTzDvEhDwmU0EMvURGP0HHdQBOaWLSdqvtwCaNZjQ
fYz0tIiywX8Em/UPaIOE2kXLc99fzmXUoaPcmr2XCIekBpizs8j0yRosBafm06OusFUPO0BUWMA7
J+jxLnuVppl4cEeOJeJ/rs5bEC3EAVi/Tp/s1zMTmbqvkqgJtSCGHaiy31GxhQ4CCVxgVy+xLwtp
0tVxsihk+s5rvwUHQyoAn5N7WU4aPrCdKTHxZOXUSFxCoj5fYNVBZ54nBNoUmJG+Qdj9T1e8zsRH
uhSLslZcOh02BZCOQ8XAhBCtFrrIxnGdTvcGBLFPo60QfB711iWeqQJhydgw8XY3gkC+tKP4ui/t
OfExZd2f36KpBZVQ9q8W1q6oVKCpyGbMdipeZDk6eItjLmrY/H8T9DX7xdhYVcRunF7gWKWwye0d
vssILtNU0h9WCDhlLXo7qeG5Ojp/oeo0D6k94NR0uX4l3J4qhjJIsJbL+s1Zc5EizoJd2WyDnGdj
QZK+fxVCmg3b4F38NTH0RUeV4jK+PpEbg9YfLIuu5i11q7any73zcwgZ+QASzLzSVhdhEJ443E/n
N4pNKdedeb2P3YvwjaA/pOrRwWN+jGRHB7WlG8duSf6lCcJCi6b+P0/nwOZ6ho5YYXDN2tMFD89U
+Zv/DjUFTrYiciPw5Nve49gEhkJPf8dVuT7dX9CdGE4rLNC08dOR0m9xL70PlSr/pLdaORsjIaMT
mw3lUpeJCyR2m20BRQWPZwXddQu1qxbvGIa2M/qksd6qrTm1E2pLaECBX09P2QTH1tJU7JyasTSq
Fb9PAm6QTLLFowXbgOXEOQnzmZnPl90OBsmtuLmQohP1ZN87hHsRpjtuMqiNA4P5FHxwxe7yWLLt
UttG9+tozVkHhfENF/xZzh3mlm+ya1xUoIJTaDCahilXJ2cIZe+GV/u9x+8woV/6PnR84kn7zG0z
r0HoLyd6cop3S8F2xtG0dFQQ/0bkZVjo7OD2PLFYdxxMF4knZvUmvrQN00feeJ3wG0TAGoLQyO9/
c1ukFJ7dor6yKmGBv+eADWXZrh2kNdg+Fj2sdky3Edpe9hk8nwigUpSw7aHPrZ1ETU1ZnAfKpc5k
emNHTsmgGuDeHpCx46tKjZM7cu5IbZpBb7JdT7RL3rzrtmmBjqRSzaLAgfaYQI1NdAP6JV52f1cr
QnX+DztoWdjdicRlcymad2hF6s9WRVkAYaZvP+RKZOf1r+4KIjm0feQU1VXoYaetMjEAq0Q4irYM
IEScrjqB65tvd8wjR20NhCITDZC155/sICUBObL/dz18p5+7P12WSPDpenDHxxms3XoX0hr6Slmw
V4TVPXP7pBJPnX0mIBJpU0cn4a8NxdSdzqCvzpsSY4xFY6nQ1Xv/S6VBsQfvQplPfx+CTrzKRZz3
jX+sF29x9NjNNKmIYNMKmVntoQm2qlwJ5hKmRGyP95xlPvS++4x9uup83mePTII4B5TfTv19OwO5
g+N+XOmYyC//rMRC+4GqC4XYFmpqMLon72+EeiBfpstLDD4GjI8p0/X7EMab+QaXAU8/nutGu3GA
d2/hb0FpPQZ08FRcjqzPcYsnDELz5QUUNB628duimyxU/ENEkCP76RDBK/fegmFwnlobNiHIHM4y
bbgOAx1xRfqPB4KMviw81d7kllNChlL/PNNC1hXJ30IiciRj3fbQu7MD0MVTZuGSgc6kqz5dy+TT
656IJAZPD+mmHFQ7OJfEgg7T2inwmWIFavtqOebLZtPId1E4rj3ZRRrLYZbmwWtXD6yFB2NisyYL
zvzSDE8GLCO2l6iQWTmQHFL5G+IZIztXubfKCmEXNXR5dxAX0FlhUqcQDnDNHpoC33JQGIxZbnMZ
NSi7d/DZWULvIi4sJaXr7jiJ+tL1DVHyNC8iNoXJ91Wjd9k9fuK5mVj/qSqCSUk9+WBdzwTzbgMA
cJ2gTFXyVh6W1qjTz6/g8dGB5XCqw+UfCb7U3h5GvU4kevnSZsz+cKTVFp6q5OhaEFV4mn+q4jOu
hk3UTRpeAh00PQ+LNAKg2xVj53MGBUmn21T4bsG3t8L9N0HE9KWp6oFjm+ozmQeLZR22Xng+Tq9G
+BbCvNWLYBRACITopoEuTMCcoCwLQCqCUKUNcsCDdnekfgNs2iQvlBajU5kywRkWEXcwPcvHr1ce
uHWRLIzibyWY9au1j4apoiGk4sTXD2BCbJQnHlp7eGb9tMt0hBkU0mFzT+ji3RkFxhN5t8CuuO2w
pdf6fuUdGYABYhWxwSaOHWwjdQ2DKhtn6aAdOhmQkO30nk8OuZGH/UgHo8APN2FXh3hnXSf9UTnu
AWHHwGQIoTfDj7aV3tPVXF+hYsdHmf4IRNERRRpPJi4s1bykT2yxCFavXEXiGxGaX9RuVVqCT906
HHpQJCh2k5z7Iht/Ht3nzegLAM2Jutgp/fWvpUIsHp+LXFCa6Z5lDtgm7UoCrLYDBZzcWW4ZS7iJ
XqbQ/gU1ZRkH6cYR+cxxsgUXgFUTtfJ36QVWCFhPXPvw7YD9K3q/CsB9iVpf3aIIpCud6uqKUHO7
Z6uzNrrngpMTw5WPQ/orOEUvUUrDYznDG6fd0QCQyMFb/Ez58avnA6csEtok5YvPO2fyPbgiBO3W
7CkUTo9GFPXZZiACNzGBovHCmgd76/01V0f9Dz6ydW5BreTrFYSrs3X0Dop60HlFSsPG2jI6fzYa
HpR5RG2S9jytBBLTndCm0W5QbBDFECOwBNHSYJdDdLNLPigylvqntfqRbkSnFGB71k42sGLlMARv
LIQIWnrghK1cyjdKEjBkm+bCvOTPZmnl7Pz2yDC33SoA8ZbaC+Ln+B9kOvCfFRpIIqePEHwE4tls
Lx3xeI2CkroIr/NSvU1Saw0tQ5DyYpm0Uojrwmw6dezj4T8piNbaxzht1xYAPFMy68Sa8+LlS56a
YRfXoTSL1h8iZhxH3VAefw+/srU6UgD48LqbW7bILFrlZUjUG12CxGHsxQAIlpcgZ66ix5kIfg+F
wsKhI9ia17D+nWu+QISSeuljppO2/lc+UrcDuNoWvi4rnBH/5ZKGw3eTbDWRoHVIoyk+qtpgHSpf
UKxeNSGN/jDFVa4Ds/1O+7SMD3q81r7nPGQHpQ6Cal/osSpp/2O8ID1V+ngVDGC9j/b1RfsR+CU7
EwINWdt6Wy4uJdrBPlgTRrB8MT51SxoO/50k+/z68CVAeRkXTaw8G36foUFEqXKzYnysCVf9v3JF
EEFHZLkjrFu24Z2z3G7adjRdDxhIMxJoZ1m0g/VKH5Vi2M1W82I2OfNDUDOFDez6FYVjeuZRC3xS
z9Tn4uwKYqDP7d9tzEoohzsIM9El4UzkWBCNzko6zeWH1mwCDGMwSC/etBhYHJ4yefVs6vmSFDN9
DmulDWztM8haBAE/0aMqMkJanppZggdo89J/647NfxUmTv05ov6TPBtLRN1BDg4hVE090NgE+SIc
A8fCt3+yaYA7MjfnGPbIe8Enyssbp+Vvu/PF+f/iNvL3RttIxMQ/PIR1W70dmwMlBJpKL/1e472l
2YtoEHAvPvt7H2wSzbadrUC8bstUpl8LexdyhSxM+5BUG2KTw9BWX5NK4Vk2u2hadNofBCTwjCq/
swNWvWFKSExUD/oUGRSZwJ/ZdTx4vbGV2gNsSJnOC608Us32m9aC2OmK/kpN3DFOPtOpgDw3ZJMx
QR0meto8nvs5oghQSQGWxtXegP0BZLDWgiEzwAZ+SGr98XWYbKWw8XpjZoQVJlpqwwxD9lDnNmvu
gYOMR+7RW5vDN0pzHeIKyURIsEjt5EhulrgYAPwL7/u7+C0AshWeJWBSwOXUjSqXbxYAKjA5JUO8
IhKqnoJduuCRv9Lv2dYY2NNo5HEsocEFISaPLeKvBRHZWu0kWOxJmi82P/fvXJga7HuqTRvIronL
gv+33hHo8fzCdI1vovkgug1NcbxQ2+MjIwaWl9ArY6N2AhtVJlAIQ/7Ovk1+p6X9kH2y66cy3OWP
+3QXCtJizDFmmXyTUe5F9mn39XAV+iFZkz3beK9XZUSZTRJpUqwwn8oe/89i99TPF1wvay8Jd7de
AHxiOzxXW0pzXhwwv72JKeAU5hXobtUmVVHJkIzAnJQUpx/1OSNNQfPN47IdwWg1z7KzeIqFJuY6
ENoVkZuqfA1KC3FawtGvKWVfqT61tPV5tlkQ9ZemfLdZq/pJhHjC6cviiFfEGK4q507cAZq8OtIX
llWZr1JsYCIaxb3/sz28wOJtVvWLNQnZhzr3aTLOSzojUFLif79rKbe097QfqQmWb0qdJiT5rsoF
XtKz84eZq2uHkG+N7jP1Oui2SuJKw/AdDYlW3Dbuz9XybHW70JHAoljzDiyT5rC46oMjQCeNRCwS
OEho7Cnu1u+eJujCnOyQU/KOTsoOkZdx4tAe/32eY/eJvXVEt9qZtHxbsEcbiAu9UZ3oYY/HOoLP
xji5kJmehkpLjvYwCUz+wb4u4D5HQ1VkltcrFGWYtKem9skklMw4gIVi4Q8U70PL74gTaT+n3XDR
4xP0p/VwOrLaD2FhTlVlZtWcgsgIshjvxUKMGD+84aPwCq0+jFkD54+ZXB4e7mqI2bN7T4iFguof
UM/vxPFrMTPX12pWE1z6qV8cyLUSUqaz8WWd/fU5/XC7a/8+Z8dDDXAz3sd2ojdLmwML70ntx0SQ
Z3vGj3xUska2nUz3i1J+buZyxsgOYU4cM4IQ7u+KuhUAzxaHmjFpXHLIibqaqmkj2oeAQFNU/9Go
51OoUJZe0woHezi1EV5jGT0TCBFl9NCMBuP8ESvkd/RfdxqNc2Ij4iXhS+mKh8NVxlSTnhLx1Cs0
t78JOuJL3fEzRdm+J5+3Bkj3RCHFesBt/7GvRbdBe6IxwLGMHGGBL6ww1DgVyzezA25TKMt17PkJ
QdtNCbchWHbrSVaZv8Xyk9KSGJODB67qxwPKGdxbkrjeLLyz6TcbwrfU5N4twtHyIcE0OHVr5arB
xwYvqxp9cKIpJsjqLxE9e6Hf8uUwdhwDqMIfwQeh3c3oUD2gFqeK9LMhfnwAM4dePzzZ4ktUbr69
9TkVlLRDT6/NU8N66tNgKBUsfCgs7X2WjuFSdtKLAQuZeeMBQ6aRorfjc6fbYsRe2xZmwjCBlSq/
j6GSXkesTJYL8LpU+WnxSxJCQ1mW34RNZdH2tpZpJfVPthovsLdKvl0CFfa0M++fwo+IDPCvwQ+7
i2HrFBkiTCeG9hzx5ozqprgvbAJ/MqS59DhloBi8H1+irsnQAWKVt30sqidrwM8HlbuyioeeRl8F
AqTrlN0DgFJ2BxEbEWjBs96lYU1Ge3+Wx0AN5mk2Gg0t1j7ky703YwsjE3V8jEpRcpl2nNRF8mYq
rJWh6Mh1uQDNntZGibogfv2m6x9fygSo+g/I4uMZf7VsfCEhiJ5sYNC86PQ6qHzrsujhTHjU04UO
dgAgRYuQmi8Z40EWPjvARD9zlFCWb4ncJB8BBLXQ6RxJuKIdXZHMsNqfPbQdH/k3M8eRh0bcr4qp
N07QP+twwdmfSrzA+dVp0U3JF/CRxBr/09zXvJ69pvIpk/CKr5/MsudQTCpAODUpt3tgK34PQ8sU
jkR6mk3eA+RDwflrjYVgq+IvRj7laWWY908TqPSP0RA3luHfkK6WUazSZfl5g9xvvA2HZNLqV5hw
s4Xdm+yBORSiqcNaVVj5GtIyRGFvVnt8CSMMbpGoGXOWK00j8melCm/A+zlswiD2iVO50dbWirwS
nhr9+T7cupxgzIx3aittKDC6MBsl/SNMta/2RbTsUubu0Ej6Wlzo2O1+PXreXN3pKF7ycVmTR+oI
0eZr7ZavwoLrZlajKv01ePKNDwe0XIDjoIlX2GZYMVGyMW8KhlCpPz0qUYPnWN6XE/0sgk+1vphc
CwI757RXD10Aze3Yuvzw4i1vI73cU20I1twJKouaAgu+RVVJWxZk00VvGSEQubLQGx670i3H5K10
swxJJ2p6dKAZskkjnCzI3THmcj7IlEH+yh5OV/jwoTW50Gp8sMZ7bJ6ZQTBlOtZoyBAOEEEj7Aja
LsZUVZLtn7V2SX/PTHRkuKhQ+1smhaH25Kn7kp3hmj1nAl/4gunCyMEIh1/xeskURPuRnK3ejuFv
zxVNTO8shrZZm2da1hbfguslU035+AokMAx4HyqLdsiO/7YtrDYovOG0qvJ2/eQFssVv95KvX2lz
fLqYajmj080vLzzJYQT5/GqLg9dIk5/EvMxvcnvzaHztjq9VZ8u2FuiEITvzcSjTDTMuorauo10W
mypHo4oN0HUDGdqTCqI1SVI5a6ME4pNGqpwIIwUcfDQus8Ij1Yp4M+BuCbJRM5xWPcMBmlOU6rVH
oNbzlLirQPaUM0F3WV2KGmniB09QDY1v8F3YVmkCg6GwwExTF2NtbOYJYgMb9Hg0t0gfRcyQCZR+
tBOkRId+ZYKNdjbN06lMkpETsNyI1WwFLw67oxR5b8YuB04rBEgdWa2sgRO+IGSlGeAPJSad4YMm
Y1CgiRkV8olTwRQxq7yIqLXkqEkRgp/MwzKyE0ArDu7FZaQ2vgP8pwilhX945HPb/VbwTer3LVqE
SSYSIF5Ji8qIcxFN7pF1TY9y9USGG7IPBkgFyvbHXW+GuOFVLk5j2vgwra/1l4sGaA5NNVxE234I
IaZXojx8LXWVdlH12nSb0c0a5Z8Id9ECpJxV3UI0M/Xt+2nFLkSwgKXIZLYwSuSu9OUXyxnslDOS
0QjZz4CFpg0mQO3+gtNyOvA5ONoFKpk2pmcCfAo92j3z2ONN1+83iPoAsB2VRGJY18THjvOd2d+j
Rqh2OiBIJqPWesIDSdU6R3RVju0qnyWyQwwM48h+gowQvM1XobbRw4dVckz4nY3M6llOpuVWyGs8
D1gKpYSvgxyvSIQ+39TSQ6NMYHIycetQ1VgJpMV8+kA26gv8DQth1dx8gEMcDApbKZ5obs4Qw+RA
4/Bwr2Pbsijb+6FBhvYXadoWdmB3+OyWtLlovbjE4cjeBbhE0I1iuwln4dUWV36mhUd4qhmQS/dX
J7k1H1FIqcS1MobzqAlP71euvdT0RPNyx/lx/Q62Wis9OyWBmzR+D87BY4eMM+Cp9EfJ9Wd3cCrQ
SnwyI1NNsTXVwV8+XJoH+IgcJqjohxbBwMIHYLqh+adP6eRtN0PO227na+UIBJJw8AWMZaqkgv4t
Soqc2Ok502JMaHzbfhIe6UG/ZUnDkXzhCIexaxqfW9IOS2qERbwgZ6KIE3OgTj3nZmOy/ha4FLct
i7FYdU6DKAE1y2CoGhColOc5T7vDiZaIQsi05rKADfan62aH4YlKmGRgk3LdKm21E/zLw/JY6brg
I2GyKSePek8mGC3/iCvWQkAiH/yaQjiWdDOgrCXGT8m8ybQQZRxj15KxxmqwWnfaxFsMzTio6JxT
vK++X3VquzWPHdXjLm4hWCtUSGVcowk7NmcJSRL9q08tKdP/62dVAUcPjoLKNxIuEbN5E5fEgi/+
KJ2PqrZ5R9Hr81C5QmMzQ0kZxD49WGWRBKV5hlC0P4fYhva42oAYpg7ls+k8pdOLwa4C4COB3i03
cQQTCvpDOtC9v3PZSwqG/R6WRWOtkMT1R3WnysBvoRW45U4wRXwF6uS2Nc+lNeNiTxr+mpMjpc2z
Agal+hVpZc3HmtRD8yy707iDTtx/gcnPfLUHNoZz0zsh33lmAUP0/ftCLVo1ZC3x58Vm8b0/gQd5
f/CodeCegr3OKpeU9HGkKmm9WVKLt5AGea8GWy7liIwny84fV9uOk2dFkLKEO0njpFersSFxf08q
VwDJTKbqMhIuH5fav02o0aaeLxwAHQ0q8d46dtgUg2t7xZjBnRR1rK6PmP/paycFVzjQt3eWmcr7
ysThCzl3cuPryzGaFtpHXj6Ir5g4R6NcXsJVPITE9FGPwpnm42E8r4ntHef54GRlaESNCXo8SOYQ
wNKf/j9DqMwTJrw0JJGhre9DfpmGEYLpfuc9ICIU448cFxCdtUf1vVHux+/VEXCEAqkyIEYJoxmY
3fXfEifFHh+XW+cfrt9gTYSAh/n9MjhkITCx9mI8U6gc2Pvu1pB2nX0OyZleSad2r0KXZO0A3Nzq
E4y8UKO28DtCPoz1qm+yj7tY955biPccoGd1Tntj9U0tOH3XGOJAlfis9GfqEtmDPirfgCDW1cnV
3ffYai6RAsYiu4EegcrGw1ec2ofxnx7URPT2zZjxMlp4+Gf4YiC+Q8vxRknCF02v0W1lmjM3v9uw
0mGIKtf4C+txwaAVP9rKh0+yHyr7ajIy0Cvjohbtn5MjQ2znzHeVET9ToBe1J7+XN08ii1JmBCp6
b0vyegOM0aq7gKn7XPNMJnXD8M4ol5ALQnzNNO39YQVcE4CD0Kz4qffJ3iPG9rDXXJ3GNwJesXg/
CXFXBFDZExU/xRAnDLrx1ctWNfC7iG7+dNpneeiqQILXmuiipJQzX4sYc+5bf6PFMh/XcnJWfDSw
WQRBe6S8HLqp96Gqo2sUIAtkeZREImhZ+eFBoB2PoRLqjyL1MPM0I4LM2XAswyDtepU4ZdltrYPO
abhzP5QAL7ArLfw2d9TZfUz1BhInS22lXcRj7bijvL4Sbg9cPUSM+CNrmF2+IFDnv41bspR5QKYS
CoUkd1BthZhDdN8HfsKDbT3rOUj8DGWP9W6YL6AtpNlwgPQb2g8Cef7ElzUrat99deCzU6/9Z4CO
00XJwtH3t8/YZXr33qZPMcFvIRP55KbKE3WwOSLWriDo0470D3K5Yt85bDFa4AtIMOwRluOK19yu
L+oPPOTZ/gkuSlV+B2Oy1ngMm8V5GFuq8EID8kDgNACSMrvsd2Nz3ZOvxz6lO9s34X6XHtgot2SP
ZPnPZ71nKZNPnuDoZDVwzBMFVWnKtHO4zEfV+2m8y47ZOrYPot3MFgKYvMTajze1CswZ11u0FNai
H+hAIpFx5hjVweSa3GqlakF5HpFPmdxF/QbW6SewqesbUcltP9GswPEWTCg4Zd8BhA+a2LHaHGH8
IzgELAMQ61M/mJKRZLGjvmtF1H2qR4w6A2ZxgLaiEEuV6sbR7+XaUN/U0KS3NIO6A+9LRAf0i3Ou
8FZtOfJUMew8FKuSOLT3/JScaGTI1M57Xii+af1S9o1n8hz+ibfQPmArDtTirO7CJPjWUzox77Nx
POP36tcKDs41xGgWtepItXjjhKlw1qcJqfryym6TFSVfF8tfU1yB6AENZa2/ZCTW0qRtUAbAt0P1
vRxe7iemV+TdU/MKDLbyg7RmiXY4cS9UkTXZCLTeLmgOsvhJII+iWRyDH4obBqBrs8C+ZcceVKex
BT6BUJt9RqG4SSjswc+oDz4BjIXnlF6RlKeMZJynzjWesTBmcYMT1958rQ9rt2WklToxF45o98lo
wq2O6myKY9lLQbFWYG3yGZM/Hurp9hUc/QSr/m/omCajgBnEGwMzv9ugrKnsdWd5J3G0r0l5koxV
PXDqmFOtTAws20/AC46qf79k7eiG4VVKeAN0LWUObAWWlaRk8FLlIRcKzBuE7elV9OzoUNmQxOLk
AOcpiqHCIjgv0ogVKnns8FKmFqGvMexXjC3asOpAMAoCuYM9ZwFQPgTExu+qjYdvtHlfuqdwwgeF
7LSFhrmtLguXQJ1d4KoHHVdc1mC4FnO9IVrxNIHTDGx0lpWX8HYjh7a2pVp1eI3WGXwxzVvYrrd+
HQ1GJlV7ATgNTIbTcbK+UYZ2YWYICmEZllpDMO0BxNvXwq2ZCOKDNBKfr+jZDZA60cnKPeTYwmuk
oEziYlLViNqX/akz4e86IZOgxV8x1SF8SprNN5RbNRE8C/IipLryhmkUMLGLmmHvs3Ei08/1xdch
qLclLz0LL3CvoOED3a93TDURL7ZRkiJ7u2cOiBRzibvxwqyqqhAd/WWXVHyBpMBMd26+kccrsNpb
mx70dGrrEuofYSlQqqwozkNMu6a1ndveDyzoQ6O6pt3ORGUXhp0R52r1DudL4W5wDsoHJhNyFxis
Zjo4LBfTaq8dph8L6uDNedmspDxdqSBYSDG4goDwfYmctAbqX/817sjuGH4OK/hSj1SRDxXp5KBS
QoZVzPmPwQzTPGQ3wlB5wbcBGmEtUJIFKxPGpEqTwdqWBb6HDV5dNAKZG9FmloExCanmNub7FFRl
6CVKRiX9+WWzP/qvNyZOdzmtt8ITuwIqnuyE6k3ne4KWbMT+/pMb5h8SNkn1bEbiX5GdpX93P4M9
E84UjPFcRJiTfgti9AwgGlGoo8ONxcSLPAsm7tBIdhqIhapvL3ResEH8po8dMEiFQxxOITSkho9j
Nh2vufNOrMTfnm1qmav5M7yLQ0FtxruZ9JhaCPtpn2hBKe60AVPugKkUF5PXb1em3LFFXBmdSKe/
hKSnw1u4Gy0267QaqekWfpIu89gVxnwgbyrUjbfDTeT0GOt5ebuhj1pcXXMYkvx2WK7RyARPoom4
z4dg69vdeI2JAHVTHQHWxOgvAyYZjvoofe08XbcJu5y5NHvW7gTgYzvjCVQR2S3KyOYMyWtYfMoc
43cGEWPHGqlUmdS3K7rKbJ02kWXVGK1BkzGEsW1ElDT/ptxytGyg7pOfY+YU3XOFb4aZ7iSGmhzh
uOII/KLw/XpemkOenIlWr9vh6JJkLLBypVC+1F24nWcfzHtXCGVaLhUg5S/DtYh/6p7u1A2sx/+8
xGaXSGEGigGLo4mpejSq3xEEVY9HY4RoPi3bK9naAxUAbX9DYF3BtFboI1TTVl8GedQlXtg4bbWr
gTKhugX0F3Jt0Stfu3jWSc3Blvzbj4yCmbuGMx4z6FWQT9LhtrVpUYPYHlOF7MrByeKY/5Fex0HG
4g4BNG184dNoIMEFxRnNMAGH4w1pE4Y+33/U5KP9xsSJY+vBBKOcd1blSzk4NFf/n3E78AOn4gkd
JZ4knrwMRRigb33DA67Pm1cPVwADHXTa2gFhVL76d+DY7l0oyX2CV4L7p657en2j98D3XyxTt4Bz
KpIuCmOg2RG69d0BgH6tFv/viWeXWSf4zfjC/e6L64iaiGVioqjZoCGgMkJdHrMOG6p26fEDlbxN
5+gKqSKdE6Cy8q+bvZr3QYTTv7Lwm36rfbw2wXcmJQv7eesIkHYd6q83sLGq087FnwXFYlKgOjYa
OwIF/1j0gHdI6BOs9Y95RIOd/qL1rpFniOtLFFvxa0UJ8URC4lANGvXW6+d6OLectKF7FF+0TFUC
5fdiUmULnsk5FJ2ub9xq+2HrmKtP3dlzg5sJYQmIy6UoLI8PeNmd2gESKgw41rvPTJEvk6JF7v7u
3+sOYslNj9z3XkJEvo1L1LkmGFsHljAQthEa77PmFj/4f+263O7gXrtjSe9NO67+d9oT+P+S5bFG
BrEa1E8yJv1FxYVviOyjsXknkZRNJ/E5YBjn5LI/MGlJmmsbfoApEABXH1hF6e1/CMrTG4UrWG10
4Y+aEqG7nUOjTWekQeKvZRwOyQ0O82O/3J9VF5xuOoiwVOYeYmVXEgbNXCMyiZ/GtsNUwM7BWLm+
bFQc5uv0s5+Jc3g4/K1XUCJi/fRGtURb7BtrXL8JGq3EK2/DCmuJzZh7gd8/0zHj2lAz8NL6/Me6
+JrTAaonELH5Dl8vSAifaZ7k5xUh1QQ1600rwUzsVZfWwLrMVjiEWRiXQ8ofabMMrUVXyfelkODy
naPRlSwltYzQebuQrRkn5g2iw01JRl2KC4TyWM3gCAg1Coo8JwQfQUu4/R1S5te5dx8Sdo3MWevs
0RCi1mzcxN98ZYkpW8usrk6O3HSCheMWYLfJLqMqJExuKyuZ6yvN0EQGrj4kPRMQmLiJHG9rvylF
/CL4k7+i0Ku7a3nrtYSjrqLfQ7XKrsJ1qfLYtVo88BTu50WbA39aZXuLO4VfRSPmg1MGpun3zMw4
X89PVf4BtI4UykRwIE6fikX0cs40DCqllyarthWU93Idv/CxnA/Sb+lgYoW0o/18Qi6qzM/kcqed
Pvx7DD6ubEQgv9uYwM/YUVIAcJdmggZ8qgWfMRuNCNvGAbPFi4f7Ew0TVcnioJm+TLYvLS/Dl37c
k50Xhkoyj2LorwiMg+lWI9xx6EdWwHd7/Je0WuujJmQrgYoj9UWJTuU7/1PDkEFeM8aFNw5GFoL4
67d6IfRfVcDPfkdzUnOgkkiEgWFBq6EX10IO8Y4SKZRKuENJegh7fDzwzlMcGccLtBDMGy8m5J8N
tpKUzvHaKeHcPXezuZoDksm3DXtB03Sol/8sOxyi6hL+FnqCtpvgSi6VN8XtRsVnREW80P7XDUEz
f2ZtA2dd6sF25XiHJlQcIHHAmJnZLELEu9LEC1sx/s8lTTJQHQ5GPUAqbEqJVB8Gf0rWcoOXK5o/
YTpGPfS57wXdXwsORt611pk/5zxS/DHVZf0JkRvqVTa0GTOBtDsbEW57JGNtvYMpsp5SahCd8+dh
2oOvj2af62jNMQSC/nQhCKY8HnqNkl+4QM9l69F6SiKaq4SJUal8f7USab1A0OYPgDUXHK8VT8kT
jNdJrZzrA3hpdOD6/ukwpnvl4DaBsH/EoBp7iDSPIdoqcACxJ9gTbvm5/qLoqPCyGRZm9Vkax80Z
IfBdWiGEeGUzhNpWcgRzJVO3NU5gVVcfnww37VaQz0GUhuKmYem+4vBUB8bRQ4iLTFw5Qhuev6If
3g7hFNM1MBS9fm8QBpKe3HivOkHsuPWA7S6baqbMlP1gwEq057ytEpzox3/uHFcTuQ7ubx/oij2M
LYUFahFnSFASt3mwYlCygvy87i8WuCgvPbMueADRbfbXvvxpTflBq1AeQtmicko8ao2tL+BNUKEe
F0n9sPDmoBCC4BhQQ3h6qypBV0g9BuYuVvmFcLYWLLn7jo4NbgKAsclJ22mK2w1mhbejzIEbdoTt
UnkgQdHdF6nCZqcVZLtm1gpzdxEVSi+E+h/e4BB1HjInYyRhf9m+REUYjGZDdRfnZfwcUGapbHMW
qbSuTIfcjAryWnRLo3WbWpMXa6AE9hWfBzRvrHHsaVvr65r4WRaLf5LOPzuvJSSfTWnbKyW/ZotU
09lykp/nh8kACB2QkFGkljp1X3ag7yPer8OOgI58Ucaib+cuGe53qW/HoWz9emTZq3SEbiyCxtzi
LhSWJVFRMHEkEN4E3Y68GC4hZvmZMUf6Sfd4oTcTbyKutBihl4+HKRkcHHqDs3p3XtW1SRDvYhCl
78ThgI9LXS4T290eXSXYrJC2Qi3pDZHkCAp0FTd0Ykx2qNrWa4ITUh4LzQIUqNROK8SL1Wac8a7F
MgF0Pj3OweJ40sClIvWq4ZQ5jmTbbHjebkepxLkVAkd7rcdRYIhvhruRKfy/xultzAexwu1UU7mN
mJ0/arzaj3v/tfEs3Obm7knLiUK7GOyjimkrngMb+NBqPGbw0B37KPGPld1CtzNgE6/Oug1g844j
Sw56XrPO0oEPHbP/kpihEhTqhMl9QlhdqCk5fAdpXj16vO6cvGAbS04CaJq2fUB7PF3nYzqfG6/k
kyA+uarJjz0qpEqS6zK70l/hKcx/Lem0/WSIg77RHx0KDSk74GOiwIO+XUlqkqFLa/4MEN4Z+znj
GH5EtVs0VQTFa3df8Bwpdr0lEQp+1UBc68/f3oSJBs7BANTB9lrxEKkhlu0/lpGRMGIp9WGT8SqF
n79Oyf4ABPn65PVLT6j/rVGftYJc/pNSGZlDoe8VmwgvW9h8RbCUlTQ/roxBW88JACebD1a8nIB5
q23JuFLAyfdabGcgFnje8pf4Y+hwiCPq2KIbGPgGgk6ahpsc2lfizr654V7c1xFY5pgm+/mFBAdS
aDeVcr/rxr9kqE9txfgnnnrBC4U1f6OtXgaeXyh11Uj1eKsZu1ktVUYS4MYLrfrUCj7vUB0tVpee
LbAs2edNkeVOFrM9OeKTok7H56/OIN99H8kIWQ0JZHCyy9OJ3YbArDa/v8QyKsx+x+w1ibct6XuI
ahWJ6QonFgZFiLbIb2fOrtv81FC4RJAvDGQPcZLb+ELDthx4m0zmBGKbgMWGcS01OMn3hNdvMs+r
T2uWxgKAfGIWpx+4Tau68NozyOQhmYa3PCKa69xPyRGqmL5CNqxWCSNq9zElYi1NKuq8OggZu/EG
ltsTusAqyFbMZtaVVf8F9v4s17VZITBq6sTQ1J7U4ZS98BnoVBfKyqm/zZKGTIF3hdEB+VpwRxtb
XRY2ZMNJBkKkvCgfV5M2jG+JQYmvPDvgh9meOgoiiDFjAGuRM+03J/LZYkFeL6pVm9NZQrCVAYhW
tI4QZmgns8jbsmnYnnW2CwW+P5LoKtHSfJHFQKSVjAZiiAp5lIWxsPF3zmraOX6usPPLVN2UZTve
WMnGXRhxUGp6LRZ18+enHsvFAlu0P+2WPBDt677/bUFr9hDuLrrQi5PsAN9ASQdilrrPHYAQusIY
9IYTufy0jebrOWxowNdujfFeyj4qs/8ZaONiDDfXschkAoa/zFBOG/XpsxQSSts2X+PvkTLqmFfi
4q+CujfQN7u8uti9sgkSIrjQ1k3D9UBEdpv7kcYXLuGX9Zp0UkfERFysKwt8siM9bXlbFTgdKAhS
QGdgsHPSsWrd+XfYBcRcMPK7CELj6PTIIXHQrScUQIFnM3FfpqXp3zHTgZ1+bvZXmxk7Op8eUCkI
kr+Dr3E2N7zZJNAK7ssumO+vHJKONJoYtLFNws/pXc5kpr/EzQRsly12f4H3VV+sod81uDR7rnLF
zgG9Sb4cXN7vmJbYxZwM18Z6xU7dAWgxHZuLHcEhFOFdMtHlQ/zO+ACxvczuts8Jb1xdltkEA0vj
wJtNviKUc1XxlqFdcHjrQkXAHrw/4neJl8jEwa7ZTPe0/LBLFxNOuVC8UFDu4CWQu5wwQcWG9XwB
nW8tMqA5I9ZKin1P/a1NArknpLIuBMGd4zvnJgyv/EK4GLeDhR3udeK7NE8PxSew9ExjqMDnf03x
0f2NGcD7C0RNaEkJXvZF/PBt7x0PD+b8YclFQ4xnPDyI28Gf6HQty2oAQViPc2669lRRqLZZt57d
6KKLKEBzylb9QXaYCYB1nQEHW3iNsJ8zrgAK21zO3oSqmCyTzJ08keFJrHNJHsJoSOf3XIF2HuE/
f7v/YW/vl6VlBc7yCWcXQcEoyUwDkkMAzBT/qv+hgCdx+BGKOHWGlSdxRJpkbsiNZUTszZVe19xH
jDkWzOw44bD3VsK3STemZw2j8aMPvNG0KFriEiKgXXKqDA0ekNQ+RGUmQIEreg6T88LEEpuQH7uu
2Uo4gq2/3br27qPbvo1G2h/GQ/97kja2OpqLLdYYHrLmm3L6tWtgWqwqvPtjqVdpgRZyMEFry8sh
aJQzfEvhl9r9l+CfKbFqBN2TE2LFJhXSfdow14evkinuahW83B8/QkbgN1D1yybvqXKV8LcWMUWs
cf4VKrfRFVyNzwj+ES0W1db6mNDG5+sHOTCRBhQQoCVZVHxdvTPqbsjY4R7+GssSHlrWydZB8wvy
GeAN8tKwj3RsQgnDAXX2cyHVu+LbSy71e6cOlD21KP9I0GpYA40aGsOiBsLjlp6vDSH9i68fM9Di
m/W2hLLDOW3PMuvJzO6x6h1HtR9WFEzls1QMmhvjsbnkOzX8y/jrsFUynTREFBPxYLZT/vlSxKj7
BBuuNskA5ud+B/3Ig/Es92x+uisnwhjA8TC8azlJWZTgdZa74L1SicqueFgPjXUZjTfSbp9pV2fP
fLiuPf5az0WXhFV8mEx8ABonjPQ12D577M/vmHmdB0pnZ17bHbuddKwFs2I3tCnXaGv+fxHaYvIH
7SqmxxUPupGY6nQo7MvpT5OD+q09TN9yEH51r9CN0GB7iB2iOmiumeyYtd/nazRVSaHp17wrRT81
GP1FTwGq8yvXx6lKPnH8HKXIbhwLPPJspzsQxVEh7VYMU3BE/SE9U4PsU8ZQOH6KjIZPvp057BAv
jnexyMyw8LrsI3wD9ONpVreEa0yAoRNnB7vkxZRoarHChcy//xaAd5/H2RmC8LtOSYp5ACsbJ1yL
AroCMZMP+4WYYFbiCWY1lHOspYjmimqH9DpnpXipwnpIfJ0j/k1RXkyP25Jp5kUJsrmjfGBCW3X2
eOZRWKLCe/HuMDjaGhUfTu16HSCkhiqW3N9FbuRzjwMjRWeu93j962cnwJJe77RKvSy+lx9BTDcI
Ch/s6FJxNv36Qw2jSn1BVYIPBjmq81vjzI9+EQBOzrAQj84W/f1Czlntt0oQ3ndOYfR7hqceZ5ML
ZmFbnEKUmg0lFwsxjBDNNv38bxPVSfxvKkDTVZ9bTT2+c4IZe+f4w7vjHwhGBnEVJmRJC3ZNwQ99
iOWMLH1fmFz6KE6izaHbNXfVPCKT6tgybWAyJ34NuFlwdX1MCqOc1PLSS47rIpaao4BvCbejeBbl
Fzs3d7E4o6dfjAXjY+axCZ1h+wJLb24jQK82XolslPlasVkNHD65oNm5l+1Qp0+CwWU4UUS11Sdt
e3X+WCRFRvLPx4Ku+LpRHS7k7OF1/QMTDkLhBWkn8gsFd0EzqEbwNuGJbfjV9u2ETkEjdnvqS31q
KoCut5XGWLuJuBygaBhMdetgsLYIlZskPUFu1Cy6bfvwBAEMX7gZp4ZpQnBDXlU/A0xZBaB/OSZ4
O6goGNRHRzaSFeV6UKSea1BJzPRN4hGrSXJ27wArbtXP3Tgg3wx58jzE/3Q1URVIWWH0GfoBET8b
pLI7AIiQBZNC62jyO+uuut/QpZQv3d1KUGgk/wgeVf1oHovgwnC2xWAabaVzrMhXOa/HSjWna3mx
cO5lHuToXze2RH3bNoLLAaHtbHruGaD0sElNC5UFIHAtjSa1DKe9aC62dEkkhldjgSujmvBt7ROr
DIl9SlExMrpjcEmz+FBXDAO6x74Za3m80gdPdTkThcaveizZsP3SKdCCIQNA/bub6SE52QvrfWsT
WnL2Bvgwd5mw74k/2oayZ5x81MmsjZKIGb3xQ5F2xoKXrIWGPCP/ufV1zy3JlTxwuKZPVyitRMtt
ZALQgk6/tocAV6LsWcstWIkCjYoHDxBwk1UDkFkbSbE4cYVr/2kR9u16bwcN5KIDFuaINgEHLlPU
pqVXxEZGD/uf3t6+G2/EOGAo6CWj3i4ISZeG3HSpQwJBHMCZ6exOsbbsZLdMCHrCqsuACfEM3Ln2
rCaPuz/P4KvY46sfVfImzGejZy6cS646KnSzAdDRMGY2w7CWI87PUZJ/0jF/AnXtexEV7jUbKcPe
5g9UkjeEnSGdYHFxqgIH2C/YVn/9mnYNkAiHaXW9K7xbCbVh98L47UB5BNz1jPNGm+NVdoo7eszF
WXiR7MjqLRG1grZa2Cug41eZ8D+N81agKF8jIn0QcyuYwgudqPXlrk8I2rU1JpIzN4NpY9Cgn4RC
/0R3Xu62rE/a2wqTmaMgniW0BMnfFmmpEj5gbeD62bldfEWjX37nHDgqoX8ZmrZTWJskZe4LZNZQ
on3Hhv5q/5rs1u8iiqYtm9QfeWt4aVj/fv8TM2e/LtB2TaE1R48Gbd/sCcy7sNGdlTIX6TrA3EGz
F4dZFM722bqqKr0KPSxJ4zIrzPCw9f0/RV7hvQaOsd2KAsyd3V3GuO94/s08wHmMFea5CgAczZJL
m0lkEoWV8uL5qvwIER2sSOQy4c6j0ak+wZEcQjppxuXIOWmrc9/73/D5TjBx3Srkh0BhfusLw7AG
RCe3HFmsbIsx3LJEwXc+dUf0EWIpK/seQ0V+KDwSPZNUkoNVTY9YeWnm56gm8kpngUzjM+h+L+PB
dFgxoMD7lHnkHegZ1189M++abrvMrlaQy5W9w10SZMxEb19bHrNRrFtL0aXSvVaYFCS1saRggosl
h8D4LCaob/YXblWA182yT8z5oQb13h88pqKR+p6Dhh2loKLBdXaG/7zYLlHjz3sNXg68c6UREZPi
SWccIZ3z61z1fyjnAYfEqsQiILjQubxXs2b47vxoqm/qje1//OFHQIIOrCZH0IXG8Y9P6VjS5X6G
sY6hCIkJa5YlHoumMpfkCVum83X6vwhZCOCqU3Re5tC50cSzhYTVqM8z1GeVF0vIVvom3gPKa5I2
Emi/suHH5xH8+h6Zbb9WvyG0P5/bVKal3wO7hxjUMceV1A4g9fhpCRPNiGJOhnVhHQegWKpbTZci
/gYmncmbRTqejDEsCBDZw3E9xoPVtEK0ELu3GJCbwmRcdPPc+F3YvwHr4EuoMnsPyPoADGbQyot5
xn295Ga0x4t2eJPhqfjtVS4dc0hDD51xt8k9oBMI3ZRI67r3ca5rRgr0apbyLeqby7dVSOvND+dy
lMOkjwaxzS2yBU56sUJ31WsIGCS62Dg+YuLwBaYTLheO21m8QJjopW08+49E7mom4Jup/TjZuUb8
NzUQEi5R0AYRIMuRs7swel3qE5yUlpgOGdkzV1vCrl9B0wMiTBO39LzWyVitb1UKLA0qj7QSiEOI
HBX8Dy9a9bRJmlcglVXmqfbeQAYco7u5f+fuvw+EDtlocfR4FyDEGdQGWHHcYQlF6CDu+QYledaX
ja0CctAHh9G8rfn4N4aioPXA8D3mzNtIwngERGq/Bftk55Fgj2g1+8Q7yZp/R8CoWkI0iczLz06c
4KW4wBSsK76hSY7fikktdrQQnqaXNtg69lpKuAdPJnHlY/WNdEVy9TNh/senbQSfT92agAG8rJb9
QE4uRIHaaTlvjzwwBbq+2kF14SV8Yoxa8grfhm7QEUuOG1O6XA9boZSI52aDUe0fxX6Qx9BCyzsC
El96lI0T8iarDp14uxM2PFXFvSnjYkoL91jVCD8IylpP+/qg6lgKB2mw6qwcsovCrqQfPC9syplx
9PsbJvvDUNDv3D/2muaT10Un24wxk8iyDyDyQSD221e4C4fUXg288zVEyBnZhk0v1qPTf6poOXw7
Zur6umLG1+ezqOZjEAQDdsEuV9M57rCqVi5BPKqcvu7KLX+pix6GTUqMAZClE8a63z+hSCX6FB0Q
oQCFEeUhYRc3jHZCTkO/S6Ifo1WfJ3nOzqZ1Zj+keXyxp/9fQgQ7ardgeR4ngnDg/ZgQtc6I+N9c
LsDn3xQbkXgPEdg/wVQs24p9qSXNfoNY9S9K+Qla3llKgzZNXANupC63SxI0C3zh5CPHYdKood9V
7meoo1t+8+WBsqSy/4sJWrRaoOQ5sIxAM2F8EPYI2g2C1YvdS1Tb2sTbDVUoOXX2UllhL1goQVxh
8JhY+e16Gc9Y8S+qqwvGY6d9ZDjyFMvKX3xfQ2QVbFdyVaHm6mzdWwZeyYKNE8/1BjDioMmuY+K4
wDiOaTCXj8qwS4WKYCGkX4R6ZwXyrEUjngVtbOxUftok5+5+fujeDiXzaiGqg3eSL3ZYnkwLJ8v9
sjHolGsKiKDiRwG+0Ym65z/A2JPoFL0HU9v2hohnk3Dof8UbtgxSB2xBMCeoAO/H9L4IqDls2wHS
6um0mwLe36jX9PRQLgpw2FRvmHN9wUWPm5gw3xMNVybr7uXvLoPik4mTETcZ411DyXGASDu6wgW4
slrx2/z/NMAVeq46xXTGZikO1ad6nb2HkbXHKk5jWmNi2U58BLMtGmsqEWoe47CPT5LOsyMIt6Z/
SEi3UmCd6qTIbS9AHmyyyvSmg4O/b4aNCIyNhDLxbEpzS4U1AE21DXVgmE18H0dn4ukl9Vtjj1Jn
y30/AS3mag5o1VliHnafIR0xc5FZ1NZRbMkRhgH4VFovd1ED5885EfefECNJGA8zEUaQ2lgNL6cN
itomF5AKoXgbXKcmiG46VI8S3MbSlo5sYcobc1Wx6xYV/Dk6UrotTe1WDNS+rKygZe47GRHamEac
lGdqfCbMajCIIsLpyg+XNfhsPkoSHbG3ohjqsnNsgvlOuUDFt1TBYPIj1BtEilwLP2z2thN7tqOx
1Ny23vAeZrxskyhg4fKH18QeXDYlzcuzGdTX0SGUGYD0n6qiMAVP+pk1dX+fg6HjVxL51aLpyyHx
Wvm/jkfMmIWojc/VkdMs8B9a9SzoYbtXINQn2duCN0TWmB4jnV0B8VDbHLcFRRipXc3GJ9M8Y1hN
iNZRyqUf3jCjIRT3LzhShRpGvOjF6LE3eojmmy9Azo3fA4Gsr5xYyqgzFWhZg+LjMhYDjDKNjlJT
yOmLJex5E0UafAFXGsTg9X5fMovbpoz5sA+IGugP3k0zu6os7EOK2Dut9ukPQozp/PsiOJJKea3x
Rx5R6HWFsBuXrUM10rPN6501kR4ixWD19flPhp6go3nnyUJZkoknXPvwJiKHuaBLA9EQBbzrOorY
ZBUwDpBWnCqecVKSX+qRPLdaYp+NDhXObDaAs/H4agYvzYRitHrg0QBrQZNglrQGcsPVRnIc3E25
YoMkzWYCb96McGJ8XYv/fAxQ8WatV36qdKbHlG5pmzrQSJY+qHRJLSomLu+CNGppuPRI3z3pi9Jn
9y+0SrhsJ2yFmRuh3sAvgJCA0nX+3yiJ1ykkXnCBTF52hn2t6/qqEhtdo2gHYpPJEycvhCgcBzj0
GxLQ3oYnIYyiy4IErgYLAmi5U41KCA51tnMrPIvS8VT2PNHIvhZcG27AE6nTIeKyhsQL1qoqRVPh
ZbXcrBmis3KLWOtcSfcmeEc4ArXd6CvGOyeROHMxiPe3v+LWtfquaJ4/6uImrOsZ+EzNjsgqXcr+
QEh1+NpmL45qcM1jQL5V7GaAkisvlqegVaa//voKlHtBXp63KQQ3aIYySIUgqB1mu/j1BVVpFKXW
pUpySopjqMPBJ+Kg0hspu7eg3DIb0o2O71DXhBOrZSmY4ITLnyaxEfkjzR8rj+eCSmVgczCyCEXI
dZKocjK8G+TMhXbDCG9YPEoj1sQQcJyHHiY3hxdqZ0R3Hw+gMFBwsTcfDlqbdeAPQoPC2lvySY6M
R1X3U1s+61UxssreKDjdzS4KV5zNS8pw98SD1UIxKnaO8mU25vEYJrC+Q9w9Zm1S9A+GhQ7QaU2G
J8Sk9Bz4m3I/3K+nW14pOVa01Z/fYLPHBbex6ZW5TcprEW1a/AH+JSm4etHWfLHQko2ONZtRxD84
LlWWTMiLtjl2ioTP7HyXXiT5qsexJ3Rjvr1TNh08XFPsAgrxzv/E/65bH2RBvr0l4iMQOxvBXPa1
nyfu4lOnkXOxXCnqlwyd1MGa+VANnCv6n8lZPCS5QY6zi4mD92+qoGWTavd77qjUgRJoR9ScbURf
7irs8Kdvc4Ai31MWFrHWNNLApGN4+RrQ8Cwxva/G9jKc9YHyhakGFPyWQetXWqdcIv0EdYzhekyn
6l9KytdVGhLWwJfpU4DU5+qa8PFX46jEssM/XaaPSB0fwH0dTBGFd2aafqrviPUw4hzKdIk2rCCH
ofPvxjCuHLk65GlQE7PtqwbkOFdegicXgry6LGh6+nueDDKUe5JXRDgvrH0l94JMFsgivGkHhbqZ
3B869y+eZw47rgI+LRoMb5M4ghz1wBeyPLrNuM7rM8JaUl1sgmfuWvxzoQU11+yMQBcXICrwpi8e
EggT1/e2SEAnxFAe64P9QYsWAqaZMeGbureK480WXuqobaLVNUhMtcnGP/7yVNQAgKC6AbTneURa
Ws5jCto8tR6dRhYkKy0DamaDJugj9Nyaz56f36lt+2KRqWjLDgxxSkSqbZSot4or9Klq5IJXrGAv
oMdSSPfzaPZygVn56jzGKH+TNkOkhRlhI83o9FmyU/uRQNh097BeNdZ2IZgmJQ8ZqcZJfOgskbmp
fLz4L9KsSUjn2IpeqCTNbw0rGnT9/7sx+N2O8F3SYxva4SqUOYwne0KW17XhJdEAxwyTp8Msddjr
ZtOajJgqMr+Q79V97Jv03pu9S1q9wytVqnZhexXqWPKtaIRwyZrFxLHl0ArZa9JxylEpYCYPGMpH
MQ5ouxZbj/Z8fOn+Iu4A/fu2QxbIxU8IHtzs1ImzhzPvU2bXCwR8TbJiqbQmCZqkFyEw9Kn5R0u/
0ekzAvLEmh1r/7aSlPQlmHkWIMknWWGxF0evtH4Qo39leGtgRl49F/s3a/mfEWPAcc0cSPenQRgp
uX1A9C4cIuMrBqESNfrbF3Enw6m8CHTFYUqq640YFPO0ZdOK8m62TRNWIa1kLTEbrY4IgUEOT7HX
bzLgdxVQIzY4rebQDmL35lN5duNXeqh3680QJ0stOFGCPEWeBBAz+C1upMsok2zMPH+3mIsU2FVb
0azi4AnHSt+2zSuCmH+v1JKxmsBvjR0fsfbB/JGtzhpjN10dRkEp8+yu5aAnzHVG8pk7VQ9lIPFy
AVArs0/UbtfSXZe76VqGlZoK+J3KLAs4c6OjgpJWLJ6bonNxNokuvd/0eXFdw6giG8DsyG3hnfB5
UQB1gbmAnarVRQp4yUE5QOYY8DZh/FiW+dlZD8ikmGl0jsZ79EnFyCld+XE+H13N6DWjFD4uMZvq
/H5BdsrzBnnfExQCsPdBMJhH/vPrrlPzDcAXQwEf17Su0vGZjIBU8QCEoXMLzEdiEELUVQ+IqSH/
z6Iuz/tXy6F4/PiSnOTa0+ZMtGCGcChHpATCPx/xy2eFRGopH7RqHVGKzEx/xSE60H0mi0EC43lO
hEo1MS4PvANAqyXAgs8JsGR8CArVp3vG3YVvq1WPm7jBVaPTPuEuw7A381q4Zwu7lJHCcvVWLyVI
sInXd/dpe1thBQZTGq96aQqJw1L9Ywf71JO4/bX5pMdScAhQLgcAqwrrFL3NAc05u7xiu+T8mJ9n
Eiai8MDP4M3QT/np3Sa69exRR574o7Vu6Va3kNWcyqB0v1p3BHeO80XgCtCZfwLNhUmCiQRFFwxZ
W+2IFSBkdWhyrp8LfFSe5N37fajGQKLQBsy4Ajdmt5G84i7FMD+VJZzE2F4quH+A9FimSTTNjkgG
pKrwFR51NG5hQ/hhOxtlraEwNZG6KVXZCTny9cV2hEEv0FMj+r1Htvq1sp04b29Bmm4m01wTX4J2
mChUJimedtjez9gPeafzxYpSMi4yhC7bokCba9UX3X26UgpEHCaj6PMZGxk3WZLD0XA8DgDyrEd3
4BlaoRGJrEd4TF3226/EcJOhnKaAoh8sMquiWJNdMcWJssVloTEGA1xCjnRXT0c6S2/dWpxfI/t2
agQJPaUvhKOu8saU7hFqwmpOYjYeKZT8Z4oAy0RLpvWMsf2HVCaUFzR2CMxVntGyqfArHfYRfRs5
wpO/1TB3RLCeAny23tWh3KXYgeeAnSeqFGUSM1Vkc8vQPY75YT24h3gBqon55MvvKHBKKbpWT7w7
b+r+/l4q8mXbiTvobiPOuZUXKAlSO+wT5n7tW+VCkzmnYPKth+lS5vI5NxVCATslyneudwalC5lQ
Z6Kf+ISYOqwChldKiupyMPPH+mJpVMLaASdpjGf3cuYKBTwWriZwIwYm4iyN5BBEFUJZy5aYCg03
MMTxDbeuLrN/ctJeDs218EbsDEmL27EHeFFRGTNL8ibqzrbxdJZqhsVMfrks6tVNMJ7ptJpqk5LP
JcFaI5AEsYk+pvlnZ8SWGs9PJdWCQsQVvA/vOYUDoaWP40rCKbyDpe5aUvRruGVtp9tbJdfsyVBn
3pltlx8V9KMQbvrc+aSCZYf32hKEV/lBhgI2SIBoON4V5/XaT9D7NDtTowH+9YRLGZOmyPfj/TGZ
olFJaDe4y966Xanf+/QHh5EnUeErP8Szd3Xm9z/g0IgaOHihBVjO5MhfH162ou3Cq1wC7jKA0/Ef
QCOgvIkLan9twTJq5hHJx+/WxcBZxkhQWMC3ut6rYLt9w/Lm37aTu8KV7uQFuri7ZU2u5Q2aYPbv
dQPqLTAtMktqm33jdUlp/Gh7Jmb1RFzcfAIUh7cXHegzcCVIhZT2rAkeniUkX8AhAq43iIQfjUoW
it3wg0LjeBLDtkdVKAZcAfits50ohtftl63Qrhm3iPYs+i7SKtddpomCFnTJK21SoSdeuRcHkM3u
nikc4qaTgX7rrcvr4km11WsWvvD2/PlPpZZXx0TB/x2rAKRc9f6CCecH9jcw21hpvO5ProeoZRT7
oVQ46aopVpM30wYZw0dWggX+lqm3DOUU83tTkiQnNV1ZJzQNfEtw0m7oiF7xQmADA5I/A4zH5taW
UpMl1SBzDhJ2DSqChSDSUGahYmW4qzswGad+yQiXqoV8phUVIwgsJWvhOqmZs7qJGFABx+Cgx9sd
PeJXctULsDx0iEjk1jug0AeTAAEBoJIYDxa5pCpWC31wBxTzprSkQ+prqog8ZJLGN0nOWteqWdR+
PP4ZoVvu1AF8HFvzt9k+F/0OuuEHizG6z5NdhWgiGyc2oOziY3X7nxlmG1t2I4C3iS3spyVWox5U
xZ+6D8tkI6nIlrRN4lnMFGxWqDWDEDdmbeTql8OgEDCx0f0Xon9892Px4gIzaWW85+PbCDtqNqFS
dG3sLcteAMl97UduEj7Nn0JvjIGO34+WSRzsJVsqawnFBzYlTtFhnHtQ3sr3aAC8NGSVDIJJ3t3d
aaFMFeoudEWIUevBdjQwBcCrtyeQTI/VO+6VhpPXQOJz0VWC0KUWXcf5Q/5eLyC/rluvLY7avpQn
XCHLHJrfY6yy660buWNpH6OblYl1JwEOkav0nAdXwGvrpVJh10UxQRJbQeQ+jU1Plf7xUvQ45PdB
7mVQ0ltvRk+S0g8uwa5AYePdIw6gldbAQZWr9JM5JQvmE3RroQ2RmNo6SRevBIKjHP7AAwDJVnvN
pTZY1UQYS4E9EifW1qIasXJvZNIiBU9h3H2rbjZP3Iq0TvpjuJcvwsE8JtSwwp0+d1OM9ufB/1f2
AaZkGkJDsba2JzqGY+WzTzfGxGcHH3lwjxrikzmKWkJfmVcnUUbfZVekyNd6+8yWRP0qyjkFfOYg
rQmwnpiDQVlKWyq4nzTd5CHlBGOp7hO0olixdKJ9reUbneNTm6BsMqLCY0tkV7SS4s2Zlnus72WX
O6M36lr9mVWVVuyb5e+hcVHmtjazmzkn+mBlEe00sIpId/Asm/flLiGKVH+xQd6qf0lOC7eaUsAV
pyGyx0uTZBfZHQSzOg9LJOTtXqUw3KBtmeb78Wa1un0emSsd9oSIIMrO5VjY6flxkAIeCNFyF5tg
6zYenm9c12PQN9lC5fJQMvhcRivQugriLhvPkLYQEUMUq2B+nu/OMteGmsWEt98BaNom5YdxjqvW
JdSyS1X/ItiYTZ2U65Ep9wIytgbGi2gxVrAujNZ7sgZAfFZYsNQkKEhh/pyW2s4QXKPBkDgA7vIN
3gaiop3U5cr+KuTaoXeT8J+XzoTYaG+LvpCB+GeACd5w5+yr1bbr9e0nt/0a/4x2yvWZ2yzUnPNo
j9nxRo3FZxbJWPQZngPFdwbcHLD3yUOWzu2+Ur6tmlGM7kuQfl4mplaW9HY7aL5E7CRoCrFxUmtS
nyIFQen95GVJN9nVZxaFp7FPRu5UFM8XfE+LpBFPcch/q9ZHv86Ym5L+RIBywiujuqZFyxAoVAVM
xaKVPIXmlWmgpA0gfg9WVqleeFl7zAP87Ir5deLOwBUFeaswBUy98ZOnKGT5vTxa8mD+5Qc3xh9A
j+aD0qSbhZpAT+zk4FBP9jIPD8dbtyGowt08FxZAtAy/0Dd32SMm1Ws/J1kXZNWK9vByVC6bxNOS
cNbwqRytPENGtJ365iBjpAdTyhLm+0YYJ2dLllwntum31BuKpYXZ63Tk79ItaDZfAquUaCVJDQOP
3Qnf+kxu3KGnF7H2Q3GvceP2tePYfnTe4E9RvTryGfZGApBiGrHlxgxrf48ZBe6LTvSyjNWha6+h
c5G/mWAjUFp+cS8s2mtQEugP235bQcOyobQ1fh4Cel/kq93Ls/V22YnAa+EQk132hz7AFjuuSR2T
t5ht4Xn/J7ukPw0QqdSxRE/qRHLLXD57BXDXv1fzfrENzDjWf4xKYYa3epUUUC8xfPe4bHZOplqk
VpvL/CCnUBUBhBISUVYV0YeZKi/0lc1amqmeo7CXkezOzhygK5GfH3L2bni+ryjzxduXr6FqIHU9
kBoxHr2fTzR+eIZtYEXmaBtyaTN6CHDjDBaC2usO2846aVCs5NIXj6kgi8N1QoCkyf0nj8qxNPuq
gmid4n4ksCDSPJHNgyHPr/AsSUdghpl1Syn+pEUsmIeadO/Z3VoFQ0nDXIkHBy9qas/HQtWJnzCQ
ZY9qsJkBmXOAwBl0ZWJkOr+A8cq1eWBop5TPlbInA+B1a0cocz35nucvn8GVj2Xj/FnQDEMhUZA4
AHHWEUShMkrEXsYWh152mceXrGDn4elR7s/pARbLC5maJx0qSBRirEPgj+OAMiJUKBxu2dX5Lxag
knWrKpVaXCShxyvlT37/2gDxL/0U0D4acXEI8dCYQhdWDAp+1dC+E1YI6RCKNOAddnpF9GmSgH7Q
sdGpZ/vSm8CSyR8/4xDlDsvpeftS/xoH4IY0s96PUUsJnna05SosOrR5ysnY7muUz5M5y7Wqs6uq
4jkY0VAEh7Cdor/a7h1qV1FNLVEh7KDGeGGpEYb3u4oYmSFwyGJk4aFce4NSOY1fqw1nWeyhPHAv
kH3tl2HFlW0brd56QN2VpNvDd2a0TP3jZ6ZlPlSs81ihuYqyaC4WJke/smiVTvEYPw3FFy8SLk4k
6whUDr5bh8dLJevPPrQbvoqQg2cgyUeCjy75WBidnHIm8O8KuoyV+Ko8Z3hNz6+77muO+RhqtaIq
+s2Xyf2A7vlaZucYVOuxQoLCuBE/9Y0i3GUryUP3ezCZFSLyyRKn7yzsm1No3R4whvspyCqn4Qgw
dSk9aXejTRsa9zW0GOL67M8lC3S2HTTocPvkNbAKp+ZdZnCVyvghuWVK/1KkJddT6UD9/r7sh9tL
YdlchKxtNDtvIouWqYce+tsFvMve24mbkP9mcYG7kLBT+bitHt8im/ETZqPEDBzEpTVKXuBCi2kr
KwRgvkKbdt15fp0JjI7o1V4bvBxFI1zTomwXO0xR5wzr3NLEMOJ/dWgjA806cwDn49GB+IFVK5N5
ucpSoNnREGjE39SXE9djQr3JEEv79paAwolz4le6IMODeHE3/oncXwwRdQGY/lSe1XdXUprfEfcO
ThPqwjhSQFHu/z77P75P9TU/0+qECzsOk3orN6kU49Df7xMhb+7qoHoLofqzqoBsZfbM6k0jvdQ3
m7H+nIUC8wjqAB1o0N3cSw+lAWDtlkRRBQAa8IDOfEBOFrwlWnQAB/t14MoMHNCoGfTWZnHDIBoR
8/XgIq2xfksPFfkPeOCxJtt3EVGb7KTIxcZNJnuqjkbYB6G38jLrdRy95XU0DLp0TZ12Ba5EMG77
TT4OyoqKytgWbdaLMsFGsdySP4vsRpC2aMWnN1PmTMMhv9/ZLUHeaZPuO1IkSx8mvNUSdpl209RI
E9A+hESPQkWk0hqKLU0skB9mGq0zNRtOD24TlSB5Fz4VTM4kS7Jp6dVNHSmFkZZXPQJrXOFdAevs
AO+cyA7DZLcSy4FnJZbWFcLcYRh7q/G30Rmmgaf9Gju97yHX4mkUbkAs/g2HV4C9W15aw7vjplwZ
hN0jmwAxs8zrtCnYESrS09dmNmu7zCOeZwd2xbKybALersk6zxXr9mLYVdr55xCeWqg1EgEgAUEX
8/BwgMtoH4OrhqKYovQnJwfpcRi2KPiE7TiSU1uOLf0k95r/WgRalESy8ZTRNziuoo0B7833o8mA
wBEQJAdzMVRTgwNa8Q7DvQXYoo2a0d6n6a6VtLr89Lqg7uveQi1F692L32aiol0gsTgAqNyakb/Z
Fb4nvaN8VjxvPZ5bPg68THPfuFPwYO9w+JS03ydBF1mReJ4ErEtqg48WzExS4thU8sf0K7zS7M+p
KpqrOrCLzmNQ+0Luuq7lXR2jGsPa6ATbaxp3Smhf7SDZ+VXrkoOkQmPcaP7Yaslv+JA2Tx4s+jWQ
za40p28dR3vEVhEhs7Yo+90XXIM3cpm1UBYyFaD7+//bJ+4tzjLsfR5+qkRfSDT5WRg8NzLemgzB
waa+i30SLStplftUm0devLQ1VGekK3A4JMIpFTkI7+fyu1BEpDPkwqvec4ABD+Oq7yiA6LFFfpDQ
F3Us141e8kRh1hffew+eYts8q8nih18Sl+AVAgm9UeVEpMO1cbelsXs0ZmQhSHpC14KHrLmSYixB
FT1eSxXZ5tnN2J4DmTZjwVQkF3wPw/0qPQTlGZBFBP7ni4IzXCX5JFryofvYXYjjXsdUG23waZn1
vyiQHgF9EeQQCLFD+vt8DvQr17zPZ8Vcou1cKBHMrxi9Yu8W53cnI84JMPivejhrj0ic6oVU6Sol
5jWv6O/SH+CkJL4A4odUlBxS443IwzAZz0faFxphwQnyfg3oYXrGh+r+0PCJfY4qq3D8LNf4xLLO
I1X+GRCpFEc4mAKZI2K9IERer8n+AftcLo2Z4YNza3/zEWfu90hXBzXDX82JXXJIFe7zVlfsJ+QK
/Q//pBE4DTAi62qXk/8fZCUKMAIGgOYe3KwZyDY6GBpx2lmz8L904KHVnWzpWNVZWHNU7xRgddyT
dVjzdcBo+KWj2TLM9GyKy+FDoSdIt5sUxkc3I5Mut25RXfESf1tBZPsT9F+22VI2Dm2ar651Xivk
QyXxAv3ndCrvFJaoX9BaFkCYhJWcYIIdFdj2Ix6zco5cEMv1jc+uTEpvDtGNMoqjBaDwZfzKw9aq
mHcZPjGTgtbSd/MiRa3hgKj8ZHgd6PKnJfchCat6W0A+M/fIdxCW1FkDBABHCm7wdx+dL/6us0HW
hiGTJP5AcP8G/L4FAJAuGGQiKbC9Yszkqk8+gfOSbp7gWHW4E5uh35PcN2CdmxMSqYyH6P+sw8ju
KjVi+VTnu8h/t9out0ynxHBu6sTifIPJdCdDAWibWrRnC68Eyr2gGbHnGficIvHWD96+Mq+mtp9q
7/sQNlD6SzKb28Ete3ahZBA6oWmhFFVSubYz3RKx0gVMGoqSzqYq/Gh56Ckbb0YkjkF6K3On/tfN
vyIPLAUEcNVY8cX/W68s6EEeN1/gOFK1QEStImYzbqFjwCNcAgMR7cbLl5zIEeXctS34KU3d4z7B
W0ATl3tx5Ev2jsS8b9EpjNM9nHDdtdCYvnQzgcJedGNmg0j+YgputX3m3kJHhaJPhgwImt1Cb/Ko
4jatRHIGZNvfUl39CWKJoj93Ccg2ZYeFFZPXmvIVg0VohU7JaZIEWT4Yw/9+l9mzy/KwqWWReq9k
Y3/lmLEmS20GbZkt5hVX/hrFgdDGvX/8m2OXrgGgyqrIhK02qcS1TxTqIO6HIBp8w/wtg7lm5Kag
/Cl7SFM0wFRK+Ls/SDGgqmgChgQu95ChgNpzJViWnjK1BB+SxvdRn/ydwgq4ZBm60pPiEsGuF0SD
b7vkIjIWVMqRpI/fpgqvMdmp3cIgzvMqa7rG2Sw3LwHvSc3fePSMqRl3RQWDLgDCbkWoNd6OEbij
RnmcJ3sQ6Vtfbx0DUcRd7TK0UJjpp5vAsQkOxWyarC7by1j+1zw63sJ8lqEkGpIbyypvt/XzMXOf
4FRRn7gNGCTL+GoZPNgyDoQyTyMFcY4xcDf0yqf60hNFdzxyCH3GgZWiZTXTFp1ed1C0sVKBHw6q
fNe26hOs+ZVn27Q7y8IEuOqHMfsjIp0U0wrF3EV40ln+BzDsrQQxewr0BoNTWjwJXp0AlPqDUcgZ
TfKduIzE13wQYFYOk+TJq+GN+1rpcN+d3yKpFxTY/p/t2bEDgQhKqgQKdwg5hoeAS01a5yl4rhBl
cM55EV6N7uNSY+Ds9UfJeBv4ffM8E7vbf/Hmn2lncXT6M4RQBu7N+0dpIChQR4wIOVP9NiHOKLr1
jaoWLtrO/62DTRuxLQuGyC5kbSsjFamNowI0bdXRis5tjU8SWfd9Ec5L3i/oWkR421JaV2759JhX
m2RjMfoGd4yeXO1D1/zXVwNqlSGADK6J3pI+NFC3vc0zweeM/JiKYFqJUSnunFJ6Uqmdcd0tzPOO
q4zcLvM8iGKQdqxvLL+WuDdsqoJvH4A/vAr1Ilb50PIP0B6QBi9nI7SelE6ES8FOoq36zBSdadTe
a2tsUOpoTgOJafMUqNfuq6mZDJ196/HhleSaFPUa+pNWaYU7t3WlCUElx77CRuYZCgGUXATiFarg
tJdRasdsRXkLtALjU/RW11hgjy4pHDivpkA/qdbauc1Mx5M9qxcuRVT1KoUMfTTekcNKTtLT8Y/T
5VMSUlgl7xNdOhgcQU7EznYDCQSg8XeD/6kDDNd0slc2dMfdEarNJRm5GuruYnU3acqbMvLj8v+S
im2YpX61X91lAR+qIzVeQwohf+fzLXbQ6M5pxeWeP8N9ZokUKFXTR+PHVPPpi+qWvD3BXPQqBiNm
Ur82JoLtlvHtq69QlEduw5CYgLLg/0No5REKecXII/RtgmFrbuygEjB3xaZUElYqHlNOi43pGFrW
R3lvufFKUJcwjyUkJ586FWJzJ/wkset52A1jGAR2lwIjxYpG1DtQXdrVnt5oapUqOVpzgKrahsEI
g8tboRz/mHRcqOJedUeEel76Jg+FS30ffGkI8T626ycHPIKqUYBbPxV3WTlA+tByEowWlCUCPSUo
mCUZUEPaVmtxiFtwVCdiH163xyoqWyoDAcIVzqsZbW1rK+TPf/8zqsaYIafCn7Y/JDxwaG18i01i
kyMrieQ+dHyNhaHJ+YTXBhOWPvVR1GEZmQAyMwmocoaBQwS7MZTDf4NPsx8+3KGUXL+P9WQozYWr
1J+0O9JfAUikvimDIWCNVsGMHstN8Cbc++8t2VXHOe7qmj91IyCyRl4EvYQC/p/wwGo1g1hA60MH
PYor4TKTiWXsswsIL9IORG8rOVf0Xk4+hWpIOTeSctrPTmQ0uhDaqES03M9Tuv/nnYH/uAY/6Kg0
YCMWh5bP7bNewJQOnIQUn4wx4ylqhpXex0/S+Kblu8psNTci7HpWuDV65yFIQzp8jwwo5aiyYFrl
pw9VIwKFPrdWTSiDN1F7MNLJku1K4Cwty7t4jeINqkbTh3uNnwCaMOFxKnoqj4/5T6gVqH0Qq2UV
oENCisYYYzTM4C/l8lCRXJYd+Iqg2IHFyje7j+vj3jogmiMrKkQ2nftZNeCiJHCNde2AQvziPvaZ
WdnK37QaV+MND+JAnlUgtXzve9d1I/EIq9NbA+mFYa+4yuMGhQctecyiaKcex/mffMQCKDz7u5p5
/VOQQQgsHtQ+5GqyhbYvKNxG4YD0b9+c77jLCNBOLKKeBU4lFBBCawTnnnOdmM7xx1krblMbqGkf
1QNTSVYYoAV8N1BY8jRqu9lnSo8rXmAOtQiXuRl7ApAz5/SxnyMMOz7rXkBRzQOknr07wE/LMPFd
/LHMopaGPB4d1Q55n4e0zEMtBOhZHofjgpJcE7w0hOTRI8k0xbBkN47dPPQcDlVeYBQwSlHtgvvN
JiOCemTAUgomcJn0/a7VfU9/QUQ9vrzTMkUNi3WbKUunVDg1aFp7HxbaBOed7nj4dEmaR5oyxAxf
C+TDnwge8dgq3TPaV7itIiqMOcG4XllV/2Dz9GxSIAsnHolg3Ova88RatFA6EMdrxGw8LPpndH5w
+Qn2V4hDOEGjY7cfmSPv8EyBwWcyW69QpA5MQYOyQtW7eZ5Zm2NbfDoDXa9YzSunqx3hMZrjSHeQ
9UDe4Z8Qsh4n47oEN0QNRRwzeUn07LwQFIOB59eP7C3+E5kCw/bDIS5Z2FWz1tKe9fZOEJLMxERh
PIcLsXhG7qwgo6kv1IwImuysAD9Lt1EsCBvf8EU+vyED+afoZYSUCDHnCGbZxABGbF85i6QZYU2L
AOpXQLIy1uQEr4Yk7I0Q5WmRZnAomHnVBQMaxMz2fvZm//Xyko24wdfj3h2HXO1M/NFl42a/OOig
Ye/vhv/UkA0IIPaJzwJLO1jK2KkGGY8kMocxWW0VBzj9UgULclIzZcERafE3NDi8cJN/0BQ6a41y
gXIh4klSuKA6Oy/GbKaN8TXRDcQXmNUKbqi6HjUqpfdm+BHqyaqfIMqB7THO6oNANdI7f9a1nl5K
Gg41sb4WJNNmzmnRnn3vnKsOYMIpF30We/6hDqMehTBlJfncyAi1OTQKaH9D1JXkcriH/QFg67dU
V9yiXgMR3HKbR5HLV6ouosSO4hJDFRljyvCRoPIG5gZAuh+XjqzDsyf9xOS3mYYGsforUKyA5TtM
usCrLayFZuzsjNaZH5PreC+SuxbwsnryQUWsW9CJCE9c5R4WjkO1zV0SClkBkbRxJG77W8J4+oGP
NytO8Cjaqg8keCYRqNQrRuUdFydaHEd1AZ0/0uNGewQIc3tVP8vSKbtEXWmyJY1JI5Y2kZmJZM2P
j526+zeM6DVD+MlnjMJBA5OHd1xJ694DT5KzYH4OVy62Adoq5G8wmwMhMFU0koE6LC6O98PLMR1u
8dVvBikSdC5T9i/9kQa1MrMdmtZr8S235K0v/pNheHN+Ib7b1b29WoNlHoKKRZqwkxC4jCDsymT7
QkzSWs3gcJNKbTBURjnfqcZ5UIiXsURmyY0J/eGuVbFyylkodSrJsp9Q64WTrdJV1Pm1cA5MaC7g
uluv7HGKNZUayerTLpQK1Iv7tL48KyIujMNn3xe2mPISqNraCnxr4b1i808x6aUkfoaA6psBX92X
0lPHtfoiskBOLnyceW9P3KhSZU+cbqt9g2pmf3MBMUEIhR4H3NCEgUeUwzzLhcOa75OdmFqO1vV0
z+gYpItKWoleZhe3SuPCgSTCqfKk/PCORES5QoXPqYqxPLx3r58OXLXV2Xkgt1EVjDrz8jCLLT20
p5Q/n/5r5ygySIVs3yCdmrSela+HviMdkhhpr/C7JZg+7nTG+FRzTzggysAAB40664h+ikdeNyhu
nrI4Fn4HXw9o8fEZwT10siAA+UcRGJAHkP+ht8v0s0nlEr25lzKNd0F3es/cJmpTXKPq4pP5dVc0
AsCD/KmjBMLyZfwV1hwQ+CPBudPx7Tm8DVUayhM18wVlu8vYtBfI+QFanUiJ788gZsyMxdSiUki/
HKWjY0b6VhtHexauBPRzDOaI9Rbjxy0aY9ZfYZC/wK79oTzPK/Fb3bVKpx0yZBKIeWS/3Chd9ts6
sFNwMgre64ncTrxtR9oyJQeg4Yv2Z9zGG9NMYaI21hrOJaBjXsFPQIJp8a04B1TGmXNK62jNlhuk
SV3OG3UF+whsV+81QgjbRbzocT82XJs9wpDjQB1gE9FjvoqAmlXpmNis3baxQeg1bV4acb3RfOPF
fecCq/va5xsP0JibNKTO8Ux78Ap3Mp/0+8EbmJROg+OHENa6gbW6R2UA7jplGH6iLk9HuZY6Idiu
/vTRBkSsydsQ29ROKS6S9KYEeKYue296cdYm4TsHp1Q5Iwjf5jcsltmfaH9FZs1UAI3YITWP7WME
RSimcekMaW+ZEqhpGyw0hJfb9uB1S6bMVQoRukinj+lIAr4lj+uV223Jc7/pLV1sRjFnZfmPU3fQ
YQ8XvfmKk2k9RXKNCv70Z5j2v+qM7n8Y0yfwaK4rdZZzdjFCjQOuth8OQFowEmMu/RJinFeYFqvK
Q2F20R+PTLmLjsF83JpK99fUiTYo0KCiT7JFToJxT0VwLksBsf22uBDHIfZqYDQeV9zRZ4OzPIWW
81m2l1FWzPqHYQhYID3mH52DouejVkB2me7gblQwTndIzAydkKjsH/M0v56XiA4bBd8EfCmrwq5i
obrce9MBqu2iSKwiHQLDXH15ctTJ5r37eoG9erLCRH82sWMmyFr5VJ9YAO0ww82+5pavqa//gVIl
7zQ5gz/M1UZUQBwhBayz4KnW3Imnr2pKUajqPeajUDlRFJ9wLWC44jeZzF67mWTu7v4KKQpe84Mw
X4QTlrsJjVfgUUZM8/Pz+VoWDm7uMX/iAoH1bSBqmk6Yn2ZlE+CoWUIUADtFh2dqYIba544y+vrC
ivWXCxTp9NrbmqXVpv7IADBfZ+cYkiw87GqXxFjikZi88L6YcZuvMcZCKEWIAqkZFfoY0ys9P2d7
Deefnb5XkZJOSosdBOsFPlRfAhKkiL5FVTyDHYuEG6iLC/i0Npr2MrQFSjo4AYXfxHoP75E6L6LE
lyVZaGkUw1BIsCYd8gnL3y9B7AKyiX5RBY5TsCATsTCv6FbFmj6stpICYo3VTtKUbBrQv/6pO6NH
iQLZkddWOF5MjqkeCUTPTf4zTTsb8uizBDiePoganVTiFh2CTs4EE+tTvB8p3VdOxwoKxfnpI3uB
g6dKhk0Gbkpn410V0NVBPcAz07VjsLMaVGjNv3jaqrVs620Bm/7TU5C/5XY8Hg9WsWvROHRJBH7I
7hgVrDAR/2Dr3SPl5GfC7eOwusSvsq3Cbz05IXHmxrbeL7ZVg9hqPHO9a/UhKpAFB2vejSZk/8kd
DiA/RuDzHzKUkyv6WYkUKrzVeFHYEcTWCLYA2gAFNfZvq1EnlNwksKh+nbtMq1AEehgvA6jEUIn5
EZNEAL5AYtDEvJwblYltogOZMxvie2tHfOxHBK7Vk9Uhl8WHdgZzJM9p5gnEFoFwphRNfC9rngph
HmN6fSP81aHyao7sOWkQ5tO8N47JDZ6bnrw0Gt8l+gP5LE0qsuaHDyGHuCdqJox7O/91AIojZmYR
ZZW68Zs7EIZh6KkRwcvMLWf4nTqvSu7oaLg44SIvDmvZ+Qu0yduj+c2esuKfX+3DmTX60uJNAEg2
xAy0YyQIuOottYsAam73G4bGBNVjaHpkqO8ohvUNnbg3yNcI1FTznluvHcAXN4zY7Q5u5loRbFv6
rtqM9AClzA6amok6p9t6iGh31XZv0HF749WcjJ26pKCiyg+2nOKiUQn8sVf3y71KeQ3DlfENa3wv
FRuRgNfsw+GERFxLz84B0orRJRCfXRXgR6uFUu4rx5X3Rnwfsbhxj/tn9Hdz2XkXkQ4JTKJLrkc2
LQmLXWYKvWoJbuMi9Omb2rWL8ELus++OqTCFlT/c+RkpcTYmNfho4KegGSNwLb2jlfaitojmJyTj
MVvLGqjgcdNdTWwnGKO19u+lTf0eYyuGU1Ssa/7rZ0VyPIBdpH+RRIfE+n6vrGt26Dr7sUjSigy5
8gnWBbKmT17ucOKOa5Oj3EfE8RCXVZUEVOzau6qwWaT7YCPJJ9GS/1WmsVCcXLTde/zqo72atE1k
4tiqoJ9t4YbBU4b4KfV6VJDY56dihvv8PecpesYit6pc75J2Gz8wkUqr7mxhMImKz2YA4hF0fmky
m1zmKcwa2G3idRLrkqH/FQglaCoACev65VMHDEafcsSSXCf+mO3tiOXRG5g5vdYUUWI3NYq03hUm
O5kHRGz/xB2LjIJZ0zsDekwMhPw1NF+1/pn7+W3LzogHijVYy/3o8lPYEEqVGArEoTx5qDK4JWzc
iQkiKGVvDN4qtHzpQ+flbVh0L8jIB4tzTpTDhjpC3I4rZV5z0gl+XX8oJcIDOsZAUFaEJyHaLae9
yNde9LmHA5OLFeUOIX9To4Y6SvHOqlKh7GqFHCblbkyVOd6crWSnqwhUYDLMWRXGrAW8Wd84/Zr6
pvSPS/SCyjpigzaFPizBlpCzHfbuzcZxjti070/xeh1Nof/YVo9HKq8shRLFb2rjMHtTpzlfB1jK
dvQlQsA4N0AfX7TpCTFvGaBQgmxTNfl55A4FkGj+tC+TCVHZogPzER367WlwhbF+WmIL9/vzFq7U
Urn+tYqv09jv1fwZibj4WMYjgQDwfbGlVnpevZsIpWLQBxQbKLbSRsxk5QdMJjpmwRzbnwmQZiCu
Tjc4r5G4yqHY1o4FyCVRmaAItsF5+FuwFmBCVOwhPo2MAss7r46eWQnbTx7A2QTtPItvkFwz8NSD
XPj0fIiuXTUyC+ifZa0WjcitrhEFxIEaPcVjVjR7OUXdbSlE/ivIYuyTFVcYxNYn07ARqDVWq5nI
olukfr86BKqKSnfjS/NOK54GXX+n4zXw+sgHPNu64WyL5VdcW2686zbWaWa8RjOC2XxlX6/kh9J5
eZhuKTlsiMfnsKdEreaZVbflDrACrDe6hK7bOisqCz3Tq5297svHD4sYtA/NGpC7STdUKG+klKCH
iKOVuavF1GGGDqAN1rpLXaOvGeiZt7jK4mLdEtX7vmtG8GxIJAZp8GTpm8OX+voUob4RoLXfKeox
I3Uheto+HWkqBQjHaq6FJmtsAxioZ8lRI5Q5e5olMSDWcdOdZ7fHtVFADwg7AqRsfdmVALi5a3nF
gSD/6BlAJ6jkfFJBFaSgIQ0PzBN7p67K52tQ0NvXAlcX8nA99ViM5JfNf469Q0s4qkE4PRWiCOTf
78NolyRqJUMvhlh2l+CHtoxYQO32hJwA1osk1u9rUF8Kl3j6ZOTVujj6AUBI0ngcEBffNhGhJtfs
Kv9c/xtyay6CEYKMkowNCrIXx4HFRmFuse+3mkgaovv9gBab71ni0f32EotsP5490xFuA2r4mFKb
vyp86nbqcqXfcIaCqdIwYjSdM/izj1bx9sr+8b03DeYkG5nYTiwy6UizMzVD8NUMMUPHRHSKh0kl
HPePaUEaO7oDYh+rGRQ4Y1OUpWrYXbGQLy6dWGlhGsjC5MScXfUjfhv7BXi0cAvq0VHppo3/t5pu
lvJJTQ325EBW//7xUH95pMwCKZp7rq0fQ9zBjWwUVagL8NJINXlD9IRBFiOylYs8g41y5IpyV92P
Ew5Wn8Bu6cEvRST9GUOuQfQMpTZG9aJC3rUcEPcWJcEPNsTq7lKh+Wz0SNFc0cBxB+ERXPCTP8L4
Nyj5lCsnQ7aFfIL/c0O1BAiMhtxyYapGhNb5XIn/JuhcywrTUySV4IfQUzyf8Yo2couLLwItUKMI
buSWPmt34hEQ/h3S3NDwGAvwS4vXfBiFQQ2oalgvN0CyxT7N4moEjB82u8SsNuiMOcmtet7u5ahd
Av5GalZu28gduOU1iJNDvwa/14SQHr2bZgNAE5h2j7wS6J7++9i+7wckuIp7OKWNUH6pcnRpQet5
WqiY6bC1SMpxZAqdhNuyrAdbWHQ4Dbh6ndatiz+KG1V5q5RxnHDd7pbJRHQmI3bcnY+1StXNjr6F
pw5RW6lz6ewN+TPumc+aqGWHvr9XuHUc3cYpooGhW2AcvB+XomSQIyXyocE5zCF8CIg/Au6G2vUj
aTEnPRL9/pYsfznTGjG3bF5ED1VNSDVWrdyt8CCECYtnPhlrIwxnlbo4H0qErwYiI6FCcBNsA3Be
Q/wmFcI/TTp41Et2GXaGZQAu7T/6x5ccWcw6gKUbT22kI4N5yH8JnXILKkJVhmNryz1c0yn5zGv4
qvFFNdNfkXc25SDBY8AY+sP6E+CB5lFw3OSZGPl7jPJiLtnn46bepRI7c5MNCdl25yk7oOa5B8GE
RASgjtwNm3iAIKf207bHlEUy5TlfhNg/VXEu8umyV/BPdpAlvQrJISg1FvNcNifxAG1YzcMZa9OK
SzF6aCgHqcv0nU+y8YTv//UCWlzW7qc3b+vDLOGko7i9tWkYXoAgL6CHNrzdIvNoT8wtdVslVCOT
8fH2w7jyLt/isU6UXOxAOxaHbfKmcrCs3Ru4NHAi7crair+OjTdp0EJgRdmtZE2f5j3po95kkbuh
mj8dqPaKC3k97DL9W3V2qr+moQH/F9Ka7UpvVNRl37YeMYUzTjtgZc87Z4K6B1CUba4t9nxqd/hP
UYOlEJBFJVvIFjlhZXWMZXijqpcddy0ZvD4JqYBPyot+QuizzRk+t9OKsIbpv0QrfBDzAccWt/2i
bMa9U1ZYcPxgjz1ZQSwt718W45WuqtfPtkC+n/QOK4kMwxWiGufV3zGBHR69pholkI2IoPESDfDE
1YGs9gvCIm/EpQ7UQbQRjJaDywn6y9jDqyez9KwWVKaYeD+LJ9HmAgBwx5b5eao80QleT0y52qL6
fTE80rd83YUpXI9QpJGYOQIAaMgpl4UorU09usDu4zUMe9PU5QLaHsWcuXM7bmxjYr5FNNZyYFC1
b/hDX8paJWk9BjMruWUY4944ecu4X/zdJOxwJTTB3f3XpT8GOIZ/ckuhNHpYfOy5MsrmoyAnccGS
m4pWop+Uvg7t7/AoRMJRr9AJRZ0npNoYpWzrwzriWPxeDcwIEbFmKzJezdgKquiDH4Jq4EevS9C/
5zbH+Gf3yPHPG7TvHJArWm4zB2lXGZq18oRH7gMwk4qgembOth4OI74KI2FGqBfgf5UB9HGJVHjg
jJUCXYWwOo50ThosKwTOIk5CSqj80R65WsRRthNlJ9NYmja3n5fWXVvcw7GnVfhv1kn9wvqyrZxV
HHjJfTFZEgZ2l7gsx4avuWTqT4awiVF1pTCtlDFir+t2k0YoL3GqkJDGnhWlGRLGHElsVRHr+uTG
KPyF2pcablROoY9NPpBEuyGa2FXmIihrHcIWncm3sx9dcK23Yel3JSC2XSEnbIs9h00UAF2iy1t+
3P71zSUP5qnJ84WkHVU6ZRQaIt1JJAf1nUnpdevzpzmYZcsnq/Y0y2J0t6KttgBX1q2ThfRtNMfR
VRW58GkDPcbiMztPfiy261RjyYklGwnvhO7I7vaUOWKeRaTf4XwP2nwx8f0D/PmNb9ZZA/LCBBVX
4bcYeFPUaozzZF9Vso9BkvAsFXs04iPVr695+v38Ak+tOf8lKT1tliIxR/D+xBiyzP8MlCCAFKk/
w8103xUfL5jilPRycovHaJpF1iZ4CmCaoSGWtg+/D9uCIyNz50PtVwKFWqKjndIl9Z8O7HXPI2rV
FTBp946Ub0F9iDfevHK6UxmM/mpc+pRo8NIvFrrAZWpLBMboRfqyBKIFHzMpC1Wnzh1pWasTEDJd
c5SKHUlMapvSzVLiA17d5jILNGo7w8n52qCXq+VCsDJGZbYJSfb6LIDN1T7QZN5v3s4Koh31ykrd
mMo7svObq/gZU3J6tpgKdjvQSYe7ZXk5NfL+UI4R80kf08A+ANMrYb5SZFD6C+74lUMg2DQnxW3q
sokrBCL7enTgh3qOYMfoL0gaLy0O2ph/6VTxaLo56JtJ+zbqi1E3rRQWFeaUl9j22tuBfJkMmXxj
HkSOE1zx1/XD4901y/IF3m30D1n61mvCNNHTYVWHM48beO4GZo4XtUtK3+mCpdHG6eDFPNDshrD7
St1bByEY0q/wPHPH/V3tAKcOBCtB6ZS2YW/pY62cpp9SYy7FueKMC+UrwrONbofjo0iyP4Dm/wf+
T0L/u5jRb0g36gm6l27eRgLMsj0bdNYeFZ8qE36QorijI9/5qkuwpddw9rdH7qSS+rGNxKtt2KBH
uNTUUZLYN9uMZ3x0YYbnMsW/13peTV+ota9XSBrZMEtwiFOgONaZZlTCG734ZbDJBSvan9x3HCmH
ipRvTJmgjSjAJm/VpaQrpQX3rWQ2XFjj1M7XHF+mLh4Jrq/Pa3dWdxDGdozM+o9J1W8uwfeNw64Y
SeQcj6mX98TZ5DRcRgsb4eexOZyIUG66gzfv3OCbKi/OBGfpY1yVQXs1ZvXbFcp26EaHo/LrXUgY
OkPWnYxlE5lLQEmdichxtP6BbHOfTxgcnoNZ9wj7JDyPEzsHFkCfuS7+kiD/TkgKGZMZ+tSXXr/A
M9liN3jQ5nsjao4UTumyuwTu4duIbmF/jBSNz34wQtlBiRydOEbUn6NvPszYVzO58P15eVwOIeF1
ijKhhkvVUdntdCOZDcNkDyFrq0r8g7Wi9DfgsIGm5fVTJVW2/gpFFvc2yR1MbTqIyo69jdXGYbhN
JL/qaECxVENSt15hzOx3PzVuo1vK8zEAqAi9bO9HIEOMUaXbn+gTaTc1MBiW//Ng6mB8GbumR+f9
L/QzvPJEtVDdnaahur9Hled6N1iEPQpQRHEb+uDh8TchYkerpKTWxD5X+hfsRTAAi/sd5eGwVPni
splCQbfttUJDEyWQdOWR5dFfC5MH6mtZUp8UOysdmyxZo6CEwmP0o2714rn9paiz9KVCRC9e0aM/
Owytg0gzVzKxcaLGbWG2IOx794a5yGQ1l6lTesVI5vQHVlbodu35RmfQjtywsEEbkfM+GHDoSASS
pIRv/jqPlQTJBFn7H2DIXDb4sX0L6EYqxuesccZG97H00X/Mz6Qub1TqjjaNYmGM4iKFt5SOL/Do
1w8VEgxgsvgeBaXajH/Jz6f7yVHpF2kM8mafEXMxqEhNcXdd0ugStfGnbNZSYzWmwl62BtPpwFRC
UYdjZgntHAmGJNaV/9f8f39zpYH0CfPskPa8Yb5iiEn//gU7bISlsPqzj6Qqe1Cdx9NHcgJQONh4
okwZLYFtuuESI89b4iy4rvStTAY4KI0dtG/yBU1sdocJ98OnuamjAH6ftinxIKH8ZW20IKneFiaO
Ci1lNGK1+G1HXaxGnpJwOr/0AMlpyuikXz21cYbHwCKMNnVgJ1RtgPogYd/ZPQmg33s6Aio5zkPy
3trWlaAMlHRabPqnz7nZH3vWtj2wSoR7BxT3xNcUqIjb/vf/J9+JXc/tFm8bivTaQm+OH/248DYU
xgbJNJNiGDHrdCqH0yT/sTsqSquEAFsfqNuGJIobxiEiRp3Ej8WamktbQKbwwicg+M8BVNs6VJcg
mF91+6CCPZHZXQz/p7pnCKdvGS2xW0PfzR4IX/iNy1RtkXaM4xP7ciJSrCB0KtBd9YN5sGxeIa4l
IWHsDLAAzrlpvsE4dFSaoabM5tQKpOMORKaauRWpFVeIX4LkN+ZT4JJHOoKFu3pNJeHQjp04Vw6p
q+i9ZbcCR+xq6wFOKZYpigjZDk7JOhfAw9+v1Tab+v44RveLJh/ihcZS50abxBk8EMy/8hwrbijH
W8ckledKlRXxvWkRjq/oWfKmA7X0PiDQzGL/YCWyjFtkTlpjcCKpxP9aeg3/HsBTzR4F2N8QpUvz
7TLzpnJ0nZmsLv9ZbzgACu7LhW7+TMc+CkZ4Ezhg4IIuxTDi5cGLO4W6Gd/7E6514voi5RjRuYEf
bo6rQxXs8YUAaOxaIDtZ+slbhICtfMUZAHL2jxc4eUGBxuQwER8hxOHUFYGmlzVHZW45+PCJo5M7
gqxJg7KAscZsVky8lewScqaDiWFVK2/Le0R+j0n46uMs2cFVtsIwJGykkE+5OSzviuZKmb4KHzdj
+cFsGiprpYyhT44ze38bBicvraURVuAj28Ksbja5pGRpnq26dm26Atwlb8kFYUVPimpEHgqZtwpu
ZQd9viGxmOlcfSBjgx1YA0QmGp1pohacGnmU9qYSnrdxLkLIN3ZzCDPvY6A9khzBKiCVoPQogvV6
EZ4v21GoDlqzqONk6PRDf4eJVHLkZfHlDhxRntosUuOLLFbpcZiEel8+7/Vb8inqXnR8o8FviYPo
28ZxfGNENnbcBLy+A4fAP0EQ0FfbBBGGOSw6UXwDbAlEge6omR0r/1TsSoZoEoAvJhdDt3HHnu6q
/FXgmFMLDGnRq9wIoVslMBC445COvPc17hoFM4dwTvabyCTfGSQ7jt0FCrBAzrtQGMyKPg7AmfI1
N0vswS6pC6r2oLN4pQm8sFRG7SU/6aqF5b3JokPZepbCBQNzs4D0qYaaMheK/g0Ho598UjP45BYx
1Zip+gJ5S2ELE6UO2OY03c2pTUJy65npfRNyHupL5bSRL3LdTYvD3S0HAbhPMMAYBSSk9mZmvk+C
DNrMGJjAMMb46yAWusOpJZsg4XgYCyED/y+w/48CH+r7c7xNYm3765u6QtpDd3D4XerfwPSA+ST7
XwwOY5rhYsM0csooAdsd9aJ2El5TTSGPju4yj4g1fa4gXcYv4bruzMcQ3KjkSU5e24ofkk08fSqU
iLkSXeEeC5GXw+2S6ovcFhdbs9VaDWUV967dKqqLRBHxrLEHCKanSWYX+Z7hJlFkfNHSTj2m1Aib
mxwkNsk+hQ0rvYG7kuJvOUDQynv9+O04CgKgfRdcyK+GZEfv60M1xC63HrJx7BGO4B+oGUU+0d/f
yR5O51bIioBCMbHIqB5M4n83vws9gp1FAojfKIuwZMtLYx3IAPo8Mt/xbWGbU+OhJtAn3BZPQrZ6
RdgZ+5amgwtlTQVr0n190J2/zpDRpujZqs5dIv832UAIn2V3x0XDt3oHnmLOoF2z1VzwcU+sFogW
OuyH0ToCNWKD3WJSDBKuhuGaNJho/FU+DQN55irQlaSOn+oVP3qYulUOHG2bUOkfCLHnyI23VUmm
TyQM/tpIG+qtG11um/0UCa/L/zlVM61gPVIYOijGsBZeBy2chapBfA84fcg8rjxc1U/t13GoCTFw
BL21jumNx7GcNfpuduj5rIgR4qMZCvPe7N1+mAEqPIdVJtT/WLKmhPFQGqHEVe7KlxeR8r6molpr
RHkTASfxadJoxJNw7M7YfWg1XP1JxtibIE2yaTMjs10ZJkMKrZQUWgAtrzWs6/5z+NJhQGyFq30W
/ceTllHxBXJiPtKULhdFCpQHHGS8lwXTlf7Y2UAxkXWRQyf1zEuPuOtogunoUUDx5Bx0druwoMFW
ukGRCluW9u5rpJ7hdCMnEk2x1cB99x4byBM3iBlroJYUJcb58/8PPgm5O3m4snbL+38ijy5OyN8Q
zkJEoqY3P32nGI3AheysvptMczp2Hp6WoDKBxdjX5UVI3W8k6XYIRfw2Ne6qxi5jUHH4WfovD20A
D92+6QoQW53Ftqt2l+seKXK/+mi7wsQWEgG2S4symFKUIsiIDkAdSr4OTxuqQKFnw6yZvGi8cByy
5xk9+FMk9JJCbxF2PooIgV4VNea56sGKLWyd4LlTrjDl6Nz5rQfFoZiknwJBa0lJVGWnZ4bEpheM
/Bfot+wdhmZOnqS+DvK0nfv3ZcH5ROXqZtXPrmPQVgJayGs4g/L13YQyXlByaqHAWGkg+VJbOG1i
PH/q/vbfPEca5xKioWrdtqkUa1z23qsTVd+iW6bXaM9GcPV2pxEhtSOI23lUZ2tjxsTzAm5UbtoA
+pUqYDydu2Zbj6WR8qci8Rt7wOoe/VUL4kmQraoY0ztad3tzhp+1z4EdGcg0HguTWhETIXPV2RFv
wwLO9Oc9uXhPd+QUJWpceBcGrVyHByEsR25vHnjIA0cEdRYbAANMtaSKp4paZo4LJ2pc7ycegKYT
XNfDbI2pS2IBkdosTk65HPVkdf7NCBtKfdMMIZxfxvQXCwmx1LYWhu3+2COzt1ori2EJ++i9uN1N
YXTclObB3yUDiqNH/g9H+HKQ/mSA5b4QGJGdZWgUQMh7wK6R5jAUBLw0KTXZPIkdTwr26VV7HDfr
rpM33uoEkPMTIbKJAtFyFTsaHRrgtAEJIrx7BEJOQ2vm826bHvenPCj6hOZBJTNlfL9O4cGsiCuT
xt8xTeY+3J9Dea8idfDLEpSQlj+WsR9GR+8fw75y6uxuLrbcAgixsfTnFJVAb+klQQN/e5iERbn4
PRu6iSlsVLy3XW9n8RLysFpAcJL5GV7JNo6iWReOO/uHAdcky4ZVtAsEZLp9FvkHjDcGcC7DI1sL
f99IrG1Mwiyc7g6IgfJwz5i+4Apq0EU8+x7JEgqMQjPX0Id6gC3j3hY823ZvAQMz+AgIYDSqeaOu
0xWSJpt3Q1E46J5bWxoS7/YGNkaAMvjDna5iXLJsl3hEVi2EqUnLbgbxFbnEQfum8G6KLU3igrhA
jd8vQlpbeWnBK33tLiAzHReFwbs24u4HIJAuEaT+/wrQAXuTpft92kouwe79y4z3bwJPa9b7W1FV
1RxpKbWexSKkCj0NWvaJVAMF428DqOdoNxNz76wz7eZZREpsiMHX+2Dc8V82xw/tTPpWTCqBwVbL
IyEx6AELDp1Bho6zYsu2Ba5snc2nQnCKx8M7mBKAztQX7ELg9kebCbgI5J08+mv/AF3HAcgfwn10
1jsbdFkwD87RXBTfCTI25vPYuCEVmwE/JU7CvlWXD2lOd/udB4Q+c0pbXGGbmA5KXEeG1ZCccN/y
iGzZUiX3CxvVdhtUi37Ler9P8cAgPSa3rIpvd73iz8+25mBfT1CDnUm9bR+w+T7LbPL8EgLVhVIR
iZuXULYkw2y7txq1Y8jqpdwWvTCPmIIvvCT3k962fRlW5JQVWV62fr2KJWxK/fSfhXA6yXp8pFf2
B763hO1QJNBpojVeTgDhEFaObwx9q2pIpXmKQTpBpkjqS675i/XtOtLMveFnp7X3LXPSxesfTCzS
Fxolm7QczjeT2Y+qDBSWb0W28BlPYTVtzH/bPOWqzi9Gs2T2TLx8+XRySBFN6CPEI9KTOM7wGBVH
ZLgw9bNI2MTZkfyTn5g+ls1yrQ+OclS4jgpfVvyUevIUCUOLGZpYRr+2PrtmKzdoX0vT+upgIK1z
PTlpYjVYBkOnMW+Hjbej7uu3C+CflPYqoGpXjpAu3gnZiinfDaCca7ifdoth4pG/VbkWzad63YhV
rrLOcUt/HELaFf1dErfsyVO4thK+azhbfwQauwE2cdPjafUTkUlYoQhRcIrYWOvWVDUaN7TZFFYi
G6Y4M3xdKvDSQ7QEILIm6TzluaYdBnGxmvsAhPyjmPn906CAC3NkQEtmDw6fdciPNlTPFM4QVwYa
DH4XF0IsNll43xWUsla6IMgng4rLcpxeYVUWr7x4KlvyWte7JloHWp6HK26M/pz5BR0lv/fASwLp
kN6339huKZutxiHWXvx+g0ZoVvnpOLG6AuBKd1CMtRDA0CWe7x3ghmqg48Dg7w5jCBv+GBTp8wRN
6XTUS5YuguH+h0Mu7NlS6yq4lEEIfCBE1ao41biqPdW8h3eD9KXOfW+JSZLezIenX2+B4vUtl9ob
xKJXmUXXaM7ZztRKi1nHPOE0EzRRk46b5L8MI/Wflv3X4lt8E42xuaEy8YEz1rdV1UT9szzEaMhG
lDiPH6nLlO7/jDYE9blPcz3zrY7PwxwApDwoSR7T+VHf3+e9cB9WArRrlsY/8+rSM6LM+NkEVTm3
oYoviqmhlff3r5qsuHYLjEqUHeXfvjciAONe+QP7jw4EYPHT4B4R55KgmQ5PdF1NFA9/4vZ0jIYa
nWWyVpNTwtLRq69ammhfDfvmeTdBMkOkANY7ULHB5SdaXrukCd1ko0uebsx12q1Ao+9jkLpfJVdG
gdDGlxhcwOGJGa2gcbB4SjPT3QZxcmSru/g/mVPnLjJ7+8ed6n2/Wvsaql8GNcPeuGNTSU9kIaFL
rq7TnjNGaF7QK7gOa+774Qa5MUnlFXaKY5fEoOJrfor59HOJyK5eS5m5FHwVa8mOhMFfRi9sHTjk
XV46dzhglaQjcjWx9EqQ6huqm4LyTFQp1Sxua21LeXJnwfrGtkZwU/0eNO0zsD+wNvFCQEhBFGLr
45H/RTsg4lUCKkwnQai9CJKRhCpVMC2Z6pPRawnjLDULyt8ectrJc+TNEoh5OVHka+0Pt2mrEiBD
vVuspIqloRB6JuCzL2Gm1te5meIQZtLyUEK5UJ5q62sn9j2DWTF+PU65W3enUh/jcL4lfp9rZ/Cc
f/BA9/puW7a2AwinhywXIAKoqnT5pJN+3zkGKjRDD+e0bnrwyggXWoeclDn5GdTG44hYPr+bzNHQ
xQsSr39MUJtD+WeXXGYRpHWWoWHW4t0PtZOIW1nrJ6oH9siaAVibO1MD2wiATvFgeYaJE1lg3KKi
21eTbR/c/yyuGVpRe1F/htt2ya4dHIYuvk0Fk4dSEPCK97MbczKv4d9muuyRpPRAvjQD4s5NpJ9D
bS0iyz7WZLPAAv1CDCZfRWXaUDfH7ksV1Ex/K6roalE36000eAmXVjj+1GFlYMVe3DpLviucix3z
h2GFRJkX9ldqHuJWGfdcRUiVeNxXpkxhgWVaiqDKfWhDOL7KAs/p/YX8yXVE3WUnQozsEaYnrSdV
msEpJVjujL1GHA/99A2Z//kwtswEpSdGrsM7GbBdWiZrKIAcYfdPJY8MFcsnUfswAJMVDZ66zQ3Z
Fr6J0uPqT+rMukR+8f8V8pjdpt7yNS7plSar5eEiLVL3wjicR3JW4AaqXNcHr4PRGamK+VosJyti
6hP/H/1fndkhylT5rbcJqupnKv5CKYI95CMw99GncRmsI2HOfSurnlvQXbtwfvnXmSRNFLQ3KtBA
HErg6gPbGp/CaWNxXmdudHp41WQWKV+XWpB8uOMmSToj7XL/Cj7MKYv2QUXKKzSr7ohYDc1EJQU/
Fb+ZHVi4cjgId9wvIH1HIQLYw8tKm1SHpySJd4E/6uP8B6POHTInv+3dEy+wSONv6/xtCgJMqIDK
7awm1NZ0S3W5BFjPSfwKeqCpevlZW3RHhbMjpMBPFHMspjjox8mS+fsrMgW6ujXoQgK8EFMaoHjn
mEH0IDQSFfF3knrAzhMXf7PyaRdhmMi+TpWcapcnztBqFyIi9NSHkPwVD5yWyGhN4XRk+ZspCCxm
CpubYTu4eAHmBjBGGzDT+U1oz/b7lKCE9/1fQxPRjVaXrsEJR58RoQj3yReHBj77huEhlyQjpo+G
ug0b9CsLbn7c78sWlLvQYlMdRR2kapRO/JfxxaIqitVB/TGy5d81FxQIDcND0V3ooGFRi+A3TaOu
zYYsm1t6pgnuF/k3hvcLvpYYJb7K+74q4MDlh7yrRM9Cb9UjBU+DkWG1DL6zZvuauuGMNfpBdE9h
weg/VtehivzxW/s6STQ01NMSTOQMYE/RnMz1u1qk5YaUnuwuwvgco7DCcwcOZWWOeVYOOLcOIfU6
WYrG8rhlkzSwOp1DOm6mm8+wvvTHvH9Ci5XpZXJiOMBlByr20/UfRIscTBIlxgPd8khPyKaXmUdc
GgPUsVCqvvXvElpAnz/YKDTM4jWDjDN7Wsqx6cO/N4PoBNQnfTHax9gStp4iBqiNRwM7MyPmAsRh
nNsLNV1hX0DsrNo0bb72UQ+i/RnypnKNIhAgppuh2FeCDfds94tuLj9tX8aA+PvX+GsTnTIEaoPG
dwjLYnuJ8pAdVpF2q6R2fLDaV+tP+sa6r3TxfiqFZmDyWad+MU+f09aXWbbUBnVk4VUyTLnnZjFF
emCUh48NtiXun2BHJXvLxnfvMIf6C/LN9VhytHWX3U2n/VuXU8nylNKZf3/rSGpoJMsox20SOcjU
fPQbPntcI2kCWn7M3kGSdYCFOOi1Sr5VpNEdqGhNwBAKJQMNucbDpvG1LOIpoAWb8XcQ5VqDjoO4
gQBNLMZutinLl9JQFRe1k/x0PQNvrVVw9iGhgZfW10QBoxaDuvCJlyFyIYC5n1M6Ql12BMIvVRnP
Uq7onJSaEJWbVFP1E8TADZ4q7t8eplhbA1HL6vEaaL7tExOJ8oBtWYMBx8H4g+cNke2XRQb9QOhc
4H8UsFlKaC9jdjhFlFXsRIwEFx2KfqXsGYceI3OCtNQpqWugI91wxBMP8+3MnD4D1CM231pQ7zll
E22iMTYb6zu4fT1n9gfj89gkT8Iw38CCPThH2Z3s+VQYHhi3YCZP6+OOqxnNeCvuM5l/tDTBUd04
g0ZQf88yFUAXJ+77ZFV70xikLtMQs3MKzd9ur7z46uEF9hMwSwFe4IWCBBzRlXrtfNSOsNu2PKlQ
81R6tpMq17wu7jat4fPWA6qttepxpP1oWmUSQXBPa594MMI/CPNiUeaQ6QQbUiRwHAQczSK2Gd5E
AwVXTKjNAfTfnIWhoY4aDkDH5gfPp8yCWCSqSQXZfCt8Xiz05mpovPhY1GRv6f76ttByeLPcqzyU
eCaq6vrCz7WTNxsF5f2zxqQC4yz9R5tMLVKyTMmf3VM+WL7lgr9KZDA1hiMzQ2GqGFLL6u5Q+oRc
XOWtPX8ocxgk5VeKPvJj9M6s0Z9oIEXi/p9aHJ4YbVp8WLekcbTWMLhmaoR2Rtk1jNHnMvNltVWO
fMu9knA6VvZvW1xYqN4JXmISLB1plw3e9oaeSQiNZK48RPX70l7CQfpfx9ujnnEkSHRPtplhQ/kP
C7lpGCXm5fYeetDB3gj3UKgTtuK0qGNTcrDlDqwRGy54Q4Y3RZqU+gzg3zP93phAHGqWnnYF29p2
5klygC2moThRTJpS1zVw2qe1XY7r5lMMq3mghkxA53WpYOSsCYUUZV2EP5yhA7somz/xYv4vs2cL
CphJlCrJb/q/zsRz5TBAtF4/5IqeNgMuHJMmDQ/KX/iv1cBDq8bQLtATneqxYErgtk1gokj/C4EU
vGkk+W4MrL3vZlA698jOb98JF7KqH7qY1rt7QRzet4ctLrsRmLOYm4TDMYXjJzz4M8ZO30yGN1Hl
RAn72+czJBj93XXaj9ZQFYGaLDkZ9FpJ0jdYylAITLUo4exl7v9CapcFqlo2Zg6mc//7lWbRtvFj
9LROMM/ln68GGfJzFD+B6i4oc2yESPlafRv506/RdViHUTkaRiWSe6mHHh/MdtGBl686yvFPf2L/
/bF10IFXlTfUWFbRp5FFCrJAsWYs+NddszxvEvLuaSkoHacQWjBP4vUsu1gIKE8viXUH6McQ3/4T
zR1NHWN1lOpGUrPCacXY8mAWGhsl8bBS6D70lLQYfiDbqgV+/WZYbnEo6CKUhj1vcJMa9jG/vkDy
G6RrWfSTTo8SPsWOlR3vU71T37bwUt7inP4A04cmATF/6adyuLnaTD7LDg1w7tdXPKYz6sjIFeCk
cOh0K+vimU9IWUTxLgx0OdOv2GvJwo0F6CEvwsHWQkwW0Ntszmg3R9SovpytzUjnJbrw9OrUlPbn
JLVSi8uUeL3HRMPKuNEJA0jqzIXk+NlPO+6Av5Ot+EeqqUfmZsob6gW2BtmR2bXEawQyQTb/QVTb
3ZIU6YqrUuLnILDORb13aVVd/LyyYXbM7Vm0tHOoxyt/uayCu2Ljbhrt6eiMI0xjbZBkgz4FMkM6
/gN8O8UUnrnBBnenBNN4zQHQfa+IyO/S0oLrjjRoEBSAIS6nOad8ts0sOzQo7bhRicCzY5U3gqc3
fw5rFZQaDLunWWz+BC7RiQfWpMQNiwEobk/Ok/NWYVUa1CumQAll1HRjaWF9IgjpE1b6X9aQBLl6
Uoq20riIoZf7DfN+338f2z/pZaHtvDVTDFUJWZaUHa088BJQK3G5a0EsJjhCq4NTDKzG1D2t0qmJ
EiKlb66zMq6lwTOVEximDrBlveL0R3F7/57WpR3kCxsfLoRQAod5UTpBFH+CGz1pahAKMcypyxc6
zKhkvMEokfy6Yt2S1CfwsQNq5Bb8tyPy3+nOJbDmxfzcCY/45b1lLBXflSgUtCifIOZKBbW2Pxes
5vKd7Xm5Fk3KaQvWZEJnd6KWeZDTTWYFjxOiwhWYOMHknSsHVs0rkcbq21HiXncnc0gNHoujwQC5
7MedwhdnumEwv5RtYFPP8HkQz/iT+e7ITkC0o0LjxIl6zMdVgPEUTeH4CXxiouOe8c+xVimsPZ72
GklgC5fdS3M4m1NJ/9iAIZDrUjYjHxw7sZT+e10eLlMHK4ADi6DgrU7CkU7rnrzJimiPV7IhUxxo
b9yEO40QJRmRIZl/UIQEmIClapz26fYNfSs1A7rVdUkUQFy7rc+h6H+1pfNmT5tzHpOtL+oGko6/
jHuA1KNxJSggDjg/laD/brGCxoVdhNzD3fNvEdzbEzHE0yDnrla0AYoBWiZnLPTghSNK1XfgjZCP
85nvLcNcYjdMGtOf1urQCeV+funuKzlI/hpTLhFhHR+VW3b1Bd6drPHK3eDPPitFbotDFd6120ZV
eN1yfg0NySWGRn/qR0Kdp9EJ5oDj2sBPzgziJm/A8l5W1/ONwIEiwxkHoAlb1C69cDGAAQQI/JUL
6179pa1DXuwdoORUnqWuCXO6Z5F2vo0v//cqoSrE942dLcQ9dqd/CKWeSjUvWUY7D1Poy3ffia/w
wU8d3kf84b3oKFtFEQR5+5XwSz07cb+O8ANql2F+ynJBBUNBGSaoO/N5RoXcpMINUVWMWNz/U2Ns
31tCssOAAqZStfmWMUpjF4gf/vtUDYZv1ZAlPVuZcZ4WUE0CDMIVibgnSII8X4o22MTLeQm57DX3
mtGK6N3QVlRwDhcdaRwz2lEfY7dTM3Sdm00yvsQaE1EKlcNiRuYUuPuYI0zZKvmvf7Xo9BXf+fyw
6hOGBPEFOHg7O9oIgiSM7QIqKcvzazciXVFcLNgqpqrGUL3UOdLu5ilwaC3DrjXcMBaFBeJtWhhI
wXxbiybAuHv/Ci3DsN8OWTZ2ehD3h4bKn6Uxaz8FjuaQZiO4+U7LWc0AmMkeQ6Kf4CT5dtMekrzX
jUDGcutfp6Ftr9JWU3E0HAoIb7uA69qCNAuqQ+QAko+3YWp6ng4DmKusc2dAjjeg8+Qr/Yp11a1n
/fig5CgwptxxvDdkEBTzno0rKLE2S1RiRbO21GgmHMrALuuSRJ/BfSUNMNcFPHnQ2sVTMnZ5CLvZ
hjm0B2pPhhu17+Nnl0nWk0YUD7ALEyP35ZeMIwFEtcU/xSgG9amVEaTj08A6GeSDpi8h9BJDIrWA
XVTF2YJEH/BusRjLsRSqZmma0aompqXAPfMcyGWP36EKbOAZZjL0FoinY20rLWvN8l0R1T8sDBhe
KICylx21o25FLByHemtPBm478wxlQZmajW8xP1vMZjia/QnUuPcy5ZcWAT7UPZQKi9halwZt6Da7
f0iejWRrS8UCFOYFLwimHE+EjVPTXiTQbWAyDPOOMqRRkLZjqNQA1TXJ1XE4H1Jx/1OBFebTN2zL
NrkdAMy+f0zZhmlNkEOOadBfMKo7uBpxI1yUhth14yZ1mnVoMZG7DgxPJ4GgUPoj3cal17jVyyzi
TKKPD9vRkM9eJQ7PRHreESJurircitgQDWYvjpAVSQZMPkMMXPH2CrdBRXKJPvChcfQ4TdKzJ/vQ
NXA8sbQwriEyKLOzK7QZ+PESVQwVOS5Iz7PAc4ZcoCpYDjSRmWL5U+8cJa7dXg/Omu7O1EzHmwyz
dZ1XXv8Z76ZQ9OturlF02HvXi8mODBlZqu5LmcbX1gw3//523mVKJUPf7+Je5IsZxdfdJPNPYTxS
tzfZ96fBYp0K0qvsX/EuycTEqWRGX5DtuJex7xGV0JaMcUFFrjlaDvu3OCBTGpmQNRoVQqrt0yxz
AsFQ9ZnZ3EuGQwQV25HqyqAcSUboBoIg2q3w56SYztfXa7Auf8mHmyl+tX9A29inAB2OoiMOi9MW
iXU2PT4qqEOu0kGfKurzM1wCoaT4M0+S8IwLPKG3JCbSOKB6Va2silKlJY0rqfd2FQq/nUN4ZbUa
Gy5gL1PWFXg0HWfPbNNln99niS64XSqZGMEwxzU2AO4iCrFZ4yg1XADif2XpXp/OplBJ5HIJh4TR
4GCnrSNWjk3+qPgut1QQYhi4lTHdKv4kiJkmoOWjwbTLeI84dEuixCBZtoVUFJEqCa6+H9bkFGAh
fVuh7aedM5gssqWOM017hxBwNsRQI0/i9aF7/WwWE/mH2wuJ1b+0stXA9a1AFQ26yz2HxnuaFKin
v4Jcpa/hW/MGp1iF8GE0qBzXjyBpjksda8DrZhZXWBAjBkVsPPNtPrnG022o3C/P5dD3lONo/XQv
UfTySjx1xO9LrIFMFjtF2dHyTatf/W8ww2wxesgj14y7ooDyHi6b7fKco5cG1/Ow75m1Q3pklViJ
dsYM4jYSpGPtROsIonHYY0Au5gCoTSAXT3OmpCzJSHHrZPbWGwWDSwXTaonzBbdAmgUeC/OhEA1t
nAzkRs2uAw9p/m8SUL3mfKFHMILseI2LGUwsJa9qDtKcc70v3XUAqIFEinf5mwnargDfhli2Ugzx
RnZ4/ONNy8EHz9CMGTlNkC6B4QWSDgE6Qej+dn82UTbuFz9ABqPPATUgLW2JdaJyovi0S2EFtVaj
JBO1qFnz9z8rs9PjJyRggWG+zChZan308e3zc+i468FNXpuT2KXVqigBYEYqH2+TQad4QPdGsung
ZZfMjDbEKZ6IR9LXxn3GWPwE6B+4VziTtvM5pP31xWTU8dptVEK9GzuYq8mBvt8T92WVGcFKPUKs
6Wo1YkCD01b7vJK9fhIGIWHtqJNRw8bcLZduKOScKykMbV/2RcpbQlLPvSUlrBuAPFsp1xLo88RA
dcr/43wrHHumlwwZ/rQkES+2EKwLMvZ1JdWIFnQ4KVTHDSUNkw3m/uq4li6XHvQzUd6jgCDC7Xvy
bIBeaKXIrafABZIDN3mx9n5+5mwutv7qxakDpQKrYRt21bNjOinOHD45ioKgII7CZoDhae9UlkJL
eIdx5a9d54sjf9b/5rs6dBChbZjmUIw9G4qIXTePTYjVQFjnF1mtmAbGgHJ0T4CT6x9f2giKhx56
9XwRch+arb5YHR8anoHqB8/Fxlr/b4+jaHDivqVTekmFp6pCi3QIn5ak3MEaDEQELKHki0+gfVqa
/Un7tQOMZv/iMFklMldevx2uwonHdSMAIw95CKEZyIAE2LBQlfn1rNCS8Q691PuaENyOlkT5RiOE
UHQwiRkKASJo+UKR29oQ1K4qMBiEgs/1Rcj4j1QP2Dke1J51bFHAWkEuiDIjpDxGKYuW69kYioGl
yBHCMm5VanRurJrX1Iuq+mH3DpLp0M8gvKl1NMnygdMObOffeiBeRq8PqiwCOWBo9+oHBKUIfsGC
2lr0z/Re6xGGSPHV93ugdA3P0a4qQB4GdlDV0m2B9O/J89NfsJYs0JMm0K7AxD+7+fvwTBocrXly
neVHeCRkpOcQ2uBomr1QJNgZLlfwv+2tFkxwlifzz75UUC2YTW9Rh1kdCGf9M4QImG4jJMnOB9S8
uvJJ/zZgOInU8Cw0ESbkJ5pJI2GubQi3BJfBFjRex5eUFw40Pj8YIqoXa03IV4ap9i+OPYMvjwxJ
01oqV1Tse9OMBf+SsCBfBC/ElKu8iKVcpmb5V7h7mM4OTIa0AwrSWwJge/uqn9quYdGYvJHQUEw/
bQ/yHl9Zx5ECQlMud00FyDcRHBTHHvTE1S7lnSFdcKSN+aOY/rXufEBTv/Z+3DsCa1gFjsg8r7zj
sjxGLRioXsmAb+b2cr46VKsZ0b6i24X33Peqv1EmwVoLg08v6mBXp4/u/1oQ2BQ62Y9DNyB/LZMu
53p6Fyp5CAnGrilgHIhSr/Jxfmqyoss9QAw1ox5ZWCbv+UXjvl2QLyiCnM97aV9oLduWeLsKK5FL
R1wJJCdkpYAoPLds7wNDj7fpTZMkh1I2GT+Lc5PgsMTsPXDuH8ZHp/g3fy2s0vdRjtdww38Vd9vj
TeRhW2lXr4SrcRdSKVXPDE9dAeEYnG2QFXi7wjQqQSga6V1KsIpYBjrQf1KGUl7i9aRCKNSjYbmm
B9schFtO2PEAfowr6K04Aey9+BkI2qHVHS9Z8NQKxqyrDHosFCeuJuSujFQSnd7tbi1297AMSUFw
rWyiyYilzGu6E/29t6tAWvkmMc2BbAuZgqXyWaHe/MxnBwX+JOgbKU66CqxQjy2poDfuDrwNeyx3
oHrw0+PdlbCl/Hux0jUvX2jfBpkYSX2lZKMQEqs4WaSOtDHwQcKJcQllGK4TGeRCH0thWTLImMCS
dJ7WPVNZokuyfZ4FlUA0KsuyxL+625jeZEka56gs+rE4kfU59ZOgweVQlGuiS/Ig9fKPHxZYaVoz
Yjoh/aatiiarqlm3oBSDsYeiUEc/vJA5LPsiqnVw5alUCiKFuPqzGZw/FqgzMpOIjo5bZNPLD4bY
ar+Cyovbpjyh/Zsz90VhIrV/81EZaevnC7lOfHp56Rq6Py15hMUqBtIeCohqj0KEtIKqYnfslPih
AQ9hqF+FLdeVxUUSxIpLNsL8WiEQKkzh+TTGQ+ut/05STRlCLJRPdrzLy3Ot7iybtbmqLnkZBUYv
2JOLq50ade7T3OhBVEtjLvZgnITYHnUatcPS2ZKPP3SYz0A8PGKx9vd6+jF8nlTIf8oynpPlyaHe
KSr7ptJ/A4g34XmXLAWkOQ4lucMebOs8E33T3SIvz2FIt3rfJCITHijfCT4j3SihYT2oeRuhVYbw
7hugf5tIPHDz0m4yeir/Ul22GbtYyfirSLsb/SgAdCfczYCgUyEVacuI467st7+70hHCAOyUmseI
uhQJebPg5yy3cnu6LAcQyrf/94efMfHfLaXPIaUd4feJTrnIhfaspLEvt4IN8Yh53n0QZm2YJldS
mU/hgJOC/ue0G14mHW+3/R9FbQdNNXKPH7UM16DpzRh6ohu99ls/pNacnX+XPfO3vYxsIC5GwD9w
LuJ8KPaIJcQPv6fpPBA7L+eToTl3b0ugRczVrPpBPi4qSGfyc/ZvY6D8tS5DzLhWkQLpH3dYiKcr
AgsnvCt46fWAH1uJxDoCmvaWrGF3JPewA2BbsLXY+rEMwR9VBM6SmuEpKuDpXS4Ka+2wyAhQthEQ
10qHeLDOeJvc1InBTnoNm+rD5sRe7uujp0wzymnvXg97KMkehAhvYFOqhAMavvlwyAEAxWOJWyGV
yT6TyBAW8nUj+UiuWWjGHPWemAySFIwZbnasfNFw+muwfHggt4ljzzQljrro2Ql0TJ00WW8HKphi
gYo/JPqAH6rkFg3oUDYufUI174M//Piv4fJlyA5VGY+Y6ql3aG9pI9Cs+MYuWcX92OmxhrMGpgGY
GCqreaDtJpyLoGmyPp3kSTJe2mRlsmcK6o/D7+W9cO0d8VpU+F45mRJkGw3f1cnhqGCsSNPpaSGt
itz+UMV/YChCPYrClDkuhgWZKT+vgzsCXmXUBVPgbMuqQEkXcut+WDyZKQQWnaVX48I/0qArsE52
nY/DM47IWxqh7sgo3/q73X2QKhaHbLu7aJwSq0eFKirjrGRXPKjDPrQ56JVsKqYn9XW9m3wCLMpw
6XD1XI0icu5gLeV0YmjDSf4Z+GqQSIhNeS4enmYrNwIpcFyJUOrtRxcGbNyyf4zPtwsl/1cnbBg2
bv1vL8ZyKt0Whx7yliOXAjaFe5JABEEHiwop9i4vGrzjrCQ1uKqXDmPSF2e8cF7FJ/ebGjERKAfE
7clwRFq2MzjWlIewFmyZ861/cZm6rRi2RmBO49B11ab84mA5QQ9S35usFHi/Qy2UVu/74OZio0mB
8zjx83oDok+gl3D+LMMqzy4R/QvfRdCKTz8JjESZVC9/SPvvzl4jLyy984QWylVz0fJOcafrwbD9
rX8IE7AL91uRxDIfsgK96ZthLOYqATxvKVta1jZs0/39lpuLqemwBsm0Kzj8W1qznVUtIX9WQJJw
kqnSlcah76OZnbbIBUGmPh6RTqYr+hDywrxXm+HP0MEaH+3y/3ZjuijIKewLSb1eycP5sfwKJa3r
boGcL2UUKQnkkiU8yfiwzU7wc5ny6MNWx6yij4sx1BLXI7vrZgm/XTf15WvDLQM0kQy9W/oyzHpT
t2C3/ytoMoIZxhvI6JGi4qtTCdyYEMIpwqCakAO0Lp8my6T+urKEgNFPQ8lxCetpjUwdmCyuuAVt
OJbqfLrRD3S9OV/x3eAqNlbUix7y1Joec2ddCKKjq5eCypcILZOCOZdLUX2PzEUBNEvp+bUJk3bk
v9IiXrLrEIIwsZ7E4Rssf2HafFrwKpYbQ7jdThHeLFlNMasB0+cGVFofw2hb6oSvGGyT0iK4Fcvj
KP30RMDQueBW4tSSRLLjlhWcnMcvXQ8GKRMTL2XH/uGq2vGyrfkwlcTmjAWliEznYj8iK4zflkdy
bcx889JkZozeTAe9Xw/Wxpj8TwThaNePQRqTPGU2PGqFFnGbTdkXJwotEwFGdzUtIrqvtr+z7Vlb
8Yv4kggbfzIyFKw+AdRD+QjzTNB4USMHgMrRfOfVhGABo7gTOK23t2xIIkd5efHK7EeXjNCThFj8
gs2nyYFoZ1y+zqhXpWZVe+YakcYzN2YneWUDzTWtOCPsLYlZQEYw+Mf6aVGA8aRChoSLdQQi+FDM
gGbtSHlq4y8IeaLrjnW/7TqUiaUwTZBnEJpwBkzN5wROltdfeRBPlH4myGinM95WFc47y8jAjWn5
3JIzo7i7HT/RNS2vvBFfT9i8z5q7X2ItaabQjbYMHu0zVKZdZ6Rf36PsV3b1GLo9yl1V1mjg3OPV
MqTDSwbpC+QUVXl6vNCpCPCmOgOK/W4TGlc/T8WtY24EObrjIjFTH8/P7P6k1j+jQ4lZr8OPGp4w
wucr0KacOmz2skN0VXbEt5P/oO3ht6B3UCmdpNEJiDaht4o6ra5274f0awWwnK8yVGtRyhrB9SlL
2VPMTgfzGmF0BrslZntwKVi18r17xOLAiLox1/Z7f1+npZRMeEEYK5jVtRTmR7HzM+PQdXwd+Hq+
XOpPEnS+bNXuP7cck9MnKaVmf1TWuEfnW117a4J8TtUkzjqXvy5eRS5wjHhuhoG2CtYdNj5xDIjt
GaPjfVQwI7K3OG01f1A4C0Xe3K/rOtXGgSSnF+SkWZNHu+q+TDvajgqoza/vcpahN81l6ypx82iB
6J4aUqbckm8K4AwfQV8qN1cS+StiLRgnn4nlWqz2YveLX9afe4e2TeOV/kBRpW+plo9XosNX0Bd6
kREfsz/gLHExckEx2rN+6FAbo//9xiEROtHmMgnREDS0T6NAqOzQCr3eYxo+v7NWjKdD9BVx1rFQ
kM35xPkhtzwwGnRhx8f6+E901EQ80APHcOnlimKgGehat1XYP1EcNIaTxQsmtqpOk7Vwlj0b8lMk
2cBRpOGdAwK+EmKDFakQTVdbZ1O3BFBoKYVgVwh4/8vTXBdSbEPgiOdMOCj45/D+qPzIA0+l8G54
W4fqtYf4OG57qMWwxuAyMuVMorLYxtaBNxiVn93Ck06zSkKaRoaKmFPY4RyN+3en7tQqq3D41+jk
m7oBlT+w0/0EVrH9uskICZQ59dMac91VmK7VXv2y4d2LhFQqpFKhRfFjMGcaeDehWnuaytrjvCwe
sOgMIq6YS4guhuQ826q/Z6l4YRr4Z/n7o8dDtua1B1tlAlCRR0bshS/JIpdrQ8oCQ+oR1AHrnv2a
nQrHB8NuvfGdBJuovFqeZb1bUKnZ9ZSW3t/zBKZ9wFmF95Ie+VzNyYWJch7lmxefMDmfne/SSsDL
GnU/q+/7GMcEbXZ+gdmjh4tb8VGGjEtz2fUKHMsM6KyJrb2zP1F5RGrRDDeE38EPFuYxPkHe4giD
csWxGNc3YFj5d3iDWCtv5XJJe/xJ5NG4ygrSn9p8ulkfDjYQFi1zjm6J2d8S+1+ICOb+KX3JZP/i
VANk/7N+D4izi4OxtTyftiwmjC1rMy3HL3eTLrocWrN8CJ+hEI1K1zrAVr+57zMg34GSiEH98aqL
Vd8amyxAoG1bxIkWuD9n4El5NokBtZHan0ONX6o/54nwlA39vfEuogvsbuXR6aZFRg3tas2tvCJb
E5UR19u22m+iq6TjFDF0dT649jhMRs8pEZRiPhw3vXuEd+KXE+6tONNUiBbiVYOOgfxxxjivCL3W
wMo3yJvnc5YcLQqDbZP8cWXz5x6JhHP2tFzQXoNqoXBP60nM+nBpPuEwNOjy3OO8GWaSiYBaLSCh
gnStbeGaYhxPo0kjhFDusAC/ps6TphxKOiQcCXupwhHByVEMzjrbIPDrR9Iyn/9x/FA/L/pJUTWM
VQ7krHk2Fr8MVP22pvIaRYNyFmA3ZyH+CWfWt1lCC++m3d8JYEJoG2J+JGmf+zlLRSvGMSh3CYND
2q8Hlrg/bTDtX+4x9TnF6He6QneDfcjlFUTjzoO1JSqFBcCAWCMQgiv3NqSf/vYnv9BYReEiU4QQ
3V0/qvbeC3o2gzIm8AveMz7hblUlsijAI2MOfowz/KkJRNslbhaDu2+k4hqjzErZw25debt5WKKR
elwi/2W6qT1AcIq9CLP4YfgifD3d6mfWH5wff305izG9oacOWX/9zZusxBj177cosod9Tg5eDlmx
EotTh5vEF3Y8CF9Yyu2ATCPfh8rGcfrhRVl5o5WiD5lmtyZKjwDRorslBultJbkYS5OyoenZ8pTN
tk9oAdatmYSvbsHiuFFA0mfq6TEJW1NlMiNyNE3h+gg9+sHWdeehKO01lJKJSaihnpbkJ55ADdVM
pYL8foHafwgezOAY/XZLhLOp3mDUDGTzFdO7ft57aikCqedoQVQqkdn90RUoPYRnQxxqtLEIaO5K
mOOkrTtYxDCWGiuxod32DQLuVl+wxcJW7qrOw0JtXBwLUEfvvSptGivYcjjpNXlPPvXMPFKCQ58m
eB4GWFbsvU+89g26mUZ4IJlpy8PPpEzbx2S2YYUhZZLM/032HAxzeyZ337x1MatTzU8iLTRAkptL
IWAhOkRq2gAYJBoP8r0gGHKZzfB/fc3fIHzi8QBsgwZye4id2zM6nznxN85PoAVOH7Gzm87tW2dZ
AU6JZDJ0YOuohvaa1d7d5ex2uEKDnAm//1/9yHvu4c3MBZByQNGX0Yu04kZt50ucJK69V3r2PnvL
2GnK1XynVk9LqGwlMfUnVUk14WAj96ZiAnk4qktc7VTd+Eh0y5TxZQKMCb434LweehHakESP66Mm
z0fAhwKT46+vkAa0RtHCyVrJmFi6S6+XQn7xbB1q6uW1g1wGJMphz4ieL48RThZAiV2MLjXRDexI
D5ottGPQgyXKOE+i7w5RklproP8dNUIFycPUKymgHHRYDMfb0rtAYm1kIONt+AY451krujMD+E/y
HDotTvRWgmsY05nsM3FGriHlOh6hpICqdUYs2OwLUu5zBM2HeojePgvmdtJjUURFFZr1wBjDx0fm
HCXK9UC+1ryr0U/qLzsWmZieduKpCpwbrgCH5OmnGTUL1U+I54kq3waZX8sZJMNlxR7jn7pLhMfa
L2HxEudAGWHPhLIprcSlPvL/vrkDZYmGLNyZtD89Y297GYE56EJSvFIAFMozf55Ie+G0Uixyr7sR
26B//OxyTaKzgR4IvWmdxtJL3R+z/Mm6qUyEDGcSqRzs6qOXjUZHa7YSCDUZ9jCapY7SROuffySD
aKyNz5kfRPmA9SxE/eDQgq+HBAbjDyY6/VIrurMN2Umz0xYcuHEPqKJOJlThbN4mXnaadE/sBZtP
F1iGN2VuJPHL2BzrjOVbk5YtyEgFc4ec3Us4oTY09080ryTSTaD76mMbmNUKPprKWxiF8SiluNoX
OZf/jcuiIy0aTiCjDWwcbkLJCxtDLqSSn7Cat3EAnmlpgWrxhYfP0wdyVY2jKIEdW+NMT4ks4B2Y
A3KVAK1gVq66jR1X8bVM2h12CH94ExdJvfBmOaid2bsj4i/dwBVLoPIq7H8/X6qLEA6f4sZjuI0u
FyyNZ6QtFngSYiUP1SG6sKZd5EvVTsEg9/p8uXaNYgJfe/ObTdTOozuhnk1Lq3AhIdk83FdDLN66
GCnnbuG1PjP3J1n/xuHHjxtZ1fjH4s2syKK1sDpgZSEokEBuLbbDu2ULb9jIaxPr2QZLl40NFTCd
CdXnkdWB0C9sKEWl3OuktJO5hH/QKsdAUUXXQyfpt+lG7IER67FMRTr+7+MveAn80LW1NI5kcmLP
GFaNXXEOpulVO+mQAfLZRWT0agmrpC/HWTE4R507RIm4pH6TTwD2UZWpmzQvm8E/XQmrqmOLL8H7
DEvrjOZECMv+yMK+1xrGwDeMwAbJ+n8Y5c7xOEias/6/nZsRZtV8aKIk9KG/GB3IMchrxfSEeJ4u
o4T5wjZFqccJdJtgI48TP+XnxczWRKxXDxR/RDADeD9HwaM3qPPAdlbMmG201pGSy5RFyPY6Jcsx
RNsj70XNcs5DQ2OWl+AT5N6laI0zJjCxNvgl49qtUKGtoBcjBJo0yMkwH8XEqA78zjNEl7bNnZfQ
yOnVZ7M4qu1/YkGvPbcwG/PyC2MhAWzGtLZwvSDOV1RVdwVLa+N43d6+ZMRoHbf5PNW49rjATCaA
Q9boz7h3k+OcLlmmTY3eN3uDk9MjfaQs8sA0cZQkOIg2P48moXw57D4ME6IYxVlNwAnBPo3P8bIK
MDceUM5Z77bFNYh1oEonXy8hwcsiVc7b8Vklll4Px4TJ942Slg46sjj96x/0DggKGk8MUnBVEGw7
gv/sTT7TSkFgh+q8hz+q/5SZ+IbvpWEVJaN3QN8YAUF7Y4fvV1zFVXOLJxZMko9QVkfQMv7zqAyU
pA+Mb5KhakNj1Bpiri9lbbR82wG2LvV9xXpUDyf80XdW3DMAbony72X938Ng/wb6X12GQ4T56+XD
QCsbs7MV5isxu66M47li9w39Xo9J1YIoX6amb90xLkMqWYi1IVJBqAv+w9awECQAVBnx/s9STgFP
2LKgAtpm3vyQEvuIW4TvJSmsO7IY3C8DsqWaSL+6ila9+OL+UMZLGo5PS9rgZB3HxJs+gwarcuUF
ENixDIWWR1W7BXmKopGmXVm0HxRngSL2S55EMAO1ORcgER7hzpFgXsHTmu5VFzadXE/ukXR92Jdc
EB91qyXckWzKdcz5mkd7j4ey3FDQvJ0FfWQz+0FXA96t+OFUlWLLruCt10RXLWp3gXDA2LBo9i92
DfowcdEYNmuOEeaWRjUTlw57xrVNDjPIbXpq9gMTOZ249LvwznhAInWwQy9CZAUqPrYFMXzW7XJr
InsSIHaJC/jojURrNp3P+hnxUp2Q1CxUyMjvhNW+2j+X9/vCShzQvXFNpQ2pgcIEBhImOoG50Non
PT7Xh7vcKENn7ADO07NE4y3Fsa9l/IeTCCm3v85A0C7o4JeUfhM28IOsJm/yNFtVVMOrSyaT+9be
V54eJ2/PL1C2yAmdiksGv9CoTgbIu6ps/BpfRLyjiRswOSgwlr39KSDgkN88+5bD7ROsRfVAOFQc
HsVwR/Z9eIPsq8HXe0hBhHPE/5LDWaPwXRDwyT24D1T9ML8PrpO6iCd7ZXYpcg1Eno8fQAzUep03
83YpoMndp5baVe+P6VmAsM9u6q0pUVFQ9gIXrt0dLcG97BR2p5WxqEg937IGr9xNKR/oPwBuaAqY
PLJ1NNNaOXs8U4MA/JlB9BLqIGkX4ZW+uV26cEPmzYR5ZJ70BQFK7liFWvhCUaZ+R5DVT1E5qk+O
IVBt5kUB9NV/MGAh2TypEMETyk/F2UDml8pDStbgAZDG/JxCpO1xfvjjTZwY8h4cmqwL04jlTYAE
JjRHIM5hGTQs+R23Evux4uxHS8j22ERCILHOuaCRDzoxnllpYTnj+3WlnIdqOPq9IrurFenAhx++
g6zrUBVsAmfChJEmeIVDnpg8AEwr1HTK0klqNkHDwjjRqg/f/WMiD74O8KYBGueWhGywHJOqrZlc
wM2SoP5tj6WwgT1f68j5YAtln8AnhJVLJTum5/uhAczMjWCN01KF2++efI75wkLqbahqTue2s/19
6vSsETA77UJW7obEUA0fSnZti78QTg/fRTTqWkF+ydY4nwwi6ezQmVlfceXD9DdPOABlBz6buVWV
2dmCmxrPajrCBR1ayWqe5rb3mZsE6JViNgyhs+2PllD6zidwXUBv9+A5AXmtUJ01rvHSdRKJ3yxk
DbI+9ZstZMnjwptTicnJdjsepa1RsGBuAwjwJqH07i1YEECLnQ5RkiphD29k/Y2vNuKmAx8UCTT2
Ch6VB6Ur2kv/sQda5QSY+0d/rJdKHhIFdD6pqvqAPGCQ94v+0TFYfe+YSB3S7fTJFveuett5WV2C
z9UOVttTsxeFXOSsQlrfjDUFxQ4mOBDDTKLvBuCJVvUqzjGmXyF/XCj2X1WbQy6Qb1ffQWI2AMKV
BJwD3qZmNLuvMQfstK8pJhMKOVc0EWXfBqH//BQrncKJzeCpbWIgh3VhjZ/AKgpo23q+OKzP0G0z
DVVJg4p6cca+7qPrmjaoEN3tVJjenPF5eMwSe4CXWlgvhSwRabrLabAd1x0jMw1aR4dmF/Fz5KiT
e1o+0DhBE2wt9XZUAIf2aTarUVZ8weEsRsOvCbt0cFrGnA81dbecEle7HoWuq+J3s9la+ZdQHdEj
Kwnfa8wwIzc6CStWtF4tzXzc/CQYYzRbnBFhu0XqXtvCU966VhNwFqFvqskWcaWT+H+d0x/QS6WR
EDkdb5qP4PXxlOa6da0VTT2DUAhxSZCbZT9vhNdIlpPokdYy3sxmEUq9HX8YlzF7/N6Zl/ySDWVn
W/inf9RiP+4LJIxXIxQIQHFPtqUUhAk3CZhCU8U6r7nXHSEQD1QfSlUs2DzXUqc5Efcu84g2k3KV
/2SPNBbPEODdFisGs0gMrzPHO+XmEW9qSvC9RRXnjs6Ehg6FsAAIv3XqnhSeD9LMQXuNtr4plhAA
YkUrish5aPfNBMlEyUl4a+hsDmCyzHM1ehb4umq1bFbg39ag2XkGasmt2ge6xboApj1OH8m17uOQ
c9DX3xH6Pk2qf3qq2IhkPbjJ3T789WUbIbboXfGcYCr47gA1FDOPnzO0D/DdWOTi71JQw5PCakPX
Elnzkgev4jNDKLLyy17bGmkjglQpGzJMXrocFvY4ZndR08FbICOizb1WxvNLUlR7VKlbf7eKmusS
Dqh0t6fcB+ORAQv0xLZaCeCRZYtkGqJVz7AY2eSe4a4OkbIJetfCfVSb6VCVDibfnphTQyYcoe8T
5WCi2HSUSoG36w32gWgK60wBgsH2vDcsHB9q4pDWaTjJNF1itZ0qCC6aHDfAV84/KWXJPlXzHwRA
PVX+W3WgdqgWVnO6RBB8/08IVQJkW7RDDJbKClEvuIh8TEWyrKi1p5vntbkZPgJYjo5rbHszrp2w
O5JgAg9bldNH6hhwP7ajL+ptrO43dUYZlktP9/HLGdQHfGsdnzgC6vcpthnwWgb3OhnL3fdm4E2W
wO2nnIoJbN8T/g8vJKj0AvPjrLbgoboMto2bX4waGmEY0/qA1yF7qedKh8JbkskFRcydjvotGF8v
E9t2hnQ9OEJoVTYrHNVBqNmrdfVX3RKbPMQHD4Qqlc8T9VJZdGMuVWi4fe030EzJPtajv3ulJSWH
+JnIAUWs78hYvlF9WTNhHscJRTvOnH6qPJXoDSrfHfGwyRniwhjpfWyNovODgQdBLD6X/r6S+kGv
APsukHEWBG9vbLs/gFZXQ/csbgPNnX8nWwut7V9zsejPRDSIq/BlIda+YRGLX6g7ZYM/HyFd3sa5
oapfMsZRUTxRDBbF0Suh+fSVifM3TG4zA0VEDQ5mtwFG0OD7ugoXsIKDWELZQXb50uc6My8S6s/V
imPHQ3lrIvzOb1J+cku69OI1Qq7NYutiNmldXg/4Ew2U5hC02p9KWLjpCMgBKr3RdDUTUfSxGNZk
q+4KJnufiBzMIplKOUzvS2mYW6uXXwc1NBGGUpISKXjE6SAed+qtjSO36av9Agx79KPVnhZrhkkO
8lApHeyCujKHV88UBiYH+ZLAcjmn1j/8eUJAWrVnamuAy5YnJa9CSBUqdWOI6D8lweyfn1DmE6/5
2BjuAPT5jyda5LmL6s3TyNwUZdjqOG9DlBHqVpTnuBwfRPJlhn53JtboaIpSF0KIwG7Rr5ssDbpR
tux+rVIptlFDo/l8dcPMCKCPKuEM9OEiuwbRN+gpbU9sLhFySM7DhZIzC/hGRSCFblKw9oj/Xh4+
lXFBKvt6346z2TFKMY41Pu5lFILJUycPcGgxxDIhJhejZMe7sykxNOMH2wWx/gORmbVhD4m05m7s
80gIgVbX45ujvPGHKzuw06DP9bZKA6Bln/DIVPyzBGwkPHFeyD/PXipiuOezvGDN9ttaYaYYznxl
gJb1k6QjhoipnANXG32YQWTJ4P5TnlNEWRxHe63O3Azsy+eHWPA974AU6ZpK4MtCTiScKDm5id1i
iR3rr4AguHnhOb3+svGrxCKPFX6zLU99KYlUyymClk2a4PqVVfJjGu9L0nu802P4cwGb1Jojav5z
cHa+x96ng785/3uZptUhye63gDoSezwoNmQzfVYOmlWiZVVpnt91NTVtP0uYIuaNOcw2lIkZ34rz
SipCoz+8jG2wWQXsvZOtZ5AHN72VWwXCcVgPbuFphgt3kBVhQhgOuXk9FrgpXvwi4pikHpYxUjwb
vW0bfPcqLrzRYGYBTvMqJbfMHBpvShJMkawM3j67fgYloYjUODT9m9q6IzO1umAmsc68WwhS0rl9
4c/+mQ91tZJT+horg2n4TFCTJlNs8Ugy8V4IWKH29C94uzJaySWZ+F/3d1dM6fQaluYjLY68/XXD
o/b8GQxUbyyYHcOaf/cwdBzCIBbNpFJHAflQnVbEcYUlJ/BJ5j/iGV0zvLFl+SyvWpD1VK0Es9Ew
PYLe++LP4XS869d1W5EutUHjc3EXs0/ljtnqH15KQ2rMdhWk4gOtCdwETaThcx0tcmzNpEqh7yiN
QvV+hk/K6D1cEmW2qMqV/dIUOpwRVUkCfHilWIVpzA+D0vWIWNYBuIp9FYFwuvg8Y626LlASfdSA
RP3KI5v9N9kcnHQcRBxNXOuZOuXhFIRCrXcoiQI8FjkB+xngBJXKLvS/W5qVW3hdMcr9tMNBg5u7
ZLA/pgfCskVLCWfrtMFVpXKSssCZVRHIJxkxx67NlL6NM9Z70uqvdFvjwon22OMnlYnz8nakrU1e
W2g2mVgxZUpEEh/VWAwsFXpLurriRpaEi9guV1cRear4CjeqHcs++m8iV+opPrJ95axkQIBe0yVX
yJsnIrlQYiDCw1lLZ3MlETLh9Vdb6LbQ9C3Kdo25gBqkPVG6oo+CFqN+5clpAsJ3WWnzxYCA0V6p
uP5e7ScUJWtTfodJFFr07Jv7EGGpuoclTBGIDMX7EJ73gNujUh9VuXCVa8Ke0ogIiX9++kYxvEqw
m9ucZxfdoePwf1m3ColvIIukChlhT1tl50gH9xJ/CuESF4vX1KtoUn3vTaoVHQ5TsAv418WuaHG2
uqk2cZnp3YY4io/w78SRgSkA127HeqFdnmV6KjrhWp5VPw/H7bFGPDHl7TkrXhQVJYLYj/ANa6pQ
Knu9w5vtP110PrU4mm+hTLX2e2m5ZuM1oU8RXbE83Yd28QGs25UyLk8X8OR4vzYw7EFbV3+wK3d6
hBxrqx0Ze1C+KhWcRdLOEg0dH2a8IJoeiItMtpe4dSCDgpvPfFJkdfSXWaT5ditQioJqvjE94HbM
/HpU/HsSTzeL2FcK8qyGvCYmUIw2GNeZJIqwSDw0OZIOept3ts0+XyD9K6qb/LFsCXdGxkn+gzVo
IXHZ0VRVI6o9lPh1mJ/6jKTmaRRAqSeCbPreqJYlI1yp1V5Do8ECCK7ucmvPaWW84MrbwUkauwwY
c88hw9fcPJKWoKSWFe1DqYp08l+9cr8LI15x6JvQpznFdRMsUAGww0XiaLIf53urrOcNouSNT2rO
ZS/0w652U+QZI5Q6K/Z6h7ynnFqiVV93Sh3168fxQL4vxjSs5YaHyb3r0wdUVxMxy7hGbvZSMndG
JOxMyYOBVaCaoYchvsbxTjD9j8jyasEls5goow957RrOMnSttRYmJIFJQFsJ1koSo2g3hFwqJah4
XnAcGOpQbzSePW17qzjs7BiIC4IbQ2AbD/JK6InxlnaDNMSvTaN7yhtj9TDs/94XDW1eJ94q20KE
JzWeqAKbR8JTYCnubjYZk4T0nMe3JFFFFAvT+ghKxDQY9Y2QA6UsRmiztKHXyJfBoCocKjR/6PC8
UPV21Wm7YumxeHZB7O+XxFnYUWKkDChS4Mm9uxR0y7QQW+gbMPTo3APm8T5lvvB4K55Hzr9bfwrX
H1+obdtBQY/k1Io7iM3r2q+R4K66N0mkxWlw9sJ7+AT9/dfeA4Y9rgxkP1swN+JQ9vThN4HxEIia
qA1rIuPj6iSDO97Gd+2P3L666NXGObATG9EQKQNz70F5D+pIYyDrmJY/1cWwFNObNVRkiFmZRXCc
m2B6c8cVaZddP63O3G5+GazIe+Lr6TzZmuMcJnDxRO3fryGhknOsJn9NbjDLtOxnqPxWDYd1K9wM
zHKrpnj6cB3PqIGavhOG6M8jXt6md3uAGYUSQyIR/KmgpXnzUPy3ojQZa0f6W26FRydx4jHfh+y9
NlzqnPYGpgDg/500fBjYUKBlP4fKaOxCMKqrpQdWuDt3pKMJO8BCtC5DbtAm+OfMAXmqhub6Qbo8
h7f4d65BK+tlFuvhwxIrJM6MXv4N3l1oc0Nh3LliiDFoBN6HAyF5JUD7bb3acS2rrJcVjcam9+E6
bOPpY9ED5IyJIIh76f8lQPhQqMpvlMhPyjm1n8s36CCV3OWtakCKPhzY9HHM/q3g1LM9YtbJY3Be
Io7NV/VJLY6hR9/Y9EVSQ88Ue+kmhYjwDHO46FvHszHmIxHoC7gISPDHgDaLZ/LbKVATMclut2Gq
Goqd5WlypBbeb6ytRtdJKN7gbrf4
`protect end_protected

